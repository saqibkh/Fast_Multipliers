module multiplier_64bits_version12(product, A, B);

    output [127:0] product;
    input [63:0] A, B;

    /*
     * Area: 89115.374260
     * Power: 77.2476mW
     * Timing: 8.51ns
     */

    wire [63:0] pp0;
    wire [63:0] pp1;
    wire [63:0] pp2;
    wire [63:0] pp3;
    wire [63:0] pp4;
    wire [63:0] pp5;
    wire [63:0] pp6;
    wire [63:0] pp7;
    wire [63:0] pp8;
    wire [63:0] pp9;
    wire [63:0] pp10;
    wire [63:0] pp11;
    wire [63:0] pp12;
    wire [63:0] pp13;
    wire [63:0] pp14;
    wire [63:0] pp15;
    wire [63:0] pp16;
    wire [63:0] pp17;
    wire [63:0] pp18;
    wire [63:0] pp19;
    wire [63:0] pp20;
    wire [63:0] pp21;
    wire [63:0] pp22;
    wire [63:0] pp23;
    wire [63:0] pp24;
    wire [63:0] pp25;
    wire [63:0] pp26;
    wire [63:0] pp27;
    wire [63:0] pp28;
    wire [63:0] pp29;
    wire [63:0] pp30;
    wire [63:0] pp31;
    wire [63:0] pp32;
    wire [63:0] pp33;
    wire [63:0] pp34;
    wire [63:0] pp35;
    wire [63:0] pp36;
    wire [63:0] pp37;
    wire [63:0] pp38;
    wire [63:0] pp39;
    wire [63:0] pp40;
    wire [63:0] pp41;
    wire [63:0] pp42;
    wire [63:0] pp43;
    wire [63:0] pp44;
    wire [63:0] pp45;
    wire [63:0] pp46;
    wire [63:0] pp47;
    wire [63:0] pp48;
    wire [63:0] pp49;
    wire [63:0] pp50;
    wire [63:0] pp51;
    wire [63:0] pp52;
    wire [63:0] pp53;
    wire [63:0] pp54;
    wire [63:0] pp55;
    wire [63:0] pp56;
    wire [63:0] pp57;
    wire [63:0] pp58;
    wire [63:0] pp59;
    wire [63:0] pp60;
    wire [63:0] pp61;
    wire [63:0] pp62;
    wire [63:0] pp63;


    assign pp0 = A[0] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp1 = A[1] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp2 = A[2] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp3 = A[3] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp4 = A[4] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp5 = A[5] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp6 = A[6] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp7 = A[7] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp8 = A[8] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp9 = A[9] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp10 = A[10] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp11 = A[11] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp12 = A[12] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp13 = A[13] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp14 = A[14] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp15 = A[15] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp16 = A[16] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp17 = A[17] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp18 = A[18] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp19 = A[19] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp20 = A[20] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp21 = A[21] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp22 = A[22] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp23 = A[23] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp24 = A[24] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp25 = A[25] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp26 = A[26] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp27 = A[27] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp28 = A[28] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp29 = A[29] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp30 = A[30] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp31 = A[31] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp32 = A[32] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp33 = A[33] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp34 = A[34] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp35 = A[35] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp36 = A[36] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp37 = A[37] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp38 = A[38] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp39 = A[39] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp40 = A[40] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp41 = A[41] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp42 = A[42] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp43 = A[43] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp44 = A[44] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp45 = A[45] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp46 = A[46] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp47 = A[47] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp48 = A[48] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp49 = A[49] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp50 = A[50] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp51 = A[51] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp52 = A[52] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp53 = A[53] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp54 = A[54] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp55 = A[55] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp56 = A[56] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp57 = A[57] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp58 = A[58] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp59 = A[59] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp60 = A[60] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp61 = A[61] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp62 = A[62] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp63 = A[63] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;


    /*Stage 1*/
    wire[3:0] s1, in1_1, in1_2;
    wire c1;
    assign in1_1 = {pp0[38],pp0[39],pp0[40],pp0[41]};
    assign in1_2 = {pp1[37],pp1[38],pp1[39],pp1[40]};
    CLA_4 KS_1(s1, c1, in1_1, in1_2);
    wire[3:0] s2, in2_1, in2_2;
    wire c2;
    assign in2_1 = {pp2[37],pp2[38],pp2[39],pp0[42]};
    assign in2_2 = {pp3[36],pp3[37],pp3[38],pp1[41]};
    CLA_4 KS_2(s2, c2, in2_1, in2_2);
    wire[3:0] s3, in3_1, in3_2;
    wire c3;
    assign in3_1 = {pp4[36],pp4[37],pp2[40],pp0[43]};
    assign in3_2 = {pp5[35],pp5[36],pp3[39],pp1[42]};
    CLA_4 KS_3(s3, c3, in3_1, in3_2);
    wire[3:0] s4, in4_1, in4_2;
    wire c4;
    assign in4_1 = {pp6[35],pp4[38],pp2[41],pp0[44]};
    assign in4_2 = {pp7[34],pp5[37],pp3[40],pp1[43]};
    CLA_4 KS_4(s4, c4, in4_1, in4_2);
    wire[3:0] s5, in5_1, in5_2;
    wire c5;
    assign in5_1 = {pp6[36],pp4[39],pp2[42],pp0[45]};
    assign in5_2 = {pp7[35],pp5[38],pp3[41],pp1[44]};
    CLA_4 KS_5(s5, c5, in5_1, in5_2);
    wire[3:0] s6, in6_1, in6_2;
    wire c6;
    assign in6_1 = {pp9[33],pp6[37],pp4[40],pp2[43]};
    assign in6_2 = {pp10[32],pp7[36],pp5[39],pp3[42]};
    CLA_4_c KS_6(s6, c6, in6_1, in6_2, pp8[34]);
    wire[3:0] s7, in7_1, in7_2;
    wire c7;
    assign in7_1 = {pp8[35],pp6[38],pp4[41],pp0[46]};
    assign in7_2 = {pp9[34],pp7[37],pp5[40],pp1[45]};
    CLA_4 KS_7(s7, c7, in7_1, in7_2);
    wire[3:0] s8, in8_1, in8_2;
    wire c8;
    assign in8_1 = {pp11[32],pp8[36],pp6[39],pp2[44]};
    assign in8_2 = {pp12[31],pp9[35],pp7[38],pp3[43]};
    CLA_4_c KS_8(s8, c8, in8_1, in8_2, pp10[33]);
    wire[3:0] s9, in9_1, in9_2;
    wire c9;
    assign in9_1 = {pp10[34],pp8[37],pp4[42],pp0[47]};
    assign in9_2 = {pp11[33],pp9[36],pp5[41],pp1[46]};
    CLA_4 KS_9(s9, c9, in9_1, in9_2);
    wire[3:0] s10, in10_1, in10_2;
    wire c10;
    assign in10_1 = {pp13[31],pp10[35],pp6[40],pp2[45]};
    assign in10_2 = {pp14[30],pp11[34],pp7[39],pp3[44]};
    CLA_4_c KS_10(s10, c10, in10_1, in10_2, pp12[32]);
    wire[3:0] s11, in11_1, in11_2;
    wire c11;
    assign in11_1 = {pp12[33],pp8[38],pp4[43],pp0[48]};
    assign in11_2 = {pp13[32],pp9[37],pp5[42],pp1[47]};
    CLA_4 KS_11(s11, c11, in11_1, in11_2);
    wire[3:0] s12, in12_1, in12_2;
    wire c12;
    assign in12_1 = {pp15[30],pp10[36],pp6[41],pp2[46]};
    assign in12_2 = {pp16[29],pp11[35],pp7[40],pp3[45]};
    CLA_4_c KS_12(s12, c12, in12_1, in12_2, pp14[31]);
    wire[3:0] s13, in13_1, in13_2;
    wire c13;
    assign in13_1 = {pp12[34],pp8[39],pp4[44],pp0[49]};
    assign in13_2 = {pp13[33],pp9[38],pp5[43],pp1[48]};
    CLA_4 KS_13(s13, c13, in13_1, in13_2);
    wire[3:0] s14, in14_1, in14_2;
    wire c14;
    assign in14_1 = {pp14[32],pp10[37],pp6[42],pp2[47]};
    assign in14_2 = {pp15[31],pp11[36],pp7[41],pp3[46]};
    CLA_4 KS_14(s14, c14, in14_1, in14_2);
    wire[3:0] s15, in15_1, in15_2;
    wire c15;
    assign in15_1 = {pp16[30],pp12[35],pp8[40],pp4[45]};
    assign in15_2 = {pp17[29],pp13[34],pp9[39],pp5[44]};
    CLA_4 KS_15(s15, c15, in15_1, in15_2);
    wire[3:0] s16, in16_1, in16_2;
    wire c16;
    assign in16_1 = {pp19[27],pp14[33],pp10[38],pp6[43]};
    assign in16_2 = {pp20[26],pp15[32],pp11[37],pp7[42]};
    CLA_4_c KS_16(s16, c16, in16_1, in16_2, pp18[28]);
    wire[3:0] s17, in17_1, in17_2;
    wire c17;
    assign in17_1 = {pp16[31],pp12[36],pp8[41],pp0[50]};
    assign in17_2 = {pp17[30],pp13[35],pp9[40],pp1[49]};
    CLA_4 KS_17(s17, c17, in17_1, in17_2);
    wire[3:0] s18, in18_1, in18_2;
    wire c18;
    assign in18_1 = {pp18[29],pp14[34],pp10[39],pp2[48]};
    assign in18_2 = {pp19[28],pp15[33],pp11[38],pp3[47]};
    CLA_4 KS_18(s18, c18, in18_1, in18_2);
    wire[3:0] s19, in19_1, in19_2;
    wire c19;
    assign in19_1 = {pp21[26],pp16[32],pp12[37],pp4[46]};
    assign in19_2 = {pp22[25],pp17[31],pp13[36],pp5[45]};
    CLA_4_c KS_19(s19, c19, in19_1, in19_2, pp20[27]);
    wire[3:0] s20, in20_1, in20_2;
    wire c20;
    assign in20_1 = {pp18[30],pp14[35],pp6[44],pp0[51]};
    assign in20_2 = {pp19[29],pp15[34],pp7[43],pp1[50]};
    CLA_4 KS_20(s20, c20, in20_1, in20_2);
    wire[3:0] s21, in21_1, in21_2;
    wire c21;
    assign in21_1 = {pp20[28],pp16[33],pp8[42],pp2[49]};
    assign in21_2 = {pp21[27],pp17[32],pp9[41],pp3[48]};
    CLA_4 KS_21(s21, c21, in21_1, in21_2);
    wire[3:0] s22, in22_1, in22_2;
    wire c22;
    assign in22_1 = {pp23[25],pp18[31],pp10[40],pp4[47]};
    assign in22_2 = {pp24[24],pp19[30],pp11[39],pp5[46]};
    CLA_4_c KS_22(s22, c22, in22_1, in22_2, pp22[26]);
    wire[3:0] s23, in23_1, in23_2;
    wire c23;
    assign in23_1 = {pp20[29],pp12[38],pp6[45],pp0[52]};
    assign in23_2 = {pp21[28],pp13[37],pp7[44],pp1[51]};
    CLA_4 KS_23(s23, c23, in23_1, in23_2);
    wire[3:0] s24, in24_1, in24_2;
    wire c24;
    assign in24_1 = {pp22[27],pp14[36],pp8[43],pp2[50]};
    assign in24_2 = {pp23[26],pp15[35],pp9[42],pp3[49]};
    CLA_4 KS_24(s24, c24, in24_1, in24_2);
    wire[3:0] s25, in25_1, in25_2;
    wire c25;
    assign in25_1 = {pp25[24],pp16[34],pp10[41],pp4[48]};
    assign in25_2 = {pp26[23],pp17[33],pp11[40],pp5[47]};
    CLA_4_c KS_25(s25, c25, in25_1, in25_2, pp24[25]);
    wire[3:0] s26, in26_1, in26_2;
    wire c26;
    assign in26_1 = {pp18[32],pp12[39],pp6[46],pp0[53]};
    assign in26_2 = {pp19[31],pp13[38],pp7[45],pp1[52]};
    CLA_4 KS_26(s26, c26, in26_1, in26_2);
    wire[3:0] s27, in27_1, in27_2;
    wire c27;
    assign in27_1 = {pp20[30],pp14[37],pp8[44],pp2[51]};
    assign in27_2 = {pp21[29],pp15[36],pp9[43],pp3[50]};
    CLA_4 KS_27(s27, c27, in27_1, in27_2);
    wire[3:0] s28, in28_1, in28_2;
    wire c28;
    assign in28_1 = {pp22[28],pp16[35],pp10[42],pp4[49]};
    assign in28_2 = {pp23[27],pp17[34],pp11[41],pp5[48]};
    CLA_4 KS_28(s28, c28, in28_1, in28_2);
    wire[3:0] s29, in29_1, in29_2;
    wire c29;
    assign in29_1 = {pp24[26],pp18[33],pp12[40],pp6[47]};
    assign in29_2 = {pp25[25],pp19[32],pp13[39],pp7[46]};
    CLA_4 KS_29(s29, c29, in29_1, in29_2);
    wire[3:0] s30, in30_1, in30_2;
    wire c30;
    assign in30_1 = {pp26[24],pp20[31],pp14[38],pp8[45]};
    assign in30_2 = {pp27[23],pp21[30],pp15[37],pp9[44]};
    CLA_4 KS_30(s30, c30, in30_1, in30_2);
    wire[3:0] s31, in31_1, in31_2;
    wire c31;
    assign in31_1 = {pp28[22],pp22[29],pp16[36],pp10[43]};
    assign in31_2 = {pp29[21],pp23[28],pp17[35],pp11[42]};
    CLA_4 KS_31(s31, c31, in31_1, in31_2);
    wire[3:0] s32, in32_1, in32_2;
    wire c32;
    assign in32_1 = {pp31[19],pp24[27],pp18[34],pp12[41]};
    assign in32_2 = {pp32[18],pp25[26],pp19[33],pp13[40]};
    CLA_4_c KS_32(s32, c32, in32_1, in32_2, pp30[20]);
    wire[3:0] s33, in33_1, in33_2;
    wire c33;
    assign in33_1 = {pp26[25],pp20[32],pp14[39],pp0[54]};
    assign in33_2 = {pp27[24],pp21[31],pp15[38],pp1[53]};
    CLA_4 KS_33(s33, c33, in33_1, in33_2);
    wire[3:0] s34, in34_1, in34_2;
    wire c34;
    assign in34_1 = {pp28[23],pp22[30],pp16[37],pp2[52]};
    assign in34_2 = {pp29[22],pp23[29],pp17[36],pp3[51]};
    CLA_4 KS_34(s34, c34, in34_1, in34_2);
    wire[3:0] s35, in35_1, in35_2;
    wire c35;
    assign in35_1 = {pp31[20],pp24[28],pp18[35],pp4[50]};
    assign in35_2 = {pp32[19],pp25[27],pp19[34],pp5[49]};
    CLA_4_c KS_35(s35, c35, in35_1, in35_2, pp30[21]);
    wire[3:0] s36, in36_1, in36_2;
    wire c36;
    assign in36_1 = {pp26[26],pp20[33],pp6[48],pp0[55]};
    assign in36_2 = {pp27[25],pp21[32],pp7[47],pp1[54]};
    CLA_4 KS_36(s36, c36, in36_1, in36_2);
    wire[3:0] s37, in37_1, in37_2;
    wire c37;
    assign in37_1 = {pp28[24],pp22[31],pp8[46],pp2[53]};
    assign in37_2 = {pp29[23],pp23[30],pp9[45],pp3[52]};
    CLA_4 KS_37(s37, c37, in37_1, in37_2);
    wire[3:0] s38, in38_1, in38_2;
    wire c38;
    assign in38_1 = {pp30[22],pp24[29],pp10[44],pp4[51]};
    assign in38_2 = {pp31[21],pp25[28],pp11[43],pp5[50]};
    CLA_4 KS_38(s38, c38, in38_1, in38_2);
    wire[3:0] s39, in39_1, in39_2;
    wire c39;
    assign in39_1 = {pp33[19],pp26[27],pp12[42],pp6[49]};
    assign in39_2 = {pp34[18],pp27[26],pp13[41],pp7[48]};
    CLA_4_c KS_39(s39, c39, in39_1, in39_2, pp32[20]);
    wire[3:0] s40, in40_1, in40_2;
    wire c40;
    assign in40_1 = {pp28[25],pp14[40],pp8[47],pp0[56]};
    assign in40_2 = {pp29[24],pp15[39],pp9[46],pp1[55]};
    CLA_4 KS_40(s40, c40, in40_1, in40_2);
    wire[3:0] s41, in41_1, in41_2;
    wire c41;
    assign in41_1 = {pp30[23],pp16[38],pp10[45],pp2[54]};
    assign in41_2 = {pp31[22],pp17[37],pp11[44],pp3[53]};
    CLA_4 KS_41(s41, c41, in41_1, in41_2);
    wire[3:0] s42, in42_1, in42_2;
    wire c42;
    assign in42_1 = {pp32[21],pp18[36],pp12[43],pp4[52]};
    assign in42_2 = {pp33[20],pp19[35],pp13[42],pp5[51]};
    CLA_4 KS_42(s42, c42, in42_1, in42_2);
    wire[3:0] s43, in43_1, in43_2;
    wire c43;
    assign in43_1 = {pp35[18],pp20[34],pp14[41],pp6[50]};
    assign in43_2 = {pp36[17],pp21[33],pp15[40],pp7[49]};
    CLA_4_c KS_43(s43, c43, in43_1, in43_2, pp34[19]);
    wire[3:0] s44, in44_1, in44_2;
    wire c44;
    assign in44_1 = {pp22[32],pp16[39],pp8[48],pp0[57]};
    assign in44_2 = {pp23[31],pp17[38],pp9[47],pp1[56]};
    CLA_4 KS_44(s44, c44, in44_1, in44_2);
    wire[3:0] s45, in45_1, in45_2;
    wire c45;
    assign in45_1 = {pp24[30],pp18[37],pp10[46],pp2[55]};
    assign in45_2 = {pp25[29],pp19[36],pp11[45],pp3[54]};
    CLA_4 KS_45(s45, c45, in45_1, in45_2);
    wire[3:0] s46, in46_1, in46_2;
    wire c46;
    assign in46_1 = {pp26[28],pp20[35],pp12[44],pp4[53]};
    assign in46_2 = {pp27[27],pp21[34],pp13[43],pp5[52]};
    CLA_4 KS_46(s46, c46, in46_1, in46_2);
    wire[3:0] s47, in47_1, in47_2;
    wire c47;
    assign in47_1 = {pp28[26],pp22[33],pp14[42],pp6[51]};
    assign in47_2 = {pp29[25],pp23[32],pp15[41],pp7[50]};
    CLA_4 KS_47(s47, c47, in47_1, in47_2);
    wire[3:0] s48, in48_1, in48_2;
    wire c48;
    assign in48_1 = {pp30[24],pp24[31],pp16[40],pp8[49]};
    assign in48_2 = {pp31[23],pp25[30],pp17[39],pp9[48]};
    CLA_4 KS_48(s48, c48, in48_1, in48_2);
    wire[3:0] s49, in49_1, in49_2;
    wire c49;
    assign in49_1 = {pp32[22],pp26[29],pp18[38],pp10[47]};
    assign in49_2 = {pp33[21],pp27[28],pp19[37],pp11[46]};
    CLA_4 KS_49(s49, c49, in49_1, in49_2);
    wire[3:0] s50, in50_1, in50_2;
    wire c50;
    assign in50_1 = {pp34[20],pp28[27],pp20[36],pp12[45]};
    assign in50_2 = {pp35[19],pp29[26],pp21[35],pp13[44]};
    CLA_4 KS_50(s50, c50, in50_1, in50_2);
    wire[3:0] s51, in51_1, in51_2;
    wire c51;
    assign in51_1 = {pp36[18],pp30[25],pp22[34],pp14[43]};
    assign in51_2 = {pp37[17],pp31[24],pp23[33],pp15[42]};
    CLA_4 KS_51(s51, c51, in51_1, in51_2);
    wire[3:0] s52, in52_1, in52_2;
    wire c52;
    assign in52_1 = {pp38[16],pp32[23],pp24[32],pp16[41]};
    assign in52_2 = {pp39[15],pp33[22],pp25[31],pp17[40]};
    CLA_4 KS_52(s52, c52, in52_1, in52_2);
    wire[3:0] s53, in53_1, in53_2;
    wire c53;
    assign in53_1 = {pp40[14],pp34[21],pp26[30],pp18[39]};
    assign in53_2 = {pp41[13],pp35[20],pp27[29],pp19[38]};
    CLA_4 KS_53(s53, c53, in53_1, in53_2);
    wire[3:0] s54, in54_1, in54_2;
    wire c54;
    assign in54_1 = {pp42[12],pp36[19],pp28[28],pp20[37]};
    assign in54_2 = {pp43[11],pp37[18],pp29[27],pp21[36]};
    CLA_4 KS_54(s54, c54, in54_1, in54_2);
    wire[3:0] s55, in55_1, in55_2;
    wire c55;
    assign in55_1 = {pp45[9],pp38[17],pp30[26],pp22[35]};
    assign in55_2 = {pp46[8],pp39[16],pp31[25],pp23[34]};
    CLA_4_c KS_55(s55, c55, in55_1, in55_2, pp44[10]);
    wire[3:0] s56, in56_1, in56_2;
    wire c56;
    assign in56_1 = {pp40[15],pp32[24],pp24[33],pp0[58]};
    assign in56_2 = {pp41[14],pp33[23],pp25[32],pp1[57]};
    CLA_4 KS_56(s56, c56, in56_1, in56_2);
    wire[3:0] s57, in57_1, in57_2;
    wire c57;
    assign in57_1 = {pp34[22],pp26[31],pp2[56],pp0[59]};
    assign in57_2 = {pp35[21],pp27[30],pp3[55],pp1[58]};
    CLA_4 KS_57(s57, c57, in57_1, in57_2);
    wire[3:0] s58, in58_1, in58_2;
    wire c58;
    assign in58_1 = {pp36[20],pp28[29],pp4[54],pp2[57]};
    assign in58_2 = {pp37[19],pp29[28],pp5[53],pp3[56]};
    CLA_4 KS_58(s58, c58, in58_1, in58_2);
    wire[3:0] s59, in59_1, in59_2;
    wire c59;
    assign in59_1 = {pp38[18],pp30[27],pp6[52],pp4[55]};
    assign in59_2 = {pp39[17],pp31[26],pp7[51],pp5[54]};
    CLA_4 KS_59(s59, c59, in59_1, in59_2);
    wire[3:0] s60, in60_1, in60_2;
    wire c60;
    assign in60_1 = {pp40[16],pp32[25],pp8[50],pp6[53]};
    assign in60_2 = {pp41[15],pp33[24],pp9[49],pp7[52]};
    CLA_4 KS_60(s60, c60, in60_1, in60_2);
    wire[3:0] s61, in61_1, in61_2;
    wire c61;
    assign in61_1 = {pp43[13],pp34[23],pp10[48],pp8[51]};
    assign in61_2 = {pp44[12],pp35[22],pp11[47],pp9[50]};
    CLA_4_c KS_61(s61, c61, in61_1, in61_2, pp42[14]);
    wire[3:0] s62, in62_1, in62_2;
    wire c62;
    assign in62_1 = {pp36[21],pp12[46],pp10[49],pp0[60]};
    assign in62_2 = {pp37[20],pp13[45],pp11[48],pp1[59]};
    CLA_4 KS_62(s62, c62, in62_1, in62_2);
    wire[3:0] s63, in63_1, in63_2;
    wire c63;
    assign in63_1 = {pp38[19],pp14[44],pp12[47],pp2[58]};
    assign in63_2 = {pp39[18],pp15[43],pp13[46],pp3[57]};
    CLA_4 KS_63(s63, c63, in63_1, in63_2);
    wire[3:0] s64, in64_1, in64_2;
    wire c64;
    assign in64_1 = {pp40[17],pp16[42],pp14[45],pp4[56]};
    assign in64_2 = {pp41[16],pp17[41],pp15[44],pp5[55]};
    CLA_4 KS_64(s64, c64, in64_1, in64_2);
    wire[3:0] s65, in65_1, in65_2;
    wire c65;
    assign in65_1 = {pp42[15],pp18[40],pp16[43],pp6[54]};
    assign in65_2 = {pp43[14],pp19[39],pp17[42],pp7[53]};
    CLA_4 KS_65(s65, c65, in65_1, in65_2);
    wire[3:0] s66, in66_1, in66_2;
    wire c66;
    assign in66_1 = {pp45[12],pp20[38],pp18[41],pp8[52]};
    assign in66_2 = {pp46[11],pp21[37],pp19[40],pp9[51]};
    CLA_4_c KS_66(s66, c66, in66_1, in66_2, pp44[13]);
    wire[3:0] s67, in67_1, in67_2;
    wire c67;
    assign in67_1 = {pp22[36],pp20[39],pp10[50],pp0[61]};
    assign in67_2 = {pp23[35],pp21[38],pp11[49],pp1[60]};
    CLA_4 KS_67(s67, c67, in67_1, in67_2);
    wire[3:0] s68, in68_1, in68_2;
    wire c68;
    assign in68_1 = {pp24[34],pp22[37],pp12[48],pp2[59]};
    assign in68_2 = {pp25[33],pp23[36],pp13[47],pp3[58]};
    CLA_4 KS_68(s68, c68, in68_1, in68_2);
    wire[3:0] s69, in69_1, in69_2;
    wire c69;
    assign in69_1 = {pp26[32],pp24[35],pp14[46],pp4[57]};
    assign in69_2 = {pp27[31],pp25[34],pp15[45],pp5[56]};
    CLA_4 KS_69(s69, c69, in69_1, in69_2);
    wire[3:0] s70, in70_1, in70_2;
    wire c70;
    assign in70_1 = {pp28[30],pp26[33],pp16[44],pp6[55]};
    assign in70_2 = {pp29[29],pp27[32],pp17[43],pp7[54]};
    CLA_4 KS_70(s70, c70, in70_1, in70_2);
    wire[3:0] s71, in71_1, in71_2;
    wire c71;
    assign in71_1 = {pp30[28],pp28[31],pp18[42],pp8[53]};
    assign in71_2 = {pp31[27],pp29[30],pp19[41],pp9[52]};
    CLA_4 KS_71(s71, c71, in71_1, in71_2);
    wire[3:0] s72, in72_1, in72_2;
    wire c72;
    assign in72_1 = {pp32[26],pp30[29],pp20[40],pp10[51]};
    assign in72_2 = {pp33[25],pp31[28],pp21[39],pp11[50]};
    CLA_4 KS_72(s72, c72, in72_1, in72_2);
    wire[3:0] s73, in73_1, in73_2;
    wire c73;
    assign in73_1 = {pp34[24],pp32[27],pp22[38],pp12[49]};
    assign in73_2 = {pp35[23],pp33[26],pp23[37],pp13[48]};
    CLA_4 KS_73(s73, c73, in73_1, in73_2);
    wire[3:0] s74, in74_1, in74_2;
    wire c74;
    assign in74_1 = {pp36[22],pp34[25],pp24[36],pp14[47]};
    assign in74_2 = {pp37[21],pp35[24],pp25[35],pp15[46]};
    CLA_4 KS_74(s74, c74, in74_1, in74_2);
    wire[3:0] s75, in75_1, in75_2;
    wire c75;
    assign in75_1 = {pp38[20],pp36[23],pp26[34],pp16[45]};
    assign in75_2 = {pp39[19],pp37[22],pp27[33],pp17[44]};
    CLA_4 KS_75(s75, c75, in75_1, in75_2);
    wire[3:0] s76, in76_1, in76_2;
    wire c76;
    assign in76_1 = {pp40[18],pp38[21],pp28[32],pp18[43]};
    assign in76_2 = {pp41[17],pp39[20],pp29[31],pp19[42]};
    CLA_4 KS_76(s76, c76, in76_1, in76_2);
    wire[3:0] s77, in77_1, in77_2;
    wire c77;
    assign in77_1 = {pp42[16],pp40[19],pp30[30],pp20[41]};
    assign in77_2 = {pp43[15],pp41[18],pp31[29],pp21[40]};
    CLA_4 KS_77(s77, c77, in77_1, in77_2);
    wire[3:0] s78, in78_1, in78_2;
    wire c78;
    assign in78_1 = {pp44[14],pp42[17],pp32[28],pp22[39]};
    assign in78_2 = {pp45[13],pp43[16],pp33[27],pp23[38]};
    CLA_4 KS_78(s78, c78, in78_1, in78_2);
    wire[3:0] s79, in79_1, in79_2;
    wire c79;
    assign in79_1 = {pp46[12],pp44[15],pp34[26],pp24[37]};
    assign in79_2 = {pp47[11],pp45[14],pp35[25],pp25[36]};
    CLA_4 KS_79(s79, c79, in79_1, in79_2);
    wire[3:0] s80, in80_1, in80_2;
    wire c80;
    assign in80_1 = {pp48[10],pp46[13],pp36[24],pp26[35]};
    assign in80_2 = {pp49[9],pp47[12],pp37[23],pp27[34]};
    CLA_4 KS_80(s80, c80, in80_1, in80_2);
    wire[0:0] s81, in81_1, in81_2;
    wire c81;
    assign in81_1 = {pp50[8]};
    assign in81_2 = {pp51[7]};
    Half_Adder KS_81(s81, c81, in81_1, in81_2);
    wire[3:0] s82, in82_1, in82_2;
    wire c82;
    assign in82_1 = {pp52[6],pp48[11],pp38[22],pp28[33]};
    assign in82_2 = {pp53[5],pp49[10],pp39[21],pp29[32]};
    CLA_4 KS_82(s82, c82, in82_1, in82_2);
    wire[0:0] s83, in83_1, in83_2;
    wire c83;
    assign in83_1 = {pp54[4]};
    assign in83_2 = {pp55[3]};
    Half_Adder KS_83(s83, c83, in83_1, in83_2);
    wire[3:0] s84, in84_1, in84_2;
    wire c84;
    assign in84_1 = {pp56[2],pp50[9],pp40[20],pp30[31]};
    assign in84_2 = {pp57[1],pp51[8],pp41[19],pp31[30]};
    CLA_4 KS_84(s84, c84, in84_1, in84_2);
    wire[0:0] s85, in85_1, in85_2;
    wire c85;
    assign in85_1 = {pp58[0]};
    assign in85_2 = {c44};
    Half_Adder KS_85(s85, c85, in85_1, in85_2);
    wire[3:0] s86, in86_1, in86_2;
    wire c86;
    assign in86_1 = {c45,pp52[7],pp42[18],pp32[29]};
    assign in86_2 = {c46,pp53[6],pp43[17],pp33[28]};
    CLA_4 KS_86(s86, c86, in86_1, in86_2);
    wire[0:0] s87, in87_1, in87_2;
    wire c87;
    assign in87_1 = {c48};
    assign in87_2 = {c49};
    Full_Adder KS_87(s87, c87, in87_1, in87_2, c47);
    wire[3:0] s88, in88_1, in88_2;
    wire c88;
    assign in88_1 = {pp44[16],pp34[27],pp0[62],pp0[63]};
    assign in88_2 = {pp45[15],pp35[26],pp1[61],pp1[62]};
    CLA_4 KS_88(s88, c88, in88_1, in88_2);
    wire[3:0] s89, in89_1, in89_2;
    wire c89;
    assign in89_1 = {pp46[14],pp36[25],pp2[60],pp2[61]};
    assign in89_2 = {pp47[13],pp37[24],pp3[59],pp3[60]};
    CLA_4 KS_89(s89, c89, in89_1, in89_2);
    wire[3:0] s90, in90_1, in90_2;
    wire c90;
    assign in90_1 = {pp48[12],pp38[23],pp4[58],pp4[59]};
    assign in90_2 = {pp49[11],pp39[22],pp5[57],pp5[58]};
    CLA_4 KS_90(s90, c90, in90_1, in90_2);
    wire[3:0] s91, in91_1, in91_2;
    wire c91;
    assign in91_1 = {pp50[10],pp40[21],pp6[56],pp6[57]};
    assign in91_2 = {pp51[9],pp41[20],pp7[55],pp7[56]};
    CLA_4 KS_91(s91, c91, in91_1, in91_2);
    wire[3:0] s92, in92_1, in92_2;
    wire c92;
    assign in92_1 = {pp53[7],pp42[19],pp8[54],pp8[55]};
    assign in92_2 = {pp54[6],pp43[18],pp9[53],pp9[54]};
    CLA_4_c KS_92(s92, c92, in92_1, in92_2, pp52[8]);
    wire[3:0] s93, in93_1, in93_2;
    wire c93;
    assign in93_1 = {pp44[17],pp10[52],pp10[53],pp1[63]};
    assign in93_2 = {pp45[16],pp11[51],pp11[52],pp2[62]};
    CLA_4 KS_93(s93, c93, in93_1, in93_2);
    wire[3:0] s94, in94_1, in94_2;
    wire c94;
    assign in94_1 = {pp46[15],pp12[50],pp12[51],pp3[61]};
    assign in94_2 = {pp47[14],pp13[49],pp13[50],pp4[60]};
    CLA_4 KS_94(s94, c94, in94_1, in94_2);
    wire[3:0] s95, in95_1, in95_2;
    wire c95;
    assign in95_1 = {pp48[13],pp14[48],pp14[49],pp5[59]};
    assign in95_2 = {pp49[12],pp15[47],pp15[48],pp6[58]};
    CLA_4 KS_95(s95, c95, in95_1, in95_2);
    wire[3:0] s96, in96_1, in96_2;
    wire c96;
    assign in96_1 = {pp50[11],pp16[46],pp16[47],pp7[57]};
    assign in96_2 = {pp51[10],pp17[45],pp17[46],pp8[56]};
    CLA_4 KS_96(s96, c96, in96_1, in96_2);
    wire[3:0] s97, in97_1, in97_2;
    wire c97;
    assign in97_1 = {pp52[9],pp18[44],pp18[45],pp9[55]};
    assign in97_2 = {pp53[8],pp19[43],pp19[44],pp10[54]};
    CLA_4 KS_97(s97, c97, in97_1, in97_2);
    wire[3:0] s98, in98_1, in98_2;
    wire c98;
    assign in98_1 = {pp55[6],pp20[42],pp20[43],pp11[53]};
    assign in98_2 = {pp56[5],pp21[41],pp21[42],pp12[52]};
    CLA_4_c KS_98(s98, c98, in98_1, in98_2, pp54[7]);
    wire[3:0] s99, in99_1, in99_2;
    wire c99;
    assign in99_1 = {pp22[40],pp22[41],pp13[51],pp2[63]};
    assign in99_2 = {pp23[39],pp23[40],pp14[50],pp3[62]};
    CLA_4 KS_99(s99, c99, in99_1, in99_2);
    wire[3:0] s100, in100_1, in100_2;
    wire c100;
    assign in100_1 = {pp24[38],pp24[39],pp15[49],pp4[61]};
    assign in100_2 = {pp25[37],pp25[38],pp16[48],pp5[60]};
    CLA_4 KS_100(s100, c100, in100_1, in100_2);
    wire[3:0] s101, in101_1, in101_2;
    wire c101;
    assign in101_1 = {pp26[36],pp26[37],pp17[47],pp6[59]};
    assign in101_2 = {pp27[35],pp27[36],pp18[46],pp7[58]};
    CLA_4 KS_101(s101, c101, in101_1, in101_2);
    wire[3:0] s102, in102_1, in102_2;
    wire c102;
    assign in102_1 = {pp28[34],pp28[35],pp19[45],pp8[57]};
    assign in102_2 = {pp29[33],pp29[34],pp20[44],pp9[56]};
    CLA_4 KS_102(s102, c102, in102_1, in102_2);
    wire[3:0] s103, in103_1, in103_2;
    wire c103;
    assign in103_1 = {pp30[32],pp30[33],pp21[43],pp10[55]};
    assign in103_2 = {pp31[31],pp31[32],pp22[42],pp11[54]};
    CLA_4 KS_103(s103, c103, in103_1, in103_2);
    wire[3:0] s104, in104_1, in104_2;
    wire c104;
    assign in104_1 = {pp32[30],pp32[31],pp23[41],pp12[53]};
    assign in104_2 = {pp33[29],pp33[30],pp24[40],pp13[52]};
    CLA_4 KS_104(s104, c104, in104_1, in104_2);
    wire[3:0] s105, in105_1, in105_2;
    wire c105;
    assign in105_1 = {pp34[28],pp34[29],pp25[39],pp14[51]};
    assign in105_2 = {pp35[27],pp35[28],pp26[38],pp15[50]};
    CLA_4 KS_105(s105, c105, in105_1, in105_2);
    wire[3:0] s106, in106_1, in106_2;
    wire c106;
    assign in106_1 = {pp36[26],pp36[27],pp27[37],pp16[49]};
    assign in106_2 = {pp37[25],pp37[26],pp28[36],pp17[48]};
    CLA_4 KS_106(s106, c106, in106_1, in106_2);
    wire[3:0] s107, in107_1, in107_2;
    wire c107;
    assign in107_1 = {pp38[24],pp38[25],pp29[35],pp18[47]};
    assign in107_2 = {pp39[23],pp39[24],pp30[34],pp19[46]};
    CLA_4 KS_107(s107, c107, in107_1, in107_2);
    wire[3:0] s108, in108_1, in108_2;
    wire c108;
    assign in108_1 = {pp40[22],pp40[23],pp31[33],pp20[45]};
    assign in108_2 = {pp41[21],pp41[22],pp32[32],pp21[44]};
    CLA_4 KS_108(s108, c108, in108_1, in108_2);
    wire[3:0] s109, in109_1, in109_2;
    wire c109;
    assign in109_1 = {pp42[20],pp42[21],pp33[31],pp22[43]};
    assign in109_2 = {pp43[19],pp43[20],pp34[30],pp23[42]};
    CLA_4 KS_109(s109, c109, in109_1, in109_2);
    wire[3:0] s110, in110_1, in110_2;
    wire c110;
    assign in110_1 = {pp44[18],pp44[19],pp35[29],pp24[41]};
    assign in110_2 = {pp45[17],pp45[18],pp36[28],pp25[40]};
    CLA_4 KS_110(s110, c110, in110_1, in110_2);
    wire[3:0] s111, in111_1, in111_2;
    wire c111;
    assign in111_1 = {pp46[16],pp46[17],pp37[27],pp26[39]};
    assign in111_2 = {pp47[15],pp47[16],pp38[26],pp27[38]};
    CLA_4 KS_111(s111, c111, in111_1, in111_2);
    wire[3:0] s112, in112_1, in112_2;
    wire c112;
    assign in112_1 = {pp48[14],pp48[15],pp39[25],pp28[37]};
    assign in112_2 = {pp49[13],pp49[14],pp40[24],pp29[36]};
    CLA_4 KS_112(s112, c112, in112_1, in112_2);
    wire[3:0] s113, in113_1, in113_2;
    wire c113;
    assign in113_1 = {pp50[12],pp50[13],pp41[23],pp30[35]};
    assign in113_2 = {pp51[11],pp51[12],pp42[22],pp31[34]};
    CLA_4 KS_113(s113, c113, in113_1, in113_2);
    wire[3:0] s114, in114_1, in114_2;
    wire c114;
    assign in114_1 = {pp52[10],pp52[11],pp43[21],pp32[33]};
    assign in114_2 = {pp53[9],pp53[10],pp44[20],pp33[32]};
    CLA_4 KS_114(s114, c114, in114_1, in114_2);
    wire[0:0] s115, in115_1, in115_2;
    wire c115;
    assign in115_1 = {pp54[8]};
    assign in115_2 = {pp55[7]};
    Half_Adder KS_115(s115, c115, in115_1, in115_2);
    wire[3:0] s116, in116_1, in116_2;
    wire c116;
    assign in116_1 = {pp56[6],pp54[9],pp45[19],pp34[31]};
    assign in116_2 = {pp57[5],pp55[8],pp46[18],pp35[30]};
    CLA_4 KS_116(s116, c116, in116_1, in116_2);
    wire[0:0] s117, in117_1, in117_2;
    wire c117;
    assign in117_1 = {pp58[4]};
    assign in117_2 = {pp59[3]};
    Half_Adder KS_117(s117, c117, in117_1, in117_2);
    wire[3:0] s118, in118_1, in118_2;
    wire c118;
    assign in118_1 = {pp60[2],pp56[7],pp47[17],pp36[29]};
    assign in118_2 = {pp61[1],pp57[6],pp48[16],pp37[28]};
    CLA_4 KS_118(s118, c118, in118_1, in118_2);
    wire[0:0] s119, in119_1, in119_2;
    wire c119;
    assign in119_1 = {pp62[0]};
    assign in119_2 = {c67};
    Half_Adder KS_119(s119, c119, in119_1, in119_2);
    wire[3:0] s120, in120_1, in120_2;
    wire c120;
    assign in120_1 = {c68,pp58[5],pp49[15],pp38[27]};
    assign in120_2 = {c69,pp59[4],pp50[14],pp39[26]};
    CLA_4 KS_120(s120, c120, in120_1, in120_2);
    wire[0:0] s121, in121_1, in121_2;
    wire c121;
    assign in121_1 = {c70};
    assign in121_2 = {c71};
    Half_Adder KS_121(s121, c121, in121_1, in121_2);
    wire[3:0] s122, in122_1, in122_2;
    wire c122;
    assign in122_1 = {c72,pp60[3],pp51[13],pp40[25]};
    assign in122_2 = {c73,pp61[2],pp52[12],pp41[24]};
    CLA_4 KS_122(s122, c122, in122_1, in122_2);
    wire[0:0] s123, in123_1, in123_2;
    wire c123;
    assign in123_1 = {c74};
    assign in123_2 = {c75};
    Half_Adder KS_123(s123, c123, in123_1, in123_2);
    wire[3:0] s124, in124_1, in124_2;
    wire c124;
    assign in124_1 = {c76,pp62[1],pp53[11],pp42[23]};
    assign in124_2 = {c77,pp63[0],pp54[10],pp43[22]};
    CLA_4 KS_124(s124, c124, in124_1, in124_2);
    wire[0:0] s125, in125_1, in125_2;
    wire c125;
    assign in125_1 = {c78};
    assign in125_2 = {c79};
    Half_Adder KS_125(s125, c125, in125_1, in125_2);
    wire[3:0] s126, in126_1, in126_2;
    wire c126;
    assign in126_1 = {c80,s88[3],pp55[9],pp44[21]};
    assign in126_2 = {c82,s89[3],pp56[8],pp45[20]};
    CLA_4 KS_126(s126, c126, in126_1, in126_2);
    wire[0:0] s127, in127_1, in127_2;
    wire c127;
    assign in127_1 = {c84};
    assign in127_2 = {c86};
    Half_Adder KS_127(s127, c127, in127_1, in127_2);
    wire[3:0] s128, in128_1, in128_2;
    wire c128;
    assign in128_1 = {s89[2],s90[3],pp57[7],pp46[19]};
    assign in128_2 = {s90[2],s91[3],pp58[6],pp47[18]};
    CLA_4_c KS_128(s128, c128, in128_1, in128_2, s88[2]);
    wire[3:0] s129, in129_1, in129_2;
    wire c129;
    assign in129_1 = {pp60[4],pp48[17],pp3[63],pp4[63]};
    assign in129_2 = {pp61[3],pp49[16],pp4[62],pp5[62]};
    CLA_4_c KS_129(s129, c129, in129_1, in129_2, pp59[5]);
    wire[3:0] s130, in130_1, in130_2;
    wire c130;
    assign in130_1 = {pp50[15],pp5[61],pp6[61],pp5[63]};
    assign in130_2 = {pp51[14],pp6[60],pp7[60],pp6[62]};
    CLA_4 KS_130(s130, c130, in130_1, in130_2);
    wire[3:0] s131, in131_1, in131_2;
    wire c131;
    assign in131_1 = {pp52[13],pp7[59],pp8[59],pp7[61]};
    assign in131_2 = {pp53[12],pp8[58],pp9[58],pp8[60]};
    CLA_4 KS_131(s131, c131, in131_1, in131_2);
    wire[3:0] s132, in132_1, in132_2;
    wire c132;
    assign in132_1 = {pp54[11],pp9[57],pp10[57],pp9[59]};
    assign in132_2 = {pp55[10],pp10[56],pp11[56],pp10[58]};
    CLA_4 KS_132(s132, c132, in132_1, in132_2);
    wire[3:0] s133, in133_1, in133_2;
    wire c133;
    assign in133_1 = {pp56[9],pp11[55],pp12[55],pp11[57]};
    assign in133_2 = {pp57[8],pp12[54],pp13[54],pp12[56]};
    CLA_4 KS_133(s133, c133, in133_1, in133_2);
    wire[3:0] s134, in134_1, in134_2;
    wire c134;
    assign in134_1 = {pp59[6],pp13[53],pp14[53],pp13[55]};
    assign in134_2 = {pp60[5],pp14[52],pp15[52],pp14[54]};
    CLA_4_c KS_134(s134, c134, in134_1, in134_2, pp58[7]);
    wire[3:0] s135, in135_1, in135_2;
    wire c135;
    assign in135_1 = {pp15[51],pp16[51],pp15[53],pp6[63]};
    assign in135_2 = {pp16[50],pp17[50],pp16[52],pp7[62]};
    CLA_4 KS_135(s135, c135, in135_1, in135_2);
    wire[3:0] s136, in136_1, in136_2;
    wire c136;
    assign in136_1 = {pp17[49],pp18[49],pp17[51],pp8[61]};
    assign in136_2 = {pp18[48],pp19[48],pp18[50],pp9[60]};
    CLA_4 KS_136(s136, c136, in136_1, in136_2);
    wire[3:0] s137, in137_1, in137_2;
    wire c137;
    assign in137_1 = {pp19[47],pp20[47],pp19[49],pp10[59]};
    assign in137_2 = {pp20[46],pp21[46],pp20[48],pp11[58]};
    CLA_4 KS_137(s137, c137, in137_1, in137_2);
    wire[3:0] s138, in138_1, in138_2;
    wire c138;
    assign in138_1 = {pp21[45],pp22[45],pp21[47],pp12[57]};
    assign in138_2 = {pp22[44],pp23[44],pp22[46],pp13[56]};
    CLA_4 KS_138(s138, c138, in138_1, in138_2);
    wire[3:0] s139, in139_1, in139_2;
    wire c139;
    assign in139_1 = {pp23[43],pp24[43],pp23[45],pp14[55]};
    assign in139_2 = {pp24[42],pp25[42],pp24[44],pp15[54]};
    CLA_4 KS_139(s139, c139, in139_1, in139_2);
    wire[3:0] s140, in140_1, in140_2;
    wire c140;
    assign in140_1 = {pp25[41],pp26[41],pp25[43],pp16[53]};
    assign in140_2 = {pp26[40],pp27[40],pp26[42],pp17[52]};
    CLA_4 KS_140(s140, c140, in140_1, in140_2);
    wire[3:0] s141, in141_1, in141_2;
    wire c141;
    assign in141_1 = {pp27[39],pp28[39],pp27[41],pp18[51]};
    assign in141_2 = {pp28[38],pp29[38],pp28[40],pp19[50]};
    CLA_4 KS_141(s141, c141, in141_1, in141_2);
    wire[3:0] s142, in142_1, in142_2;
    wire c142;
    assign in142_1 = {pp29[37],pp30[37],pp29[39],pp20[49]};
    assign in142_2 = {pp30[36],pp31[36],pp30[38],pp21[48]};
    CLA_4 KS_142(s142, c142, in142_1, in142_2);
    wire[3:0] s143, in143_1, in143_2;
    wire c143;
    assign in143_1 = {pp31[35],pp32[35],pp31[37],pp22[47]};
    assign in143_2 = {pp32[34],pp33[34],pp32[36],pp23[46]};
    CLA_4 KS_143(s143, c143, in143_1, in143_2);
    wire[3:0] s144, in144_1, in144_2;
    wire c144;
    assign in144_1 = {pp33[33],pp34[33],pp33[35],pp24[45]};
    assign in144_2 = {pp34[32],pp35[32],pp34[34],pp25[44]};
    CLA_4 KS_144(s144, c144, in144_1, in144_2);
    wire[3:0] s145, in145_1, in145_2;
    wire c145;
    assign in145_1 = {pp35[31],pp36[31],pp35[33],pp26[43]};
    assign in145_2 = {pp36[30],pp37[30],pp36[32],pp27[42]};
    CLA_4 KS_145(s145, c145, in145_1, in145_2);
    wire[3:0] s146, in146_1, in146_2;
    wire c146;
    assign in146_1 = {pp37[29],pp38[29],pp37[31],pp28[41]};
    assign in146_2 = {pp38[28],pp39[28],pp38[30],pp29[40]};
    CLA_4 KS_146(s146, c146, in146_1, in146_2);
    wire[3:0] s147, in147_1, in147_2;
    wire c147;
    assign in147_1 = {pp39[27],pp40[27],pp39[29],pp30[39]};
    assign in147_2 = {pp40[26],pp41[26],pp40[28],pp31[38]};
    CLA_4 KS_147(s147, c147, in147_1, in147_2);
    wire[3:0] s148, in148_1, in148_2;
    wire c148;
    assign in148_1 = {pp41[25],pp42[25],pp41[27],pp32[37]};
    assign in148_2 = {pp42[24],pp43[24],pp42[26],pp33[36]};
    CLA_4 KS_148(s148, c148, in148_1, in148_2);
    wire[3:0] s149, in149_1, in149_2;
    wire c149;
    assign in149_1 = {pp43[23],pp44[23],pp43[25],pp34[35]};
    assign in149_2 = {pp44[22],pp45[22],pp44[24],pp35[34]};
    CLA_4 KS_149(s149, c149, in149_1, in149_2);
    wire[3:0] s150, in150_1, in150_2;
    wire c150;
    assign in150_1 = {pp45[21],pp46[21],pp45[23],pp36[33]};
    assign in150_2 = {pp46[20],pp47[20],pp46[22],pp37[32]};
    CLA_4 KS_150(s150, c150, in150_1, in150_2);
    wire[3:0] s151, in151_1, in151_2;
    wire c151;
    assign in151_1 = {pp47[19],pp48[19],pp47[21],pp38[31]};
    assign in151_2 = {pp48[18],pp49[18],pp48[20],pp39[30]};
    CLA_4 KS_151(s151, c151, in151_1, in151_2);
    wire[0:0] s152, in152_1, in152_2;
    wire c152;
    assign in152_1 = {pp49[17]};
    assign in152_2 = {pp50[16]};
    Half_Adder KS_152(s152, c152, in152_1, in152_2);
    wire[3:0] s153, in153_1, in153_2;
    wire c153;
    assign in153_1 = {pp51[15],pp50[17],pp49[19],pp40[29]};
    assign in153_2 = {pp52[14],pp51[16],pp50[18],pp41[28]};
    CLA_4 KS_153(s153, c153, in153_1, in153_2);
    wire[0:0] s154, in154_1, in154_2;
    wire c154;
    assign in154_1 = {pp53[13]};
    assign in154_2 = {pp54[12]};
    Half_Adder KS_154(s154, c154, in154_1, in154_2);
    wire[1:0] s155, in155_1, in155_2;
    wire c155;
    assign in155_1 = {pp55[11],pp52[15]};
    assign in155_2 = {pp56[10],pp53[14]};
    CLA_2 KS_155(s155, c155, in155_1, in155_2);
    wire[0:0] s156, in156_1, in156_2;
    wire c156;
    assign in156_1 = {pp57[9]};
    assign in156_2 = {pp58[8]};
    Half_Adder KS_156(s156, c156, in156_1, in156_2);
    wire[3:0] s157, in157_1, in157_2;
    wire c157;
    assign in157_1 = {pp59[7],pp54[13],pp51[17],pp42[27]};
    assign in157_2 = {pp60[6],pp55[12],pp52[16],pp43[26]};
    CLA_4 KS_157(s157, c157, in157_1, in157_2);
    wire[0:0] s158, in158_1, in158_2;
    wire c158;
    assign in158_1 = {pp61[5]};
    assign in158_2 = {pp62[4]};
    Half_Adder KS_158(s158, c158, in158_1, in158_2);
    wire[1:0] s159, in159_1, in159_2;
    wire c159;
    assign in159_1 = {pp63[3],pp56[11]};
    assign in159_2 = {c99,pp57[10]};
    CLA_2 KS_159(s159, c159, in159_1, in159_2);
    wire[0:0] s160, in160_1, in160_2;
    wire c160;
    assign in160_1 = {c100};
    assign in160_2 = {c101};
    Half_Adder KS_160(s160, c160, in160_1, in160_2);
    wire[3:0] s161, in161_1, in161_2;
    wire c161;
    assign in161_1 = {c102,pp58[9],pp53[15],pp44[25]};
    assign in161_2 = {c103,pp59[8],pp54[14],pp45[24]};
    CLA_4 KS_161(s161, c161, in161_1, in161_2);
    wire[0:0] s162, in162_1, in162_2;
    wire c162;
    assign in162_1 = {c104};
    assign in162_2 = {c105};
    Half_Adder KS_162(s162, c162, in162_1, in162_2);
    wire[1:0] s163, in163_1, in163_2;
    wire c163;
    assign in163_1 = {c106,pp60[7]};
    assign in163_2 = {c107,pp61[6]};
    CLA_2 KS_163(s163, c163, in163_1, in163_2);
    wire[0:0] s164, in164_1, in164_2;
    wire c164;
    assign in164_1 = {c108};
    assign in164_2 = {c109};
    Half_Adder KS_164(s164, c164, in164_1, in164_2);
    wire[3:0] s165, in165_1, in165_2;
    wire c165;
    assign in165_1 = {c110,pp62[5],pp55[13],pp46[23]};
    assign in165_2 = {c111,pp63[4],pp56[12],pp47[22]};
    CLA_4 KS_165(s165, c165, in165_1, in165_2);
    wire[0:0] s166, in166_1, in166_2;
    wire c166;
    assign in166_1 = {c112};
    assign in166_2 = {c113};
    Half_Adder KS_166(s166, c166, in166_1, in166_2);
    wire[1:0] s167, in167_1, in167_2;
    wire c167;
    assign in167_1 = {c114,s129[3]};
    assign in167_2 = {c116,s130[2]};
    CLA_2 KS_167(s167, c167, in167_1, in167_2);
    wire[0:0] s168, in168_1, in168_2;
    wire c168;
    assign in168_1 = {c118};
    assign in168_2 = {c120};
    Half_Adder KS_168(s168, c168, in168_1, in168_2);
    wire[3:0] s169, in169_1, in169_2;
    wire c169;
    assign in169_1 = {c122,s131[2],pp57[11],pp48[21]};
    assign in169_2 = {c124,s132[2],pp58[10],pp49[20]};
    CLA_4 KS_169(s169, c169, in169_1, in169_2);
    wire[0:0] s170, in170_1, in170_2;
    wire c170;
    assign in170_1 = {c126};
    assign in170_2 = {c128};
    Half_Adder KS_170(s170, c170, in170_1, in170_2);
    wire[1:0] s171, in171_1, in171_2;
    wire c171;
    assign in171_1 = {s129[2],s133[2]};
    assign in171_2 = {s130[1],s134[2]};
    CLA_2 KS_171(s171, c171, in171_1, in171_2);
    wire[0:0] s172, in172_1, in172_2;
    wire c172;
    assign in172_1 = {s131[1]};
    assign in172_2 = {s132[1]};
    Half_Adder KS_172(s172, c172, in172_1, in172_2);
    wire[3:0] s173, in173_1, in173_2;
    wire c173;
    assign in173_1 = {s134[1],s135[1],pp59[9],pp50[19]};
    assign in173_2 = {s135[0],s136[1],pp60[8],pp51[18]};
    CLA_4_c KS_173(s173, c173, in173_1, in173_2, s133[1]);
    wire[3:0] s174, in174_1, in174_2;
    wire c174;
    assign in174_1 = {pp53[16],pp7[63],pp8[63],pp9[63]};
    assign in174_2 = {pp54[15],pp8[62],pp9[62],pp10[62]};
    CLA_4_c KS_174(s174, c174, in174_1, in174_2, pp52[17]);
    wire[3:0] s175, in175_1, in175_2;
    wire c175;
    assign in175_1 = {pp9[61],pp10[61],pp11[61],pp10[63]};
    assign in175_2 = {pp10[60],pp11[60],pp12[60],pp11[62]};
    CLA_4 KS_175(s175, c175, in175_1, in175_2);
    wire[3:0] s176, in176_1, in176_2;
    wire c176;
    assign in176_1 = {pp11[59],pp12[59],pp13[59],pp12[61]};
    assign in176_2 = {pp12[58],pp13[58],pp14[58],pp13[60]};
    CLA_4 KS_176(s176, c176, in176_1, in176_2);
    wire[3:0] s177, in177_1, in177_2;
    wire c177;
    assign in177_1 = {pp13[57],pp14[57],pp15[57],pp14[59]};
    assign in177_2 = {pp14[56],pp15[56],pp16[56],pp15[58]};
    CLA_4 KS_177(s177, c177, in177_1, in177_2);
    wire[3:0] s178, in178_1, in178_2;
    wire c178;
    assign in178_1 = {pp15[55],pp16[55],pp17[55],pp16[57]};
    assign in178_2 = {pp16[54],pp17[54],pp18[54],pp17[56]};
    CLA_4 KS_178(s178, c178, in178_1, in178_2);
    wire[3:0] s179, in179_1, in179_2;
    wire c179;
    assign in179_1 = {pp17[53],pp18[53],pp19[53],pp18[55]};
    assign in179_2 = {pp18[52],pp19[52],pp20[52],pp19[54]};
    CLA_4 KS_179(s179, c179, in179_1, in179_2);
    wire[3:0] s180, in180_1, in180_2;
    wire c180;
    assign in180_1 = {pp19[51],pp20[51],pp21[51],pp20[53]};
    assign in180_2 = {pp20[50],pp21[50],pp22[50],pp21[52]};
    CLA_4 KS_180(s180, c180, in180_1, in180_2);
    wire[3:0] s181, in181_1, in181_2;
    wire c181;
    assign in181_1 = {pp21[49],pp22[49],pp23[49],pp22[51]};
    assign in181_2 = {pp22[48],pp23[48],pp24[48],pp23[50]};
    CLA_4 KS_181(s181, c181, in181_1, in181_2);
    wire[3:0] s182, in182_1, in182_2;
    wire c182;
    assign in182_1 = {pp23[47],pp24[47],pp25[47],pp24[49]};
    assign in182_2 = {pp24[46],pp25[46],pp26[46],pp25[48]};
    CLA_4 KS_182(s182, c182, in182_1, in182_2);
    wire[3:0] s183, in183_1, in183_2;
    wire c183;
    assign in183_1 = {pp25[45],pp26[45],pp27[45],pp26[47]};
    assign in183_2 = {pp26[44],pp27[44],pp28[44],pp27[46]};
    CLA_4 KS_183(s183, c183, in183_1, in183_2);
    wire[3:0] s184, in184_1, in184_2;
    wire c184;
    assign in184_1 = {pp27[43],pp28[43],pp29[43],pp28[45]};
    assign in184_2 = {pp28[42],pp29[42],pp30[42],pp29[44]};
    CLA_4 KS_184(s184, c184, in184_1, in184_2);
    wire[3:0] s185, in185_1, in185_2;
    wire c185;
    assign in185_1 = {pp29[41],pp30[41],pp31[41],pp30[43]};
    assign in185_2 = {pp30[40],pp31[40],pp32[40],pp31[42]};
    CLA_4 KS_185(s185, c185, in185_1, in185_2);
    wire[3:0] s186, in186_1, in186_2;
    wire c186;
    assign in186_1 = {pp31[39],pp32[39],pp33[39],pp32[41]};
    assign in186_2 = {pp32[38],pp33[38],pp34[38],pp33[40]};
    CLA_4 KS_186(s186, c186, in186_1, in186_2);
    wire[3:0] s187, in187_1, in187_2;
    wire c187;
    assign in187_1 = {pp33[37],pp34[37],pp35[37],pp34[39]};
    assign in187_2 = {pp34[36],pp35[36],pp36[36],pp35[38]};
    CLA_4 KS_187(s187, c187, in187_1, in187_2);
    wire[3:0] s188, in188_1, in188_2;
    wire c188;
    assign in188_1 = {pp35[35],pp36[35],pp37[35],pp36[37]};
    assign in188_2 = {pp36[34],pp37[34],pp38[34],pp37[36]};
    CLA_4 KS_188(s188, c188, in188_1, in188_2);
    wire[3:0] s189, in189_1, in189_2;
    wire c189;
    assign in189_1 = {pp37[33],pp38[33],pp39[33],pp38[35]};
    assign in189_2 = {pp38[32],pp39[32],pp40[32],pp39[34]};
    CLA_4 KS_189(s189, c189, in189_1, in189_2);
    wire[3:0] s190, in190_1, in190_2;
    wire c190;
    assign in190_1 = {pp39[31],pp40[31],pp41[31],pp40[33]};
    assign in190_2 = {pp40[30],pp41[30],pp42[30],pp41[32]};
    CLA_4 KS_190(s190, c190, in190_1, in190_2);
    wire[3:0] s191, in191_1, in191_2;
    wire c191;
    assign in191_1 = {pp41[29],pp42[29],pp43[29],pp42[31]};
    assign in191_2 = {pp42[28],pp43[28],pp44[28],pp43[30]};
    CLA_4 KS_191(s191, c191, in191_1, in191_2);
    wire[1:0] s192, in192_1, in192_2;
    wire c192;
    assign in192_1 = {pp43[27],pp44[27]};
    assign in192_2 = {pp44[26],pp45[26]};
    CLA_2 KS_192(s192, c192, in192_1, in192_2);
    wire[0:0] s193, in193_1, in193_2;
    wire c193;
    assign in193_1 = {pp45[25]};
    assign in193_2 = {pp46[24]};
    Half_Adder KS_193(s193, c193, in193_1, in193_2);
    wire[3:0] s194, in194_1, in194_2;
    wire c194;
    assign in194_1 = {pp47[23],pp46[25],pp45[27],pp44[29]};
    assign in194_2 = {pp48[22],pp47[24],pp46[26],pp45[28]};
    CLA_4 KS_194(s194, c194, in194_1, in194_2);
    wire[0:0] s195, in195_1, in195_2;
    wire c195;
    assign in195_1 = {pp49[21]};
    assign in195_2 = {pp50[20]};
    Half_Adder KS_195(s195, c195, in195_1, in195_2);
    wire[1:0] s196, in196_1, in196_2;
    wire c196;
    assign in196_1 = {pp51[19],pp48[23]};
    assign in196_2 = {pp52[18],pp49[22]};
    CLA_2 KS_196(s196, c196, in196_1, in196_2);
    wire[0:0] s197, in197_1, in197_2;
    wire c197;
    assign in197_1 = {pp53[17]};
    assign in197_2 = {pp54[16]};
    Half_Adder KS_197(s197, c197, in197_1, in197_2);
    wire[2:0] s198, in198_1, in198_2;
    wire c198;
    assign in198_1 = {pp55[15],pp50[21],pp47[25]};
    assign in198_2 = {pp56[14],pp51[20],pp48[24]};
    CLA_3 KS_198(s198, c198, in198_1, in198_2);
    wire[0:0] s199, in199_1, in199_2;
    wire c199;
    assign in199_1 = {pp57[13]};
    assign in199_2 = {pp58[12]};
    Half_Adder KS_199(s199, c199, in199_1, in199_2);
    wire[1:0] s200, in200_1, in200_2;
    wire c200;
    assign in200_1 = {pp59[11],pp52[19]};
    assign in200_2 = {pp60[10],pp53[18]};
    CLA_2 KS_200(s200, c200, in200_1, in200_2);
    wire[0:0] s201, in201_1, in201_2;
    wire c201;
    assign in201_1 = {pp61[9]};
    assign in201_2 = {pp62[8]};
    Half_Adder KS_201(s201, c201, in201_1, in201_2);
    wire[3:0] s202, in202_1, in202_2;
    wire c202;
    assign in202_1 = {pp63[7],pp54[17],pp49[23],pp46[27]};
    assign in202_2 = {c135,pp55[16],pp50[22],pp47[26]};
    CLA_4 KS_202(s202, c202, in202_1, in202_2);
    wire[0:0] s203, in203_1, in203_2;
    wire c203;
    assign in203_1 = {c136};
    assign in203_2 = {c137};
    Half_Adder KS_203(s203, c203, in203_1, in203_2);
    wire[1:0] s204, in204_1, in204_2;
    wire c204;
    assign in204_1 = {c138,pp56[15]};
    assign in204_2 = {c139,pp57[14]};
    CLA_2 KS_204(s204, c204, in204_1, in204_2);
    wire[0:0] s205, in205_1, in205_2;
    wire c205;
    assign in205_1 = {c140};
    assign in205_2 = {c141};
    Half_Adder KS_205(s205, c205, in205_1, in205_2);
    wire[2:0] s206, in206_1, in206_2;
    wire c206;
    assign in206_1 = {c142,pp58[13],pp51[21]};
    assign in206_2 = {c143,pp59[12],pp52[20]};
    CLA_3 KS_206(s206, c206, in206_1, in206_2);
    wire[0:0] s207, in207_1, in207_2;
    wire c207;
    assign in207_1 = {c144};
    assign in207_2 = {c145};
    Half_Adder KS_207(s207, c207, in207_1, in207_2);
    wire[1:0] s208, in208_1, in208_2;
    wire c208;
    assign in208_1 = {c146,pp60[11]};
    assign in208_2 = {c147,pp61[10]};
    CLA_2 KS_208(s208, c208, in208_1, in208_2);
    wire[0:0] s209, in209_1, in209_2;
    wire c209;
    assign in209_1 = {c148};
    assign in209_2 = {c149};
    Half_Adder KS_209(s209, c209, in209_1, in209_2);
    wire[3:0] s210, in210_1, in210_2;
    wire c210;
    assign in210_1 = {c150,pp62[9],pp53[19],pp48[25]};
    assign in210_2 = {c151,pp63[8],pp54[18],pp49[24]};
    CLA_4 KS_210(s210, c210, in210_1, in210_2);
    wire[0:0] s211, in211_1, in211_2;
    wire c211;
    assign in211_1 = {c153};
    assign in211_2 = {c157};
    Half_Adder KS_211(s211, c211, in211_1, in211_2);
    wire[1:0] s212, in212_1, in212_2;
    wire c212;
    assign in212_1 = {c161,s174[2]};
    assign in212_2 = {c165,s175[1]};
    CLA_2 KS_212(s212, c212, in212_1, in212_2);
    wire[0:0] s213, in213_1, in213_2;
    wire c213;
    assign in213_1 = {c169};
    assign in213_2 = {c173};
    Half_Adder KS_213(s213, c213, in213_1, in213_2);
    wire[2:0] s214, in214_1, in214_2;
    wire c214;
    assign in214_1 = {s175[0],s176[1],pp55[17]};
    assign in214_2 = {s176[0],s177[1],pp56[16]};
    CLA_3_c KS_214(s214, c214, in214_1, in214_2, s174[1]);
    wire[3:0] s215, in215_1, in215_2;
    wire c215;
    assign in215_1 = {pp11[63],pp12[63],pp13[63],pp14[63]};
    assign in215_2 = {pp12[62],pp13[62],pp14[62],pp15[62]};
    CLA_4 KS_215(s215, c215, in215_1, in215_2);
    wire[3:0] s216, in216_1, in216_2;
    wire c216;
    assign in216_1 = {pp13[61],pp14[61],pp15[61],pp16[61]};
    assign in216_2 = {pp14[60],pp15[60],pp16[60],pp17[60]};
    CLA_4 KS_216(s216, c216, in216_1, in216_2);
    wire[3:0] s217, in217_1, in217_2;
    wire c217;
    assign in217_1 = {pp15[59],pp16[59],pp17[59],pp18[59]};
    assign in217_2 = {pp16[58],pp17[58],pp18[58],pp19[58]};
    CLA_4 KS_217(s217, c217, in217_1, in217_2);
    wire[3:0] s218, in218_1, in218_2;
    wire c218;
    assign in218_1 = {pp17[57],pp18[57],pp19[57],pp20[57]};
    assign in218_2 = {pp18[56],pp19[56],pp20[56],pp21[56]};
    CLA_4 KS_218(s218, c218, in218_1, in218_2);
    wire[3:0] s219, in219_1, in219_2;
    wire c219;
    assign in219_1 = {pp19[55],pp20[55],pp21[55],pp22[55]};
    assign in219_2 = {pp20[54],pp21[54],pp22[54],pp23[54]};
    CLA_4 KS_219(s219, c219, in219_1, in219_2);
    wire[3:0] s220, in220_1, in220_2;
    wire c220;
    assign in220_1 = {pp21[53],pp22[53],pp23[53],pp24[53]};
    assign in220_2 = {pp22[52],pp23[52],pp24[52],pp25[52]};
    CLA_4 KS_220(s220, c220, in220_1, in220_2);
    wire[3:0] s221, in221_1, in221_2;
    wire c221;
    assign in221_1 = {pp23[51],pp24[51],pp25[51],pp26[51]};
    assign in221_2 = {pp24[50],pp25[50],pp26[50],pp27[50]};
    CLA_4 KS_221(s221, c221, in221_1, in221_2);
    wire[3:0] s222, in222_1, in222_2;
    wire c222;
    assign in222_1 = {pp25[49],pp26[49],pp27[49],pp28[49]};
    assign in222_2 = {pp26[48],pp27[48],pp28[48],pp29[48]};
    CLA_4 KS_222(s222, c222, in222_1, in222_2);
    wire[3:0] s223, in223_1, in223_2;
    wire c223;
    assign in223_1 = {pp27[47],pp28[47],pp29[47],pp30[47]};
    assign in223_2 = {pp28[46],pp29[46],pp30[46],pp31[46]};
    CLA_4 KS_223(s223, c223, in223_1, in223_2);
    wire[3:0] s224, in224_1, in224_2;
    wire c224;
    assign in224_1 = {pp29[45],pp30[45],pp31[45],pp32[45]};
    assign in224_2 = {pp30[44],pp31[44],pp32[44],pp33[44]};
    CLA_4 KS_224(s224, c224, in224_1, in224_2);
    wire[3:0] s225, in225_1, in225_2;
    wire c225;
    assign in225_1 = {pp31[43],pp32[43],pp33[43],pp34[43]};
    assign in225_2 = {pp32[42],pp33[42],pp34[42],pp35[42]};
    CLA_4 KS_225(s225, c225, in225_1, in225_2);
    wire[3:0] s226, in226_1, in226_2;
    wire c226;
    assign in226_1 = {pp33[41],pp34[41],pp35[41],pp36[41]};
    assign in226_2 = {pp34[40],pp35[40],pp36[40],pp37[40]};
    CLA_4 KS_226(s226, c226, in226_1, in226_2);
    wire[3:0] s227, in227_1, in227_2;
    wire c227;
    assign in227_1 = {pp35[39],pp36[39],pp37[39],pp38[39]};
    assign in227_2 = {pp36[38],pp37[38],pp38[38],pp39[38]};
    CLA_4 KS_227(s227, c227, in227_1, in227_2);
    wire[2:0] s228, in228_1, in228_2;
    wire c228;
    assign in228_1 = {pp37[37],pp38[37],pp39[37]};
    assign in228_2 = {pp38[36],pp39[36],pp40[36]};
    CLA_3 KS_228(s228, c228, in228_1, in228_2);
    wire[1:0] s229, in229_1, in229_2;
    wire c229;
    assign in229_1 = {pp39[35],pp40[35]};
    assign in229_2 = {pp40[34],pp41[34]};
    CLA_2 KS_229(s229, c229, in229_1, in229_2);
    wire[0:0] s230, in230_1, in230_2;
    wire c230;
    assign in230_1 = {pp41[33]};
    assign in230_2 = {pp42[32]};
    Half_Adder KS_230(s230, c230, in230_1, in230_2);
    wire[3:0] s231, in231_1, in231_2;
    wire c231;
    assign in231_1 = {pp43[31],pp42[33],pp41[35],pp40[37]};
    assign in231_2 = {pp44[30],pp43[32],pp42[34],pp41[36]};
    CLA_4 KS_231(s231, c231, in231_1, in231_2);
    wire[0:0] s232, in232_1, in232_2;
    wire c232;
    assign in232_1 = {pp45[29]};
    assign in232_2 = {pp46[28]};
    Half_Adder KS_232(s232, c232, in232_1, in232_2);
    wire[1:0] s233, in233_1, in233_2;
    wire c233;
    assign in233_1 = {pp47[27],pp44[31]};
    assign in233_2 = {pp48[26],pp45[30]};
    CLA_2 KS_233(s233, c233, in233_1, in233_2);
    wire[0:0] s234, in234_1, in234_2;
    wire c234;
    assign in234_1 = {pp49[25]};
    assign in234_2 = {pp50[24]};
    Half_Adder KS_234(s234, c234, in234_1, in234_2);
    wire[2:0] s235, in235_1, in235_2;
    wire c235;
    assign in235_1 = {pp51[23],pp46[29],pp43[33]};
    assign in235_2 = {pp52[22],pp47[28],pp44[32]};
    CLA_3 KS_235(s235, c235, in235_1, in235_2);
    wire[0:0] s236, in236_1, in236_2;
    wire c236;
    assign in236_1 = {pp53[21]};
    assign in236_2 = {pp54[20]};
    Half_Adder KS_236(s236, c236, in236_1, in236_2);
    wire[1:0] s237, in237_1, in237_2;
    wire c237;
    assign in237_1 = {pp55[19],pp48[27]};
    assign in237_2 = {pp56[18],pp49[26]};
    CLA_2 KS_237(s237, c237, in237_1, in237_2);
    wire[0:0] s238, in238_1, in238_2;
    wire c238;
    assign in238_1 = {pp57[17]};
    assign in238_2 = {pp58[16]};
    Half_Adder KS_238(s238, c238, in238_1, in238_2);
    wire[3:0] s239, in239_1, in239_2;
    wire c239;
    assign in239_1 = {pp59[15],pp50[25],pp45[31],pp42[35]};
    assign in239_2 = {pp60[14],pp51[24],pp46[30],pp43[34]};
    CLA_4 KS_239(s239, c239, in239_1, in239_2);
    wire[0:0] s240, in240_1, in240_2;
    wire c240;
    assign in240_1 = {pp61[13]};
    assign in240_2 = {pp62[12]};
    Half_Adder KS_240(s240, c240, in240_1, in240_2);
    wire[1:0] s241, in241_1, in241_2;
    wire c241;
    assign in241_1 = {pp63[11],pp52[23]};
    assign in241_2 = {c175,pp53[22]};
    CLA_2 KS_241(s241, c241, in241_1, in241_2);
    wire[0:0] s242, in242_1, in242_2;
    wire c242;
    assign in242_1 = {c176};
    assign in242_2 = {c177};
    Half_Adder KS_242(s242, c242, in242_1, in242_2);
    wire[2:0] s243, in243_1, in243_2;
    wire c243;
    assign in243_1 = {c178,pp54[21],pp47[29]};
    assign in243_2 = {c179,pp55[20],pp48[28]};
    CLA_3 KS_243(s243, c243, in243_1, in243_2);
    wire[0:0] s244, in244_1, in244_2;
    wire c244;
    assign in244_1 = {c180};
    assign in244_2 = {c181};
    Half_Adder KS_244(s244, c244, in244_1, in244_2);
    wire[1:0] s245, in245_1, in245_2;
    wire c245;
    assign in245_1 = {c182,pp56[19]};
    assign in245_2 = {c183,pp57[18]};
    CLA_2 KS_245(s245, c245, in245_1, in245_2);
    wire[0:0] s246, in246_1, in246_2;
    wire c246;
    assign in246_1 = {c184};
    assign in246_2 = {c185};
    Half_Adder KS_246(s246, c246, in246_1, in246_2);
    wire[3:0] s247, in247_1, in247_2;
    wire c247;
    assign in247_1 = {c186,pp58[17],pp49[27],pp44[33]};
    assign in247_2 = {c187,pp59[16],pp50[26],pp45[32]};
    CLA_4 KS_247(s247, c247, in247_1, in247_2);
    wire[0:0] s248, in248_1, in248_2;
    wire c248;
    assign in248_1 = {c189};
    assign in248_2 = {c190};
    Full_Adder KS_248(s248, c248, in248_1, in248_2, c188);
    wire[3:0] s249, in249_1, in249_2;
    wire c249;
    assign in249_1 = {pp15[63],pp16[63],pp17[63],pp18[63]};
    assign in249_2 = {pp16[62],pp17[62],pp18[62],pp19[62]};
    CLA_4 KS_249(s249, c249, in249_1, in249_2);
    wire[3:0] s250, in250_1, in250_2;
    wire c250;
    assign in250_1 = {pp17[61],pp18[61],pp19[61],pp20[61]};
    assign in250_2 = {pp18[60],pp19[60],pp20[60],pp21[60]};
    CLA_4 KS_250(s250, c250, in250_1, in250_2);
    wire[3:0] s251, in251_1, in251_2;
    wire c251;
    assign in251_1 = {pp19[59],pp20[59],pp21[59],pp22[59]};
    assign in251_2 = {pp20[58],pp21[58],pp22[58],pp23[58]};
    CLA_4 KS_251(s251, c251, in251_1, in251_2);
    wire[3:0] s252, in252_1, in252_2;
    wire c252;
    assign in252_1 = {pp21[57],pp22[57],pp23[57],pp24[57]};
    assign in252_2 = {pp22[56],pp23[56],pp24[56],pp25[56]};
    CLA_4 KS_252(s252, c252, in252_1, in252_2);
    wire[3:0] s253, in253_1, in253_2;
    wire c253;
    assign in253_1 = {pp23[55],pp24[55],pp25[55],pp26[55]};
    assign in253_2 = {pp24[54],pp25[54],pp26[54],pp27[54]};
    CLA_4 KS_253(s253, c253, in253_1, in253_2);
    wire[3:0] s254, in254_1, in254_2;
    wire c254;
    assign in254_1 = {pp25[53],pp26[53],pp27[53],pp28[53]};
    assign in254_2 = {pp26[52],pp27[52],pp28[52],pp29[52]};
    CLA_4 KS_254(s254, c254, in254_1, in254_2);
    wire[3:0] s255, in255_1, in255_2;
    wire c255;
    assign in255_1 = {pp27[51],pp28[51],pp29[51],pp30[51]};
    assign in255_2 = {pp28[50],pp29[50],pp30[50],pp31[50]};
    CLA_4 KS_255(s255, c255, in255_1, in255_2);
    wire[3:0] s256, in256_1, in256_2;
    wire c256;
    assign in256_1 = {pp29[49],pp30[49],pp31[49],pp32[49]};
    assign in256_2 = {pp30[48],pp31[48],pp32[48],pp33[48]};
    CLA_4 KS_256(s256, c256, in256_1, in256_2);
    wire[3:0] s257, in257_1, in257_2;
    wire c257;
    assign in257_1 = {pp31[47],pp32[47],pp33[47],pp34[47]};
    assign in257_2 = {pp32[46],pp33[46],pp34[46],pp35[46]};
    CLA_4 KS_257(s257, c257, in257_1, in257_2);
    wire[2:0] s258, in258_1, in258_2;
    wire c258;
    assign in258_1 = {pp33[45],pp34[45],pp35[45]};
    assign in258_2 = {pp34[44],pp35[44],pp36[44]};
    CLA_3 KS_258(s258, c258, in258_1, in258_2);
    wire[1:0] s259, in259_1, in259_2;
    wire c259;
    assign in259_1 = {pp35[43],pp36[43]};
    assign in259_2 = {pp36[42],pp37[42]};
    CLA_2 KS_259(s259, c259, in259_1, in259_2);
    wire[0:0] s260, in260_1, in260_2;
    wire c260;
    assign in260_1 = {pp37[41]};
    assign in260_2 = {pp38[40]};
    Half_Adder KS_260(s260, c260, in260_1, in260_2);
    wire[3:0] s261, in261_1, in261_2;
    wire c261;
    assign in261_1 = {pp39[39],pp38[41],pp37[43],pp36[45]};
    assign in261_2 = {pp40[38],pp39[40],pp38[42],pp37[44]};
    CLA_4 KS_261(s261, c261, in261_1, in261_2);
    wire[0:0] s262, in262_1, in262_2;
    wire c262;
    assign in262_1 = {pp41[37]};
    assign in262_2 = {pp42[36]};
    Half_Adder KS_262(s262, c262, in262_1, in262_2);
    wire[1:0] s263, in263_1, in263_2;
    wire c263;
    assign in263_1 = {pp43[35],pp40[39]};
    assign in263_2 = {pp44[34],pp41[38]};
    CLA_2 KS_263(s263, c263, in263_1, in263_2);
    wire[0:0] s264, in264_1, in264_2;
    wire c264;
    assign in264_1 = {pp45[33]};
    assign in264_2 = {pp46[32]};
    Half_Adder KS_264(s264, c264, in264_1, in264_2);
    wire[2:0] s265, in265_1, in265_2;
    wire c265;
    assign in265_1 = {pp47[31],pp42[37],pp39[41]};
    assign in265_2 = {pp48[30],pp43[36],pp40[40]};
    CLA_3 KS_265(s265, c265, in265_1, in265_2);
    wire[0:0] s266, in266_1, in266_2;
    wire c266;
    assign in266_1 = {pp49[29]};
    assign in266_2 = {pp50[28]};
    Half_Adder KS_266(s266, c266, in266_1, in266_2);
    wire[1:0] s267, in267_1, in267_2;
    wire c267;
    assign in267_1 = {pp51[27],pp44[35]};
    assign in267_2 = {pp52[26],pp45[34]};
    CLA_2 KS_267(s267, c267, in267_1, in267_2);
    wire[0:0] s268, in268_1, in268_2;
    wire c268;
    assign in268_1 = {pp53[25]};
    assign in268_2 = {pp54[24]};
    Half_Adder KS_268(s268, c268, in268_1, in268_2);
    wire[3:0] s269, in269_1, in269_2;
    wire c269;
    assign in269_1 = {pp55[23],pp46[33],pp41[39],pp38[43]};
    assign in269_2 = {pp56[22],pp47[32],pp42[38],pp39[42]};
    CLA_4 KS_269(s269, c269, in269_1, in269_2);
    wire[0:0] s270, in270_1, in270_2;
    wire c270;
    assign in270_1 = {pp57[21]};
    assign in270_2 = {pp58[20]};
    Half_Adder KS_270(s270, c270, in270_1, in270_2);
    wire[1:0] s271, in271_1, in271_2;
    wire c271;
    assign in271_1 = {pp59[19],pp48[31]};
    assign in271_2 = {pp60[18],pp49[30]};
    CLA_2 KS_271(s271, c271, in271_1, in271_2);
    wire[0:0] s272, in272_1, in272_2;
    wire c272;
    assign in272_1 = {pp61[17]};
    assign in272_2 = {pp62[16]};
    Half_Adder KS_272(s272, c272, in272_1, in272_2);
    wire[2:0] s273, in273_1, in273_2;
    wire c273;
    assign in273_1 = {pp63[15],pp50[29],pp43[37]};
    assign in273_2 = {c215,pp51[28],pp44[36]};
    CLA_3 KS_273(s273, c273, in273_1, in273_2);
    wire[0:0] s274, in274_1, in274_2;
    wire c274;
    assign in274_1 = {c217};
    assign in274_2 = {c218};
    Full_Adder KS_274(s274, c274, in274_1, in274_2, c216);
    wire[3:0] s275, in275_1, in275_2;
    wire c275;
    assign in275_1 = {pp19[63],pp20[63],pp21[63],pp22[63]};
    assign in275_2 = {pp20[62],pp21[62],pp22[62],pp23[62]};
    CLA_4 KS_275(s275, c275, in275_1, in275_2);
    wire[3:0] s276, in276_1, in276_2;
    wire c276;
    assign in276_1 = {pp21[61],pp22[61],pp23[61],pp24[61]};
    assign in276_2 = {pp22[60],pp23[60],pp24[60],pp25[60]};
    CLA_4 KS_276(s276, c276, in276_1, in276_2);
    wire[3:0] s277, in277_1, in277_2;
    wire c277;
    assign in277_1 = {pp23[59],pp24[59],pp25[59],pp26[59]};
    assign in277_2 = {pp24[58],pp25[58],pp26[58],pp27[58]};
    CLA_4 KS_277(s277, c277, in277_1, in277_2);
    wire[3:0] s278, in278_1, in278_2;
    wire c278;
    assign in278_1 = {pp25[57],pp26[57],pp27[57],pp28[57]};
    assign in278_2 = {pp26[56],pp27[56],pp28[56],pp29[56]};
    CLA_4 KS_278(s278, c278, in278_1, in278_2);
    wire[3:0] s279, in279_1, in279_2;
    wire c279;
    assign in279_1 = {pp27[55],pp28[55],pp29[55],pp30[55]};
    assign in279_2 = {pp28[54],pp29[54],pp30[54],pp31[54]};
    CLA_4 KS_279(s279, c279, in279_1, in279_2);
    wire[2:0] s280, in280_1, in280_2;
    wire c280;
    assign in280_1 = {pp29[53],pp30[53],pp31[53]};
    assign in280_2 = {pp30[52],pp31[52],pp32[52]};
    CLA_3 KS_280(s280, c280, in280_1, in280_2);
    wire[1:0] s281, in281_1, in281_2;
    wire c281;
    assign in281_1 = {pp31[51],pp32[51]};
    assign in281_2 = {pp32[50],pp33[50]};
    CLA_2 KS_281(s281, c281, in281_1, in281_2);
    wire[0:0] s282, in282_1, in282_2;
    wire c282;
    assign in282_1 = {pp33[49]};
    assign in282_2 = {pp34[48]};
    Half_Adder KS_282(s282, c282, in282_1, in282_2);
    wire[3:0] s283, in283_1, in283_2;
    wire c283;
    assign in283_1 = {pp35[47],pp34[49],pp33[51],pp32[53]};
    assign in283_2 = {pp36[46],pp35[48],pp34[50],pp33[52]};
    CLA_4 KS_283(s283, c283, in283_1, in283_2);
    wire[0:0] s284, in284_1, in284_2;
    wire c284;
    assign in284_1 = {pp37[45]};
    assign in284_2 = {pp38[44]};
    Half_Adder KS_284(s284, c284, in284_1, in284_2);
    wire[1:0] s285, in285_1, in285_2;
    wire c285;
    assign in285_1 = {pp39[43],pp36[47]};
    assign in285_2 = {pp40[42],pp37[46]};
    CLA_2 KS_285(s285, c285, in285_1, in285_2);
    wire[0:0] s286, in286_1, in286_2;
    wire c286;
    assign in286_1 = {pp41[41]};
    assign in286_2 = {pp42[40]};
    Half_Adder KS_286(s286, c286, in286_1, in286_2);
    wire[2:0] s287, in287_1, in287_2;
    wire c287;
    assign in287_1 = {pp43[39],pp38[45],pp35[49]};
    assign in287_2 = {pp44[38],pp39[44],pp36[48]};
    CLA_3 KS_287(s287, c287, in287_1, in287_2);
    wire[0:0] s288, in288_1, in288_2;
    wire c288;
    assign in288_1 = {pp45[37]};
    assign in288_2 = {pp46[36]};
    Half_Adder KS_288(s288, c288, in288_1, in288_2);
    wire[1:0] s289, in289_1, in289_2;
    wire c289;
    assign in289_1 = {pp47[35],pp40[43]};
    assign in289_2 = {pp48[34],pp41[42]};
    CLA_2 KS_289(s289, c289, in289_1, in289_2);
    wire[0:0] s290, in290_1, in290_2;
    wire c290;
    assign in290_1 = {pp49[33]};
    assign in290_2 = {pp50[32]};
    Half_Adder KS_290(s290, c290, in290_1, in290_2);
    wire[3:0] s291, in291_1, in291_2;
    wire c291;
    assign in291_1 = {pp52[30],pp42[41],pp37[47],pp34[51]};
    assign in291_2 = {pp53[29],pp43[40],pp38[46],pp35[50]};
    CLA_4_c KS_291(s291, c291, in291_1, in291_2, pp51[31]);
    wire[3:0] s292, in292_1, in292_2;
    wire c292;
    assign in292_1 = {pp23[63],pp24[63],pp25[63],pp26[63]};
    assign in292_2 = {pp24[62],pp25[62],pp26[62],pp27[62]};
    CLA_4 KS_292(s292, c292, in292_1, in292_2);
    wire[2:0] s293, in293_1, in293_2;
    wire c293;
    assign in293_1 = {pp25[61],pp26[61],pp27[61]};
    assign in293_2 = {pp26[60],pp27[60],pp28[60]};
    CLA_3 KS_293(s293, c293, in293_1, in293_2);
    wire[1:0] s294, in294_1, in294_2;
    wire c294;
    assign in294_1 = {pp27[59],pp28[59]};
    assign in294_2 = {pp28[58],pp29[58]};
    CLA_2 KS_294(s294, c294, in294_1, in294_2);
    wire[0:0] s295, in295_1, in295_2;
    wire c295;
    assign in295_1 = {pp29[57]};
    assign in295_2 = {pp30[56]};
    Half_Adder KS_295(s295, c295, in295_1, in295_2);
    wire[3:0] s296, in296_1, in296_2;
    wire c296;
    assign in296_1 = {pp31[55],pp30[57],pp29[59],pp28[61]};
    assign in296_2 = {pp32[54],pp31[56],pp30[58],pp29[60]};
    CLA_4 KS_296(s296, c296, in296_1, in296_2);
    wire[0:0] s297, in297_1, in297_2;
    wire c297;
    assign in297_1 = {pp33[53]};
    assign in297_2 = {pp34[52]};
    Half_Adder KS_297(s297, c297, in297_1, in297_2);
    wire[1:0] s298, in298_1, in298_2;
    wire c298;
    assign in298_1 = {pp35[51],pp32[55]};
    assign in298_2 = {pp36[50],pp33[54]};
    CLA_2 KS_298(s298, c298, in298_1, in298_2);
    wire[0:0] s299, in299_1, in299_2;
    wire c299;
    assign in299_1 = {pp37[49]};
    assign in299_2 = {pp38[48]};
    Half_Adder KS_299(s299, c299, in299_1, in299_2);
    wire[2:0] s300, in300_1, in300_2;
    wire c300;
    assign in300_1 = {pp40[46],pp34[53],pp31[57]};
    assign in300_2 = {pp41[45],pp35[52],pp32[56]};
    CLA_3_c KS_300(s300, c300, in300_1, in300_2, pp39[47]);
    wire[0:0] s301, in301_1, in301_2;
    wire c301;
    assign in301_1 = {pp27[63]};
    assign in301_2 = {pp28[62]};
    Half_Adder KS_301(s301, c301, in301_1, in301_2);

    /*Stage 2*/
    wire[3:0] s302, in302_1, in302_2;
    wire c302;
    assign in302_1 = {pp0[23],pp0[24],pp0[25],pp0[26]};
    assign in302_2 = {pp1[22],pp1[23],pp1[24],pp1[25]};
    CLA_4 KS_302(s302, c302, in302_1, in302_2);
    wire[3:0] s303, in303_1, in303_2;
    wire c303;
    assign in303_1 = {pp2[22],pp2[23],pp2[24],pp0[27]};
    assign in303_2 = {pp3[21],pp3[22],pp3[23],pp1[26]};
    CLA_4 KS_303(s303, c303, in303_1, in303_2);
    wire[3:0] s304, in304_1, in304_2;
    wire c304;
    assign in304_1 = {pp4[21],pp4[22],pp2[25],pp0[28]};
    assign in304_2 = {pp5[20],pp5[21],pp3[24],pp1[27]};
    CLA_4 KS_304(s304, c304, in304_1, in304_2);
    wire[3:0] s305, in305_1, in305_2;
    wire c305;
    assign in305_1 = {pp6[20],pp4[23],pp2[26],pp0[29]};
    assign in305_2 = {pp7[19],pp5[22],pp3[25],pp1[28]};
    CLA_4 KS_305(s305, c305, in305_1, in305_2);
    wire[3:0] s306, in306_1, in306_2;
    wire c306;
    assign in306_1 = {pp6[21],pp4[24],pp2[27],pp0[30]};
    assign in306_2 = {pp7[20],pp5[23],pp3[26],pp1[29]};
    CLA_4 KS_306(s306, c306, in306_1, in306_2);
    wire[3:0] s307, in307_1, in307_2;
    wire c307;
    assign in307_1 = {pp9[18],pp6[22],pp4[25],pp2[28]};
    assign in307_2 = {pp10[17],pp7[21],pp5[24],pp3[27]};
    CLA_4_c KS_307(s307, c307, in307_1, in307_2, pp8[19]);
    wire[3:0] s308, in308_1, in308_2;
    wire c308;
    assign in308_1 = {pp8[20],pp6[23],pp4[26],pp0[31]};
    assign in308_2 = {pp9[19],pp7[22],pp5[25],pp1[30]};
    CLA_4 KS_308(s308, c308, in308_1, in308_2);
    wire[3:0] s309, in309_1, in309_2;
    wire c309;
    assign in309_1 = {pp11[17],pp8[21],pp6[24],pp2[29]};
    assign in309_2 = {pp12[16],pp9[20],pp7[23],pp3[28]};
    CLA_4_c KS_309(s309, c309, in309_1, in309_2, pp10[18]);
    wire[3:0] s310, in310_1, in310_2;
    wire c310;
    assign in310_1 = {pp10[19],pp8[22],pp4[27],pp0[32]};
    assign in310_2 = {pp11[18],pp9[21],pp5[26],pp1[31]};
    CLA_4 KS_310(s310, c310, in310_1, in310_2);
    wire[3:0] s311, in311_1, in311_2;
    wire c311;
    assign in311_1 = {pp13[16],pp10[20],pp6[25],pp2[30]};
    assign in311_2 = {pp14[15],pp11[19],pp7[24],pp3[29]};
    CLA_4_c KS_311(s311, c311, in311_1, in311_2, pp12[17]);
    wire[3:0] s312, in312_1, in312_2;
    wire c312;
    assign in312_1 = {pp12[18],pp8[23],pp4[28],pp0[33]};
    assign in312_2 = {pp13[17],pp9[22],pp5[27],pp1[32]};
    CLA_4 KS_312(s312, c312, in312_1, in312_2);
    wire[3:0] s313, in313_1, in313_2;
    wire c313;
    assign in313_1 = {pp15[15],pp10[21],pp6[26],pp2[31]};
    assign in313_2 = {pp16[14],pp11[20],pp7[25],pp3[30]};
    CLA_4_c KS_313(s313, c313, in313_1, in313_2, pp14[16]);
    wire[3:0] s314, in314_1, in314_2;
    wire c314;
    assign in314_1 = {pp12[19],pp8[24],pp4[29],pp0[34]};
    assign in314_2 = {pp13[18],pp9[23],pp5[28],pp1[33]};
    CLA_4 KS_314(s314, c314, in314_1, in314_2);
    wire[3:0] s315, in315_1, in315_2;
    wire c315;
    assign in315_1 = {pp14[17],pp10[22],pp6[27],pp2[32]};
    assign in315_2 = {pp15[16],pp11[21],pp7[26],pp3[31]};
    CLA_4 KS_315(s315, c315, in315_1, in315_2);
    wire[3:0] s316, in316_1, in316_2;
    wire c316;
    assign in316_1 = {pp16[15],pp12[20],pp8[25],pp4[30]};
    assign in316_2 = {pp17[14],pp13[19],pp9[24],pp5[29]};
    CLA_4 KS_316(s316, c316, in316_1, in316_2);
    wire[3:0] s317, in317_1, in317_2;
    wire c317;
    assign in317_1 = {pp19[12],pp14[18],pp10[23],pp6[28]};
    assign in317_2 = {pp20[11],pp15[17],pp11[22],pp7[27]};
    CLA_4_c KS_317(s317, c317, in317_1, in317_2, pp18[13]);
    wire[3:0] s318, in318_1, in318_2;
    wire c318;
    assign in318_1 = {pp16[16],pp12[21],pp8[26],pp0[35]};
    assign in318_2 = {pp17[15],pp13[20],pp9[25],pp1[34]};
    CLA_4 KS_318(s318, c318, in318_1, in318_2);
    wire[3:0] s319, in319_1, in319_2;
    wire c319;
    assign in319_1 = {pp18[14],pp14[19],pp10[24],pp2[33]};
    assign in319_2 = {pp19[13],pp15[18],pp11[23],pp3[32]};
    CLA_4 KS_319(s319, c319, in319_1, in319_2);
    wire[3:0] s320, in320_1, in320_2;
    wire c320;
    assign in320_1 = {pp21[11],pp16[17],pp12[22],pp4[31]};
    assign in320_2 = {pp22[10],pp17[16],pp13[21],pp5[30]};
    CLA_4_c KS_320(s320, c320, in320_1, in320_2, pp20[12]);
    wire[3:0] s321, in321_1, in321_2;
    wire c321;
    assign in321_1 = {pp18[15],pp14[20],pp6[29],pp0[36]};
    assign in321_2 = {pp19[14],pp15[19],pp7[28],pp1[35]};
    CLA_4 KS_321(s321, c321, in321_1, in321_2);
    wire[3:0] s322, in322_1, in322_2;
    wire c322;
    assign in322_1 = {pp20[13],pp16[18],pp8[27],pp2[34]};
    assign in322_2 = {pp21[12],pp17[17],pp9[26],pp3[33]};
    CLA_4 KS_322(s322, c322, in322_1, in322_2);
    wire[3:0] s323, in323_1, in323_2;
    wire c323;
    assign in323_1 = {pp23[10],pp18[16],pp10[25],pp4[32]};
    assign in323_2 = {pp24[9],pp19[15],pp11[24],pp5[31]};
    CLA_4_c KS_323(s323, c323, in323_1, in323_2, pp22[11]);
    wire[3:0] s324, in324_1, in324_2;
    wire c324;
    assign in324_1 = {pp20[14],pp12[23],pp6[30],pp0[37]};
    assign in324_2 = {pp21[13],pp13[22],pp7[29],pp1[36]};
    CLA_4 KS_324(s324, c324, in324_1, in324_2);
    wire[3:0] s325, in325_1, in325_2;
    wire c325;
    assign in325_1 = {pp22[12],pp14[21],pp8[28],pp2[35]};
    assign in325_2 = {pp23[11],pp15[20],pp9[27],pp3[34]};
    CLA_4 KS_325(s325, c325, in325_1, in325_2);
    wire[3:0] s326, in326_1, in326_2;
    wire c326;
    assign in326_1 = {pp25[9],pp16[19],pp10[26],pp4[33]};
    assign in326_2 = {pp26[8],pp17[18],pp11[25],pp5[32]};
    CLA_4_c KS_326(s326, c326, in326_1, in326_2, pp24[10]);
    wire[3:0] s327, in327_1, in327_2;
    wire c327;
    assign in327_1 = {pp18[17],pp12[24],pp6[31],pp2[36]};
    assign in327_2 = {pp19[16],pp13[23],pp7[30],pp3[35]};
    CLA_4 KS_327(s327, c327, in327_1, in327_2);
    wire[3:0] s328, in328_1, in328_2;
    wire c328;
    assign in328_1 = {pp20[15],pp14[22],pp8[29],pp4[34]};
    assign in328_2 = {pp21[14],pp15[21],pp9[28],pp5[33]};
    CLA_4 KS_328(s328, c328, in328_1, in328_2);
    wire[3:0] s329, in329_1, in329_2;
    wire c329;
    assign in329_1 = {pp22[13],pp16[20],pp10[27],pp6[32]};
    assign in329_2 = {pp23[12],pp17[19],pp11[26],pp7[31]};
    CLA_4 KS_329(s329, c329, in329_1, in329_2);
    wire[3:0] s330, in330_1, in330_2;
    wire c330;
    assign in330_1 = {pp24[11],pp18[18],pp12[25],pp8[30]};
    assign in330_2 = {pp25[10],pp19[17],pp13[24],pp9[29]};
    CLA_4 KS_330(s330, c330, in330_1, in330_2);
    wire[3:0] s331, in331_1, in331_2;
    wire c331;
    assign in331_1 = {pp26[9],pp20[16],pp14[23],pp10[28]};
    assign in331_2 = {pp27[8],pp21[15],pp15[22],pp11[27]};
    CLA_4 KS_331(s331, c331, in331_1, in331_2);
    wire[3:0] s332, in332_1, in332_2;
    wire c332;
    assign in332_1 = {pp28[7],pp22[14],pp16[21],pp12[26]};
    assign in332_2 = {pp29[6],pp23[13],pp17[20],pp13[25]};
    CLA_4 KS_332(s332, c332, in332_1, in332_2);
    wire[3:0] s333, in333_1, in333_2;
    wire c333;
    assign in333_1 = {pp31[4],pp24[12],pp18[19],pp14[24]};
    assign in333_2 = {pp32[3],pp25[11],pp19[18],pp15[23]};
    CLA_4_c KS_333(s333, c333, in333_1, in333_2, pp30[5]);
    wire[3:0] s334, in334_1, in334_2;
    wire c334;
    assign in334_1 = {pp26[10],pp20[17],pp16[22],pp4[35]};
    assign in334_2 = {pp27[9],pp21[16],pp17[21],pp5[34]};
    CLA_4 KS_334(s334, c334, in334_1, in334_2);
    wire[3:0] s335, in335_1, in335_2;
    wire c335;
    assign in335_1 = {pp28[8],pp22[15],pp18[20],pp6[33]};
    assign in335_2 = {pp29[7],pp23[14],pp19[19],pp7[32]};
    CLA_4 KS_335(s335, c335, in335_1, in335_2);
    wire[3:0] s336, in336_1, in336_2;
    wire c336;
    assign in336_1 = {pp31[5],pp24[13],pp20[18],pp8[31]};
    assign in336_2 = {pp32[4],pp25[12],pp21[17],pp9[30]};
    CLA_4_c KS_336(s336, c336, in336_1, in336_2, pp30[6]);
    wire[3:0] s337, in337_1, in337_2;
    wire c337;
    assign in337_1 = {pp26[11],pp22[16],pp10[29],pp6[34]};
    assign in337_2 = {pp27[10],pp23[15],pp11[28],pp7[33]};
    CLA_4 KS_337(s337, c337, in337_1, in337_2);
    wire[3:0] s338, in338_1, in338_2;
    wire c338;
    assign in338_1 = {pp28[9],pp24[14],pp12[27],pp8[32]};
    assign in338_2 = {pp29[8],pp25[13],pp13[26],pp9[31]};
    CLA_4 KS_338(s338, c338, in338_1, in338_2);
    wire[3:0] s339, in339_1, in339_2;
    wire c339;
    assign in339_1 = {pp30[7],pp26[12],pp14[25],pp10[30]};
    assign in339_2 = {pp31[6],pp27[11],pp15[24],pp11[29]};
    CLA_4 KS_339(s339, c339, in339_1, in339_2);
    wire[3:0] s340, in340_1, in340_2;
    wire c340;
    assign in340_1 = {pp33[4],pp28[10],pp16[23],pp12[28]};
    assign in340_2 = {pp34[3],pp29[9],pp17[22],pp13[27]};
    CLA_4_c KS_340(s340, c340, in340_1, in340_2, pp32[5]);
    wire[3:0] s341, in341_1, in341_2;
    wire c341;
    assign in341_1 = {pp30[8],pp18[21],pp14[26],pp8[33]};
    assign in341_2 = {pp31[7],pp19[20],pp15[25],pp9[32]};
    CLA_4 KS_341(s341, c341, in341_1, in341_2);
    wire[3:0] s342, in342_1, in342_2;
    wire c342;
    assign in342_1 = {pp32[6],pp20[19],pp16[24],pp10[31]};
    assign in342_2 = {pp33[5],pp21[18],pp17[23],pp11[30]};
    CLA_4 KS_342(s342, c342, in342_1, in342_2);
    wire[3:0] s343, in343_1, in343_2;
    wire c343;
    assign in343_1 = {pp35[3],pp22[17],pp18[22],pp12[29]};
    assign in343_2 = {pp36[2],pp23[16],pp19[21],pp13[28]};
    CLA_4_c KS_343(s343, c343, in343_1, in343_2, pp34[4]);
    wire[3:0] s344, in344_1, in344_2;
    wire c344;
    assign in344_1 = {pp24[15],pp20[20],pp14[27],pp11[31]};
    assign in344_2 = {pp25[14],pp21[19],pp15[26],pp12[30]};
    CLA_4 KS_344(s344, c344, in344_1, in344_2);
    wire[3:0] s345, in345_1, in345_2;
    wire c345;
    assign in345_1 = {pp26[13],pp22[18],pp16[25],pp13[29]};
    assign in345_2 = {pp27[12],pp23[17],pp17[24],pp14[28]};
    CLA_4 KS_345(s345, c345, in345_1, in345_2);
    wire[3:0] s346, in346_1, in346_2;
    wire c346;
    assign in346_1 = {pp28[11],pp24[16],pp18[23],pp15[27]};
    assign in346_2 = {pp29[10],pp25[15],pp19[22],pp16[26]};
    CLA_4 KS_346(s346, c346, in346_1, in346_2);
    wire[3:0] s347, in347_1, in347_2;
    wire c347;
    assign in347_1 = {pp30[9],pp26[14],pp20[21],pp17[25]};
    assign in347_2 = {pp31[8],pp27[13],pp21[20],pp18[24]};
    CLA_4 KS_347(s347, c347, in347_1, in347_2);
    wire[3:0] s348, in348_1, in348_2;
    wire c348;
    assign in348_1 = {pp32[7],pp28[12],pp22[19],pp19[23]};
    assign in348_2 = {pp33[6],pp29[11],pp23[18],pp20[22]};
    CLA_4 KS_348(s348, c348, in348_1, in348_2);
    wire[3:0] s349, in349_1, in349_2;
    wire c349;
    assign in349_1 = {pp34[5],pp30[10],pp24[17],pp21[21]};
    assign in349_2 = {pp35[4],pp31[9],pp25[16],pp22[20]};
    CLA_4 KS_349(s349, c349, in349_1, in349_2);
    wire[3:0] s350, in350_1, in350_2;
    wire c350;
    assign in350_1 = {pp36[3],pp32[8],pp26[15],pp23[19]};
    assign in350_2 = {pp37[2],pp33[7],pp27[14],pp24[18]};
    CLA_4 KS_350(s350, c350, in350_1, in350_2);
    wire[3:0] s351, in351_1, in351_2;
    wire c351;
    assign in351_1 = {pp38[1],pp34[6],pp28[13],pp25[17]};
    assign in351_2 = {pp39[0],pp35[5],pp29[12],pp26[16]};
    CLA_4 KS_351(s351, c351, in351_1, in351_2);
    wire[3:0] s352, in352_1, in352_2;
    wire c352;
    assign in352_1 = {s1[1],pp36[4],pp30[11],pp27[15]};
    assign in352_2 = {s2[0],pp37[3],pp31[10],pp28[14]};
    CLA_4 KS_352(s352, c352, in352_1, in352_2);
    wire[3:0] s353, in353_1, in353_2;
    wire c353;
    assign in353_1 = {c327,pp38[2],pp32[9],pp29[13]};
    assign in353_2 = {c328,pp39[1],pp33[8],pp30[12]};
    CLA_4 KS_353(s353, c353, in353_1, in353_2);
    wire[3:0] s354, in354_1, in354_2;
    wire c354;
    assign in354_1 = {c330,pp40[0],pp34[7],pp31[11]};
    assign in354_2 = {c331,s1[2],pp35[6],pp32[10]};
    CLA_4_c KS_354(s354, c354, in354_1, in354_2, c329);
    wire[3:0] s355, in355_1, in355_2;
    wire c355;
    assign in355_1 = {pp36[5],pp33[9],pp13[30],pp15[29]};
    assign in355_2 = {pp37[4],pp34[8],pp14[29],pp16[28]};
    CLA_4 KS_355(s355, c355, in355_1, in355_2);
    wire[3:0] s356, in356_1, in356_2;
    wire c356;
    assign in356_1 = {pp38[3],pp35[7],pp15[28],pp17[27]};
    assign in356_2 = {pp39[2],pp36[6],pp16[27],pp18[26]};
    CLA_4 KS_356(s356, c356, in356_1, in356_2);
    wire[3:0] s357, in357_1, in357_2;
    wire c357;
    assign in357_1 = {pp40[1],pp37[5],pp17[26],pp19[25]};
    assign in357_2 = {pp41[0],pp38[4],pp18[25],pp20[24]};
    CLA_4 KS_357(s357, c357, in357_1, in357_2);
    wire[3:0] s358, in358_1, in358_2;
    wire c358;
    assign in358_1 = {s2[2],pp39[3],pp19[24],pp21[23]};
    assign in358_2 = {s3[1],pp40[2],pp20[23],pp22[22]};
    CLA_4_c KS_358(s358, c358, in358_1, in358_2, s1[3]);
    wire[3:0] s359, in359_1, in359_2;
    wire c359;
    assign in359_1 = {pp41[1],pp21[22],pp23[21],pp17[28]};
    assign in359_2 = {pp42[0],pp22[21],pp24[20],pp18[27]};
    CLA_4 KS_359(s359, c359, in359_1, in359_2);
    wire[3:0] s360, in360_1, in360_2;
    wire c360;
    assign in360_1 = {s2[3],pp23[20],pp25[19],pp19[26]};
    assign in360_2 = {s3[2],pp24[19],pp26[18],pp20[25]};
    CLA_4_c KS_360(s360, c360, in360_1, in360_2, c1);
    wire[3:0] s361, in361_1, in361_2;
    wire c361;
    assign in361_1 = {pp25[18],pp27[17],pp21[24],pp21[25]};
    assign in361_2 = {pp26[17],pp28[16],pp22[23],pp22[24]};
    CLA_4 KS_361(s361, c361, in361_1, in361_2);
    wire[3:0] s362, in362_1, in362_2;
    wire c362;
    assign in362_1 = {pp27[16],pp29[15],pp23[22],pp23[23]};
    assign in362_2 = {pp28[15],pp30[14],pp24[21],pp24[22]};
    CLA_4 KS_362(s362, c362, in362_1, in362_2);
    wire[3:0] s363, in363_1, in363_2;
    wire c363;
    assign in363_1 = {pp29[14],pp31[13],pp25[20],pp25[21]};
    assign in363_2 = {pp30[13],pp32[12],pp26[19],pp26[20]};
    CLA_4 KS_363(s363, c363, in363_1, in363_2);
    wire[3:0] s364, in364_1, in364_2;
    wire c364;
    assign in364_1 = {pp31[12],pp33[11],pp27[18],pp27[19]};
    assign in364_2 = {pp32[11],pp34[10],pp28[17],pp28[18]};
    CLA_4 KS_364(s364, c364, in364_1, in364_2);
    wire[3:0] s365, in365_1, in365_2;
    wire c365;
    assign in365_1 = {pp33[10],pp35[9],pp29[16],pp29[17]};
    assign in365_2 = {pp34[9],pp36[8],pp30[15],pp30[16]};
    CLA_4 KS_365(s365, c365, in365_1, in365_2);
    wire[3:0] s366, in366_1, in366_2;
    wire c366;
    assign in366_1 = {pp35[8],pp37[7],pp31[14],pp31[15]};
    assign in366_2 = {pp36[7],pp38[6],pp32[13],pp32[14]};
    CLA_4 KS_366(s366, c366, in366_1, in366_2);
    wire[3:0] s367, in367_1, in367_2;
    wire c367;
    assign in367_1 = {pp37[6],pp39[5],pp33[12],pp33[13]};
    assign in367_2 = {pp38[5],pp40[4],pp34[11],pp34[12]};
    CLA_4 KS_367(s367, c367, in367_1, in367_2);
    wire[3:0] s368, in368_1, in368_2;
    wire c368;
    assign in368_1 = {pp39[4],pp41[3],pp35[10],pp35[11]};
    assign in368_2 = {pp40[3],pp42[2],pp36[9],pp36[10]};
    CLA_4 KS_368(s368, c368, in368_1, in368_2);
    wire[3:0] s369, in369_1, in369_2;
    wire c369;
    assign in369_1 = {pp41[2],pp43[1],pp37[8],pp37[9]};
    assign in369_2 = {pp42[1],pp44[0],pp38[7],pp38[8]};
    CLA_4 KS_369(s369, c369, in369_1, in369_2);
    wire[3:0] s370, in370_1, in370_2;
    wire c370;
    assign in370_1 = {pp43[0],c3,pp39[6],pp39[7]};
    assign in370_2 = {c2,s4[3],pp40[5],pp40[6]};
    CLA_4 KS_370(s370, c370, in370_1, in370_2);
    wire[0:0] s371, in371_1, in371_2;
    wire c371;
    assign in371_1 = {s3[3]};
    assign in371_2 = {s4[2]};
    Half_Adder KS_371(s371, c371, in371_1, in371_2);
    wire[3:0] s372, in372_1, in372_2;
    wire c372;
    assign in372_1 = {s5[1],s5[2],pp41[4],pp41[5]};
    assign in372_2 = {s6[1],s6[2],pp42[3],pp42[4]};
    CLA_4 KS_372(s372, c372, in372_1, in372_2);
    wire[0:0] s373, in373_1, in373_2;
    wire c373;
    assign in373_1 = {s7[0]};
    assign in373_2 = {s8[0]};
    Half_Adder KS_373(s373, c373, in373_1, in373_2);
    wire[3:0] s374, in374_1, in374_2;
    wire c374;
    assign in374_1 = {c344,s7[1],pp43[2],pp43[3]};
    assign in374_2 = {c345,s8[1],pp44[1],pp44[2]};
    CLA_4 KS_374(s374, c374, in374_1, in374_2);
    wire[0:0] s375, in375_1, in375_2;
    wire c375;
    assign in375_1 = {c346};
    assign in375_2 = {c347};
    Half_Adder KS_375(s375, c375, in375_1, in375_2);
    wire[3:0] s376, in376_1, in376_2;
    wire c376;
    assign in376_1 = {c348,s9[0],pp45[0],pp45[1]};
    assign in376_2 = {c349,s10[0],c4,pp46[0]};
    CLA_4 KS_376(s376, c376, in376_1, in376_2);
    wire[0:0] s377, in377_1, in377_2;
    wire c377;
    assign in377_1 = {c350};
    assign in377_2 = {c351};
    Half_Adder KS_377(s377, c377, in377_1, in377_2);
    wire[3:0] s378, in378_1, in378_2;
    wire c378;
    assign in378_1 = {c352,s355[3],s5[3],c5};
    assign in378_2 = {c353,s356[3],s6[3],c6};
    CLA_4 KS_378(s378, c378, in378_1, in378_2);
    wire[0:0] s379, in379_1, in379_2;
    wire c379;
    assign in379_1 = {s355[2]};
    assign in379_2 = {s356[2]};
    Full_Adder KS_379(s379, c379, in379_1, in379_2, c354);
    wire[3:0] s380, in380_1, in380_2;
    wire c380;
    assign in380_1 = {s7[2],s7[3],pp23[24],pp25[23]};
    assign in380_2 = {s8[2],s8[3],pp24[23],pp26[22]};
    CLA_4 KS_380(s380, c380, in380_1, in380_2);
    wire[3:0] s381, in381_1, in381_2;
    wire c381;
    assign in381_1 = {s10[1],s9[2],pp25[22],pp27[21]};
    assign in381_2 = {s11[0],s10[2],pp26[21],pp28[20]};
    CLA_4_c KS_381(s381, c381, in381_1, in381_2, s9[1]);
    wire[3:0] s382, in382_1, in382_2;
    wire c382;
    assign in382_1 = {s11[1],pp27[20],pp29[19],pp27[22]};
    assign in382_2 = {s12[1],pp28[19],pp30[18],pp28[21]};
    CLA_4 KS_382(s382, c382, in382_1, in382_2);
    wire[3:0] s383, in383_1, in383_2;
    wire c383;
    assign in383_1 = {pp29[18],pp31[17],pp29[20],pp33[17]};
    assign in383_2 = {pp30[17],pp32[16],pp30[19],pp34[16]};
    CLA_4 KS_383(s383, c383, in383_1, in383_2);
    wire[3:0] s384, in384_1, in384_2;
    wire c384;
    assign in384_1 = {pp31[16],pp33[15],pp31[18],pp35[15]};
    assign in384_2 = {pp32[15],pp34[14],pp32[17],pp36[14]};
    CLA_4 KS_384(s384, c384, in384_1, in384_2);
    wire[3:0] s385, in385_1, in385_2;
    wire c385;
    assign in385_1 = {pp33[14],pp35[13],pp33[16],pp37[13]};
    assign in385_2 = {pp34[13],pp36[12],pp34[15],pp38[12]};
    CLA_4 KS_385(s385, c385, in385_1, in385_2);
    wire[3:0] s386, in386_1, in386_2;
    wire c386;
    assign in386_1 = {pp35[12],pp37[11],pp35[14],pp39[11]};
    assign in386_2 = {pp36[11],pp38[10],pp36[13],pp40[10]};
    CLA_4 KS_386(s386, c386, in386_1, in386_2);
    wire[3:0] s387, in387_1, in387_2;
    wire c387;
    assign in387_1 = {pp37[10],pp39[9],pp37[12],pp41[9]};
    assign in387_2 = {pp38[9],pp40[8],pp38[11],pp42[8]};
    CLA_4 KS_387(s387, c387, in387_1, in387_2);
    wire[3:0] s388, in388_1, in388_2;
    wire c388;
    assign in388_1 = {pp39[8],pp41[7],pp39[10],pp43[7]};
    assign in388_2 = {pp40[7],pp42[6],pp40[9],pp44[6]};
    CLA_4 KS_388(s388, c388, in388_1, in388_2);
    wire[3:0] s389, in389_1, in389_2;
    wire c389;
    assign in389_1 = {pp41[6],pp43[5],pp41[8],pp45[5]};
    assign in389_2 = {pp42[5],pp44[4],pp42[7],pp46[4]};
    CLA_4 KS_389(s389, c389, in389_1, in389_2);
    wire[3:0] s390, in390_1, in390_2;
    wire c390;
    assign in390_1 = {pp43[4],pp45[3],pp43[6],pp47[3]};
    assign in390_2 = {pp44[3],pp46[2],pp44[5],pp48[2]};
    CLA_4 KS_390(s390, c390, in390_1, in390_2);
    wire[3:0] s391, in391_1, in391_2;
    wire c391;
    assign in391_1 = {pp45[2],pp47[1],pp45[4],pp49[1]};
    assign in391_2 = {pp46[1],pp48[0],pp46[3],pp50[0]};
    CLA_4 KS_391(s391, c391, in391_1, in391_2);
    wire[3:0] s392, in392_1, in392_2;
    wire c392;
    assign in392_1 = {pp47[0],c9,pp47[2],c13};
    assign in392_2 = {c7,c10,pp48[1],c14};
    CLA_4 KS_392(s392, c392, in392_1, in392_2);
    wire[3:0] s393, in393_1, in393_2;
    wire c393;
    assign in393_1 = {c8,s11[3],pp49[0],c15};
    assign in393_2 = {s9[3],s12[3],c11,c16};
    CLA_4 KS_393(s393, c393, in393_1, in393_2);
    wire[3:0] s394, in394_1, in394_2;
    wire c394;
    assign in394_1 = {s10[3],s13[2],c12,s17[3]};
    assign in394_2 = {s11[2],s14[2],s13[3],s18[3]};
    CLA_4 KS_394(s394, c394, in394_1, in394_2);
    wire[3:0] s395, in395_1, in395_2;
    wire c395;
    assign in395_1 = {s12[2],s15[2],s14[3],s19[3]};
    assign in395_2 = {s13[1],s16[2],s15[3],s20[2]};
    CLA_4 KS_395(s395, c395, in395_1, in395_2);
    wire[0:0] s396, in396_1, in396_2;
    wire c396;
    assign in396_1 = {s14[1]};
    assign in396_2 = {s15[1]};
    Half_Adder KS_396(s396, c396, in396_1, in396_2);
    wire[3:0] s397, in397_1, in397_2;
    wire c397;
    assign in397_1 = {s16[1],s17[1],s16[3],s21[2]};
    assign in397_2 = {s17[0],s18[1],s17[2],s22[2]};
    CLA_4 KS_397(s397, c397, in397_1, in397_2);
    wire[0:0] s398, in398_1, in398_2;
    wire c398;
    assign in398_1 = {s18[0]};
    assign in398_2 = {s19[0]};
    Half_Adder KS_398(s398, c398, in398_1, in398_2);
    wire[3:0] s399, in399_1, in399_2;
    wire c399;
    assign in399_1 = {c361,s19[1],s18[2],s23[1]};
    assign in399_2 = {c362,s20[0],s19[2],s24[1]};
    CLA_4 KS_399(s399, c399, in399_1, in399_2);
    wire[0:0] s400, in400_1, in400_2;
    wire c400;
    assign in400_1 = {c363};
    assign in400_2 = {c364};
    Half_Adder KS_400(s400, c400, in400_1, in400_2);
    wire[3:0] s401, in401_1, in401_2;
    wire c401;
    assign in401_1 = {c365,s21[0],s20[1],s25[1]};
    assign in401_2 = {c366,s22[0],s21[1],s26[0]};
    CLA_4 KS_401(s401, c401, in401_1, in401_2);
    wire[0:0] s402, in402_1, in402_2;
    wire c402;
    assign in402_1 = {c367};
    assign in402_2 = {c368};
    Half_Adder KS_402(s402, c402, in402_1, in402_2);
    wire[3:0] s403, in403_1, in403_2;
    wire c403;
    assign in403_1 = {c369,s380[3],s22[1],s27[0]};
    assign in403_2 = {c370,s381[3],s23[0],s28[0]};
    CLA_4 KS_403(s403, c403, in403_1, in403_2);
    wire[0:0] s404, in404_1, in404_2;
    wire c404;
    assign in404_1 = {c372};
    assign in404_2 = {c374};
    Half_Adder KS_404(s404, c404, in404_1, in404_2);
    wire[1:0] s405, in405_1, in405_2;
    wire c405;
    assign in405_1 = {c376,s382[2]};
    assign in405_2 = {c378,s383[1]};
    CLA_2 KS_405(s405, c405, in405_1, in405_2);
    wire[0:0] s406, in406_1, in406_2;
    wire c406;
    assign in406_1 = {s380[2]};
    assign in406_2 = {s381[2]};
    Half_Adder KS_406(s406, c406, in406_1, in406_2);
    wire[2:0] s407, in407_1, in407_2;
    wire c407;
    assign in407_1 = {s383[0],s384[1],s24[0]};
    assign in407_2 = {s384[0],s385[1],s25[0]};
    CLA_3_c KS_407(s407, c407, in407_1, in407_2, s382[1]);
    wire[3:0] s408, in408_1, in408_2;
    wire c408;
    assign in408_1 = {pp33[18],pp35[17],pp37[16],pp47[7]};
    assign in408_2 = {pp34[17],pp36[16],pp38[15],pp48[6]};
    CLA_4 KS_408(s408, c408, in408_1, in408_2);
    wire[3:0] s409, in409_1, in409_2;
    wire c409;
    assign in409_1 = {pp35[16],pp37[15],pp39[14],pp49[5]};
    assign in409_2 = {pp36[15],pp38[14],pp40[13],pp50[4]};
    CLA_4 KS_409(s409, c409, in409_1, in409_2);
    wire[3:0] s410, in410_1, in410_2;
    wire c410;
    assign in410_1 = {pp37[14],pp39[13],pp41[12],pp51[3]};
    assign in410_2 = {pp38[13],pp40[12],pp42[11],pp52[2]};
    CLA_4 KS_410(s410, c410, in410_1, in410_2);
    wire[3:0] s411, in411_1, in411_2;
    wire c411;
    assign in411_1 = {pp39[12],pp41[11],pp43[10],pp53[1]};
    assign in411_2 = {pp40[11],pp42[10],pp44[9],pp54[0]};
    CLA_4 KS_411(s411, c411, in411_1, in411_2);
    wire[3:0] s412, in412_1, in412_2;
    wire c412;
    assign in412_1 = {pp41[10],pp43[9],pp45[8],c26};
    assign in412_2 = {pp42[9],pp44[8],pp46[7],c27};
    CLA_4 KS_412(s412, c412, in412_1, in412_2);
    wire[3:0] s413, in413_1, in413_2;
    wire c413;
    assign in413_1 = {pp43[8],pp45[7],pp47[6],c28};
    assign in413_2 = {pp44[7],pp46[6],pp48[5],c29};
    CLA_4 KS_413(s413, c413, in413_1, in413_2);
    wire[3:0] s414, in414_1, in414_2;
    wire c414;
    assign in414_1 = {pp45[6],pp47[5],pp49[4],c30};
    assign in414_2 = {pp46[5],pp48[4],pp50[3],c31};
    CLA_4 KS_414(s414, c414, in414_1, in414_2);
    wire[3:0] s415, in415_1, in415_2;
    wire c415;
    assign in415_1 = {pp47[4],pp49[3],pp51[2],c32};
    assign in415_2 = {pp48[3],pp50[2],pp52[1],s33[3]};
    CLA_4 KS_415(s415, c415, in415_1, in415_2);
    wire[3:0] s416, in416_1, in416_2;
    wire c416;
    assign in416_1 = {pp49[2],pp51[1],pp53[0],s34[3]};
    assign in416_2 = {pp50[1],pp52[0],c23,s35[3]};
    CLA_4 KS_416(s416, c416, in416_1, in416_2);
    wire[3:0] s417, in417_1, in417_2;
    wire c417;
    assign in417_1 = {pp51[0],c20,c24,s36[2]};
    assign in417_2 = {c17,c21,c25,s37[2]};
    CLA_4 KS_417(s417, c417, in417_1, in417_2);
    wire[3:0] s418, in418_1, in418_2;
    wire c418;
    assign in418_1 = {c18,c22,s26[3],s38[2]};
    assign in418_2 = {c19,s23[3],s27[3],s39[2]};
    CLA_4 KS_418(s418, c418, in418_1, in418_2);
    wire[3:0] s419, in419_1, in419_2;
    wire c419;
    assign in419_1 = {s20[3],s24[3],s28[3],s40[1]};
    assign in419_2 = {s21[3],s25[3],s29[3],s41[1]};
    CLA_4 KS_419(s419, c419, in419_1, in419_2);
    wire[3:0] s420, in420_1, in420_2;
    wire c420;
    assign in420_1 = {s22[3],s26[2],s30[3],s42[1]};
    assign in420_2 = {s23[2],s27[2],s31[3],s43[1]};
    CLA_4 KS_420(s420, c420, in420_1, in420_2);
    wire[3:0] s421, in421_1, in421_2;
    wire c421;
    assign in421_1 = {s24[2],s28[2],s32[3],s44[0]};
    assign in421_2 = {s25[2],s29[2],s33[2],s45[0]};
    CLA_4 KS_421(s421, c421, in421_1, in421_2);
    wire[3:0] s422, in422_1, in422_2;
    wire c422;
    assign in422_1 = {s26[1],s30[2],s34[2],s46[0]};
    assign in422_2 = {s27[1],s31[2],s35[2],s47[0]};
    CLA_4 KS_422(s422, c422, in422_1, in422_2);
    wire[3:0] s423, in423_1, in423_2;
    wire c423;
    assign in423_1 = {s28[1],s32[2],s36[1],s48[0]};
    assign in423_2 = {s29[1],s33[1],s37[1],s49[0]};
    CLA_4 KS_423(s423, c423, in423_1, in423_2);
    wire[0:0] s424, in424_1, in424_2;
    wire c424;
    assign in424_1 = {s30[1]};
    assign in424_2 = {s31[1]};
    Half_Adder KS_424(s424, c424, in424_1, in424_2);
    wire[1:0] s425, in425_1, in425_2;
    wire c425;
    assign in425_1 = {s32[1],s34[1]};
    assign in425_2 = {s33[0],s35[1]};
    CLA_2 KS_425(s425, c425, in425_1, in425_2);
    wire[0:0] s426, in426_1, in426_2;
    wire c426;
    assign in426_1 = {s34[0]};
    assign in426_2 = {s35[0]};
    Half_Adder KS_426(s426, c426, in426_1, in426_2);
    wire[2:0] s427, in427_1, in427_2;
    wire c427;
    assign in427_1 = {c383,s36[0],s38[1]};
    assign in427_2 = {c384,s37[0],s39[1]};
    CLA_3 KS_427(s427, c427, in427_1, in427_2);
    wire[0:0] s428, in428_1, in428_2;
    wire c428;
    assign in428_1 = {c385};
    assign in428_2 = {c386};
    Half_Adder KS_428(s428, c428, in428_1, in428_2);
    wire[1:0] s429, in429_1, in429_2;
    wire c429;
    assign in429_1 = {c387,s38[0]};
    assign in429_2 = {c388,s39[0]};
    CLA_2 KS_429(s429, c429, in429_1, in429_2);
    wire[0:0] s430, in430_1, in430_2;
    wire c430;
    assign in430_1 = {c389};
    assign in430_2 = {c390};
    Half_Adder KS_430(s430, c430, in430_1, in430_2);
    wire[3:0] s431, in431_1, in431_2;
    wire c431;
    assign in431_1 = {c391,s408[1],s40[0],s50[0]};
    assign in431_2 = {c392,s409[1],s41[0],s51[0]};
    CLA_4 KS_431(s431, c431, in431_1, in431_2);
    wire[0:0] s432, in432_1, in432_2;
    wire c432;
    assign in432_1 = {c393};
    assign in432_2 = {c394};
    Half_Adder KS_432(s432, c432, in432_1, in432_2);
    wire[1:0] s433, in433_1, in433_2;
    wire c433;
    assign in433_1 = {c395,s410[1]};
    assign in433_2 = {c397,s411[1]};
    CLA_2 KS_433(s433, c433, in433_1, in433_2);
    wire[0:0] s434, in434_1, in434_2;
    wire c434;
    assign in434_1 = {c399};
    assign in434_2 = {c401};
    Half_Adder KS_434(s434, c434, in434_1, in434_2);
    wire[2:0] s435, in435_1, in435_2;
    wire c435;
    assign in435_1 = {c403,s412[1],s42[0]};
    assign in435_2 = {s408[0],s413[1],s43[0]};
    CLA_3 KS_435(s435, c435, in435_1, in435_2);
    wire[0:0] s436, in436_1, in436_2;
    wire c436;
    assign in436_1 = {s409[0]};
    assign in436_2 = {s410[0]};
    Half_Adder KS_436(s436, c436, in436_1, in436_2);
    wire[1:0] s437, in437_1, in437_2;
    wire c437;
    assign in437_1 = {s411[0],s414[1]};
    assign in437_2 = {s412[0],s415[1]};
    CLA_2 KS_437(s437, c437, in437_1, in437_2);
    wire[0:0] s438, in438_1, in438_2;
    wire c438;
    assign in438_1 = {s414[0]};
    assign in438_2 = {s415[0]};
    Full_Adder KS_438(s438, c438, in438_1, in438_2, s413[0]);
    wire[3:0] s439, in439_1, in439_2;
    wire c439;
    assign in439_1 = {pp42[13],pp45[11],pp47[10],c50};
    assign in439_2 = {pp43[12],pp46[10],pp48[9],c51};
    CLA_4 KS_439(s439, c439, in439_1, in439_2);
    wire[3:0] s440, in440_1, in440_2;
    wire c440;
    assign in440_1 = {pp44[11],pp47[9],pp49[8],c52};
    assign in440_2 = {pp45[10],pp48[8],pp50[7],c53};
    CLA_4 KS_440(s440, c440, in440_1, in440_2);
    wire[3:0] s441, in441_1, in441_2;
    wire c441;
    assign in441_1 = {pp46[9],pp49[7],pp51[6],c54};
    assign in441_2 = {pp47[8],pp50[6],pp52[5],c55};
    CLA_4 KS_441(s441, c441, in441_1, in441_2);
    wire[3:0] s442, in442_1, in442_2;
    wire c442;
    assign in442_1 = {pp48[7],pp51[5],pp53[4],s56[3]};
    assign in442_2 = {pp49[6],pp52[4],pp54[3],s57[2]};
    CLA_4 KS_442(s442, c442, in442_1, in442_2);
    wire[3:0] s443, in443_1, in443_2;
    wire c443;
    assign in443_1 = {pp50[5],pp53[3],pp55[2],s58[2]};
    assign in443_2 = {pp51[4],pp54[2],pp56[1],s59[2]};
    CLA_4 KS_443(s443, c443, in443_1, in443_2);
    wire[3:0] s444, in444_1, in444_2;
    wire c444;
    assign in444_1 = {pp52[3],pp55[1],pp57[0],s60[2]};
    assign in444_2 = {pp53[2],pp56[0],c40,s61[2]};
    CLA_4 KS_444(s444, c444, in444_1, in444_2);
    wire[3:0] s445, in445_1, in445_2;
    wire c445;
    assign in445_1 = {pp54[1],c36,c41,s62[1]};
    assign in445_2 = {pp55[0],c37,c42,s63[1]};
    CLA_4 KS_445(s445, c445, in445_1, in445_2);
    wire[3:0] s446, in446_1, in446_2;
    wire c446;
    assign in446_1 = {c33,c38,c43,s64[1]};
    assign in446_2 = {c34,c39,s44[3],s65[1]};
    CLA_4 KS_446(s446, c446, in446_1, in446_2);
    wire[3:0] s447, in447_1, in447_2;
    wire c447;
    assign in447_1 = {c35,s40[3],s45[3],s66[1]};
    assign in447_2 = {s36[3],s41[3],s46[3],s67[0]};
    CLA_4 KS_447(s447, c447, in447_1, in447_2);
    wire[3:0] s448, in448_1, in448_2;
    wire c448;
    assign in448_1 = {s37[3],s42[3],s47[3],s68[0]};
    assign in448_2 = {s38[3],s43[3],s48[3],s69[0]};
    CLA_4 KS_448(s448, c448, in448_1, in448_2);
    wire[3:0] s449, in449_1, in449_2;
    wire c449;
    assign in449_1 = {s39[3],s44[2],s49[3],s70[0]};
    assign in449_2 = {s40[2],s45[2],s50[3],s71[0]};
    CLA_4 KS_449(s449, c449, in449_1, in449_2);
    wire[3:0] s450, in450_1, in450_2;
    wire c450;
    assign in450_1 = {s41[2],s46[2],s51[3],s72[0]};
    assign in450_2 = {s42[2],s47[2],s52[3],s73[0]};
    CLA_4 KS_450(s450, c450, in450_1, in450_2);
    wire[3:0] s451, in451_1, in451_2;
    wire c451;
    assign in451_1 = {s43[2],s48[2],s53[3],s74[0]};
    assign in451_2 = {s44[1],s49[2],s54[3],s75[0]};
    CLA_4 KS_451(s451, c451, in451_1, in451_2);
    wire[3:0] s452, in452_1, in452_2;
    wire c452;
    assign in452_1 = {s45[1],s50[2],s55[3],s76[0]};
    assign in452_2 = {s46[1],s51[2],s56[2],s77[0]};
    CLA_4 KS_452(s452, c452, in452_1, in452_2);
    wire[3:0] s453, in453_1, in453_2;
    wire c453;
    assign in453_1 = {s47[1],s52[2],s57[1],s78[0]};
    assign in453_2 = {s48[1],s53[2],s58[1],s79[0]};
    CLA_4 KS_453(s453, c453, in453_1, in453_2);
    wire[3:0] s454, in454_1, in454_2;
    wire c454;
    assign in454_1 = {s49[1],s54[2],s59[1],s80[0]};
    assign in454_2 = {s50[1],s55[2],s60[1],s81[0]};
    CLA_4 KS_454(s454, c454, in454_1, in454_2);
    wire[0:0] s455, in455_1, in455_2;
    wire c455;
    assign in455_1 = {s51[1]};
    assign in455_2 = {s52[1]};
    Half_Adder KS_455(s455, c455, in455_1, in455_2);
    wire[1:0] s456, in456_1, in456_2;
    wire c456;
    assign in456_1 = {s53[1],s56[1]};
    assign in456_2 = {s54[1],s57[0]};
    CLA_2 KS_456(s456, c456, in456_1, in456_2);
    wire[0:0] s457, in457_1, in457_2;
    wire c457;
    assign in457_1 = {s55[1]};
    assign in457_2 = {s56[0]};
    Half_Adder KS_457(s457, c457, in457_1, in457_2);
    wire[2:0] s458, in458_1, in458_2;
    wire c458;
    assign in458_1 = {c408,s58[0],s61[1]};
    assign in458_2 = {c409,s59[0],s62[0]};
    CLA_3 KS_458(s458, c458, in458_1, in458_2);
    wire[0:0] s459, in459_1, in459_2;
    wire c459;
    assign in459_1 = {c410};
    assign in459_2 = {c411};
    Half_Adder KS_459(s459, c459, in459_1, in459_2);
    wire[1:0] s460, in460_1, in460_2;
    wire c460;
    assign in460_1 = {c412,s60[0]};
    assign in460_2 = {c413,s61[0]};
    CLA_2 KS_460(s460, c460, in460_1, in460_2);
    wire[0:0] s461, in461_1, in461_2;
    wire c461;
    assign in461_1 = {c414};
    assign in461_2 = {c415};
    Half_Adder KS_461(s461, c461, in461_1, in461_2);
    wire[3:0] s462, in462_1, in462_2;
    wire c462;
    assign in462_1 = {c416,s439[1],s63[0],s82[0]};
    assign in462_2 = {c417,s440[1],s64[0],s83[0]};
    CLA_4 KS_462(s462, c462, in462_1, in462_2);
    wire[0:0] s463, in463_1, in463_2;
    wire c463;
    assign in463_1 = {c418};
    assign in463_2 = {c419};
    Half_Adder KS_463(s463, c463, in463_1, in463_2);
    wire[1:0] s464, in464_1, in464_2;
    wire c464;
    assign in464_1 = {c420,s441[1]};
    assign in464_2 = {c421,s442[1]};
    CLA_2 KS_464(s464, c464, in464_1, in464_2);
    wire[0:0] s465, in465_1, in465_2;
    wire c465;
    assign in465_1 = {c422};
    assign in465_2 = {c423};
    Half_Adder KS_465(s465, c465, in465_1, in465_2);
    wire[2:0] s466, in466_1, in466_2;
    wire c466;
    assign in466_1 = {c431,s443[1],s65[0]};
    assign in466_2 = {s439[0],s444[1],s66[0]};
    CLA_3 KS_466(s466, c466, in466_1, in466_2);
    wire[0:0] s467, in467_1, in467_2;
    wire c467;
    assign in467_1 = {s440[0]};
    assign in467_2 = {s441[0]};
    Half_Adder KS_467(s467, c467, in467_1, in467_2);
    wire[1:0] s468, in468_1, in468_2;
    wire c468;
    assign in468_1 = {s442[0],s445[1]};
    assign in468_2 = {s443[0],s446[1]};
    CLA_2 KS_468(s468, c468, in468_1, in468_2);
    wire[0:0] s469, in469_1, in469_2;
    wire c469;
    assign in469_1 = {s445[0]};
    assign in469_2 = {s446[0]};
    Full_Adder KS_469(s469, c469, in469_1, in469_2, s444[0]);
    wire[3:0] s470, in470_1, in470_2;
    wire c470;
    assign in470_1 = {pp54[5],pp55[5],pp57[4],s91[2]};
    assign in470_2 = {pp55[4],pp56[4],pp58[3],s92[2]};
    CLA_4 KS_470(s470, c470, in470_1, in470_2);
    wire[3:0] s471, in471_1, in471_2;
    wire c471;
    assign in471_1 = {pp56[3],pp57[3],pp59[2],s93[1]};
    assign in471_2 = {pp57[2],pp58[2],pp60[1],s94[1]};
    CLA_4 KS_471(s471, c471, in471_1, in471_2);
    wire[3:0] s472, in472_1, in472_2;
    wire c472;
    assign in472_1 = {pp58[1],pp59[1],pp61[0],s95[1]};
    assign in472_2 = {pp59[0],pp60[0],c62,s96[1]};
    CLA_4 KS_472(s472, c472, in472_1, in472_2);
    wire[3:0] s473, in473_1, in473_2;
    wire c473;
    assign in473_1 = {c56,c57,c63,s97[1]};
    assign in473_2 = {s57[3],c58,c64,s98[1]};
    CLA_4 KS_473(s473, c473, in473_1, in473_2);
    wire[3:0] s474, in474_1, in474_2;
    wire c474;
    assign in474_1 = {s58[3],c59,c65,s99[0]};
    assign in474_2 = {s59[3],c60,c66,s100[0]};
    CLA_4 KS_474(s474, c474, in474_1, in474_2);
    wire[3:0] s475, in475_1, in475_2;
    wire c475;
    assign in475_1 = {s60[3],c61,s67[3],s101[0]};
    assign in475_2 = {s61[3],s62[3],s68[3],s102[0]};
    CLA_4 KS_475(s475, c475, in475_1, in475_2);
    wire[3:0] s476, in476_1, in476_2;
    wire c476;
    assign in476_1 = {s62[2],s63[3],s69[3],s103[0]};
    assign in476_2 = {s63[2],s64[3],s70[3],s104[0]};
    CLA_4 KS_476(s476, c476, in476_1, in476_2);
    wire[3:0] s477, in477_1, in477_2;
    wire c477;
    assign in477_1 = {s64[2],s65[3],s71[3],s105[0]};
    assign in477_2 = {s65[2],s66[3],s72[3],s106[0]};
    CLA_4 KS_477(s477, c477, in477_1, in477_2);
    wire[3:0] s478, in478_1, in478_2;
    wire c478;
    assign in478_1 = {s66[2],s67[2],s73[3],s107[0]};
    assign in478_2 = {s67[1],s68[2],s74[3],s108[0]};
    CLA_4 KS_478(s478, c478, in478_1, in478_2);
    wire[3:0] s479, in479_1, in479_2;
    wire c479;
    assign in479_1 = {s68[1],s69[2],s75[3],s109[0]};
    assign in479_2 = {s69[1],s70[2],s76[3],s110[0]};
    CLA_4 KS_479(s479, c479, in479_1, in479_2);
    wire[3:0] s480, in480_1, in480_2;
    wire c480;
    assign in480_1 = {s70[1],s71[2],s77[3],s111[0]};
    assign in480_2 = {s71[1],s72[2],s78[3],s112[0]};
    CLA_4 KS_480(s480, c480, in480_1, in480_2);
    wire[3:0] s481, in481_1, in481_2;
    wire c481;
    assign in481_1 = {s72[1],s73[2],s79[3],s113[0]};
    assign in481_2 = {s73[1],s74[2],s80[3],s114[0]};
    CLA_4 KS_481(s481, c481, in481_1, in481_2);
    wire[3:0] s482, in482_1, in482_2;
    wire c482;
    assign in482_1 = {s74[1],s75[2],s82[3],s115[0]};
    assign in482_2 = {s75[1],s76[2],s84[3],s116[0]};
    CLA_4 KS_482(s482, c482, in482_1, in482_2);
    wire[3:0] s483, in483_1, in483_2;
    wire c483;
    assign in483_1 = {s76[1],s77[2],s86[3],s117[0]};
    assign in483_2 = {s77[1],s78[2],s88[1],s118[0]};
    CLA_4 KS_483(s483, c483, in483_1, in483_2);
    wire[3:0] s484, in484_1, in484_2;
    wire c484;
    assign in484_1 = {s78[1],s79[2],s89[1],s119[0]};
    assign in484_2 = {s79[1],s80[2],s90[1],s120[0]};
    CLA_4 KS_484(s484, c484, in484_1, in484_2);
    wire[3:0] s485, in485_1, in485_2;
    wire c485;
    assign in485_1 = {s80[1],s82[2],s91[1],s121[0]};
    assign in485_2 = {c81,s84[2],s92[1],s122[0]};
    CLA_4 KS_485(s485, c485, in485_1, in485_2);
    wire[0:0] s486, in486_1, in486_2;
    wire c486;
    assign in486_1 = {s82[1]};
    assign in486_2 = {c83};
    Half_Adder KS_486(s486, c486, in486_1, in486_2);
    wire[1:0] s487, in487_1, in487_2;
    wire c487;
    assign in487_1 = {s84[1],s86[2]};
    assign in487_2 = {c85,s88[0]};
    CLA_2 KS_487(s487, c487, in487_1, in487_2);
    wire[0:0] s488, in488_1, in488_2;
    wire c488;
    assign in488_1 = {s86[1]};
    assign in488_2 = {c87};
    Half_Adder KS_488(s488, c488, in488_1, in488_2);
    wire[2:0] s489, in489_1, in489_2;
    wire c489;
    assign in489_1 = {c439,s89[0],s93[0]};
    assign in489_2 = {c440,s90[0],s94[0]};
    CLA_3 KS_489(s489, c489, in489_1, in489_2);
    wire[0:0] s490, in490_1, in490_2;
    wire c490;
    assign in490_1 = {c441};
    assign in490_2 = {c442};
    Half_Adder KS_490(s490, c490, in490_1, in490_2);
    wire[1:0] s491, in491_1, in491_2;
    wire c491;
    assign in491_1 = {c443,s91[0]};
    assign in491_2 = {c444,s92[0]};
    CLA_2 KS_491(s491, c491, in491_1, in491_2);
    wire[0:0] s492, in492_1, in492_2;
    wire c492;
    assign in492_1 = {c445};
    assign in492_2 = {c446};
    Half_Adder KS_492(s492, c492, in492_1, in492_2);
    wire[3:0] s493, in493_1, in493_2;
    wire c493;
    assign in493_1 = {c447,s470[1],s95[0],s123[0]};
    assign in493_2 = {c448,s471[1],s96[0],s124[0]};
    CLA_4 KS_493(s493, c493, in493_1, in493_2);
    wire[0:0] s494, in494_1, in494_2;
    wire c494;
    assign in494_1 = {c449};
    assign in494_2 = {c450};
    Half_Adder KS_494(s494, c494, in494_1, in494_2);
    wire[1:0] s495, in495_1, in495_2;
    wire c495;
    assign in495_1 = {c451,s472[1]};
    assign in495_2 = {c452,s473[1]};
    CLA_2 KS_495(s495, c495, in495_1, in495_2);
    wire[0:0] s496, in496_1, in496_2;
    wire c496;
    assign in496_1 = {c453};
    assign in496_2 = {c454};
    Half_Adder KS_496(s496, c496, in496_1, in496_2);
    wire[2:0] s497, in497_1, in497_2;
    wire c497;
    assign in497_1 = {c462,s474[1],s97[0]};
    assign in497_2 = {s470[0],s475[1],s98[0]};
    CLA_3 KS_497(s497, c497, in497_1, in497_2);
    wire[0:0] s498, in498_1, in498_2;
    wire c498;
    assign in498_1 = {s471[0]};
    assign in498_2 = {s472[0]};
    Half_Adder KS_498(s498, c498, in498_1, in498_2);
    wire[1:0] s499, in499_1, in499_2;
    wire c499;
    assign in499_1 = {s473[0],s476[1]};
    assign in499_2 = {s474[0],s477[1]};
    CLA_2 KS_499(s499, c499, in499_1, in499_2);
    wire[0:0] s500, in500_1, in500_2;
    wire c500;
    assign in500_1 = {s476[0]};
    assign in500_2 = {s477[0]};
    Full_Adder KS_500(s500, c500, in500_1, in500_2, s475[0]);
    wire[3:0] s501, in501_1, in501_2;
    wire c501;
    assign in501_1 = {s92[3],pp62[2],pp61[4],s136[0]};
    assign in501_2 = {s93[2],pp63[1],pp62[3],s137[0]};
    CLA_4 KS_501(s501, c501, in501_1, in501_2);
    wire[3:0] s502, in502_1, in502_2;
    wire c502;
    assign in502_1 = {s94[2],1'b0,pp63[2],s138[0]};
    assign in502_2 = {s95[2],c88,c93,s139[0]};
    CLA_4 KS_502(s502, c502, in502_1, in502_2);
    wire[3:0] s503, in503_1, in503_2;
    wire c503;
    assign in503_1 = {s96[2],c89,c94,s140[0]};
    assign in503_2 = {s97[2],c90,c95,s141[0]};
    CLA_4 KS_503(s503, c503, in503_1, in503_2);
    wire[3:0] s504, in504_1, in504_2;
    wire c504;
    assign in504_1 = {s98[2],c91,c96,s142[0]};
    assign in504_2 = {s99[1],c92,c97,s143[0]};
    CLA_4 KS_504(s504, c504, in504_1, in504_2);
    wire[3:0] s505, in505_1, in505_2;
    wire c505;
    assign in505_1 = {s100[1],s93[3],c98,s144[0]};
    assign in505_2 = {s101[1],s94[3],s99[3],s145[0]};
    CLA_4 KS_505(s505, c505, in505_1, in505_2);
    wire[3:0] s506, in506_1, in506_2;
    wire c506;
    assign in506_1 = {s102[1],s95[3],s100[3],s146[0]};
    assign in506_2 = {s103[1],s96[3],s101[3],s147[0]};
    CLA_4 KS_506(s506, c506, in506_1, in506_2);
    wire[3:0] s507, in507_1, in507_2;
    wire c507;
    assign in507_1 = {s104[1],s97[3],s102[3],s148[0]};
    assign in507_2 = {s105[1],s98[3],s103[3],s149[0]};
    CLA_4 KS_507(s507, c507, in507_1, in507_2);
    wire[3:0] s508, in508_1, in508_2;
    wire c508;
    assign in508_1 = {s106[1],s99[2],s104[3],s150[0]};
    assign in508_2 = {s107[1],s100[2],s105[3],s151[0]};
    CLA_4 KS_508(s508, c508, in508_1, in508_2);
    wire[3:0] s509, in509_1, in509_2;
    wire c509;
    assign in509_1 = {s108[1],s101[2],s106[3],s152[0]};
    assign in509_2 = {s109[1],s102[2],s107[3],s153[0]};
    CLA_4 KS_509(s509, c509, in509_1, in509_2);
    wire[3:0] s510, in510_1, in510_2;
    wire c510;
    assign in510_1 = {s110[1],s103[2],s108[3],s154[0]};
    assign in510_2 = {s111[1],s104[2],s109[3],s155[0]};
    CLA_4 KS_510(s510, c510, in510_1, in510_2);
    wire[3:0] s511, in511_1, in511_2;
    wire c511;
    assign in511_1 = {s112[1],s105[2],s110[3],s156[0]};
    assign in511_2 = {s113[1],s106[2],s111[3],s157[0]};
    CLA_4 KS_511(s511, c511, in511_1, in511_2);
    wire[3:0] s512, in512_1, in512_2;
    wire c512;
    assign in512_1 = {s114[1],s107[2],s112[3],s158[0]};
    assign in512_2 = {c115,s108[2],s113[3],s159[0]};
    CLA_4 KS_512(s512, c512, in512_1, in512_2);
    wire[3:0] s513, in513_1, in513_2;
    wire c513;
    assign in513_1 = {s116[1],s109[2],s114[3],s160[0]};
    assign in513_2 = {c117,s110[2],s116[3],s161[0]};
    CLA_4 KS_513(s513, c513, in513_1, in513_2);
    wire[3:0] s514, in514_1, in514_2;
    wire c514;
    assign in514_1 = {s118[1],s111[2],s118[3],s162[0]};
    assign in514_2 = {c119,s112[2],s120[3],s163[0]};
    CLA_4 KS_514(s514, c514, in514_1, in514_2);
    wire[3:0] s515, in515_1, in515_2;
    wire c515;
    assign in515_1 = {s120[1],s113[2],s122[3],s164[0]};
    assign in515_2 = {c121,s114[2],s124[3],s165[0]};
    CLA_4 KS_515(s515, c515, in515_1, in515_2);
    wire[3:0] s516, in516_1, in516_2;
    wire c516;
    assign in516_1 = {s122[1],s116[2],s126[3],s166[0]};
    assign in516_2 = {c123,s118[2],s128[3],s167[0]};
    CLA_4 KS_516(s516, c516, in516_1, in516_2);
    wire[0:0] s517, in517_1, in517_2;
    wire c517;
    assign in517_1 = {s124[1]};
    assign in517_2 = {c125};
    Half_Adder KS_517(s517, c517, in517_1, in517_2);
    wire[1:0] s518, in518_1, in518_2;
    wire c518;
    assign in518_1 = {s126[1],s120[2]};
    assign in518_2 = {c127,s122[2]};
    CLA_2 KS_518(s518, c518, in518_1, in518_2);
    wire[0:0] s519, in519_1, in519_2;
    wire c519;
    assign in519_1 = {s128[1]};
    assign in519_2 = {c470};
    Half_Adder KS_519(s519, c519, in519_1, in519_2);
    wire[2:0] s520, in520_1, in520_2;
    wire c520;
    assign in520_1 = {c471,s124[2],s129[1]};
    assign in520_2 = {c472,s126[2],s130[0]};
    CLA_3 KS_520(s520, c520, in520_1, in520_2);
    wire[0:0] s521, in521_1, in521_2;
    wire c521;
    assign in521_1 = {c473};
    assign in521_2 = {c474};
    Half_Adder KS_521(s521, c521, in521_1, in521_2);
    wire[1:0] s522, in522_1, in522_2;
    wire c522;
    assign in522_1 = {c475,s128[2]};
    assign in522_2 = {c476,s129[0]};
    CLA_2 KS_522(s522, c522, in522_1, in522_2);
    wire[0:0] s523, in523_1, in523_2;
    wire c523;
    assign in523_1 = {c477};
    assign in523_2 = {c478};
    Half_Adder KS_523(s523, c523, in523_1, in523_2);
    wire[3:0] s524, in524_1, in524_2;
    wire c524;
    assign in524_1 = {c479,s501[1],s131[0],s168[0]};
    assign in524_2 = {c480,s502[1],s132[0],s169[0]};
    CLA_4 KS_524(s524, c524, in524_1, in524_2);
    wire[0:0] s525, in525_1, in525_2;
    wire c525;
    assign in525_1 = {c481};
    assign in525_2 = {c482};
    Half_Adder KS_525(s525, c525, in525_1, in525_2);
    wire[1:0] s526, in526_1, in526_2;
    wire c526;
    assign in526_1 = {c483,s503[1]};
    assign in526_2 = {c484,s504[1]};
    CLA_2 KS_526(s526, c526, in526_1, in526_2);
    wire[0:0] s527, in527_1, in527_2;
    wire c527;
    assign in527_1 = {c485};
    assign in527_2 = {c493};
    Half_Adder KS_527(s527, c527, in527_1, in527_2);
    wire[2:0] s528, in528_1, in528_2;
    wire c528;
    assign in528_1 = {s501[0],s505[1],s133[0]};
    assign in528_2 = {s502[0],s506[1],s134[0]};
    CLA_3 KS_528(s528, c528, in528_1, in528_2);
    wire[0:0] s529, in529_1, in529_2;
    wire c529;
    assign in529_1 = {s503[0]};
    assign in529_2 = {s504[0]};
    Half_Adder KS_529(s529, c529, in529_1, in529_2);
    wire[1:0] s530, in530_1, in530_2;
    wire c530;
    assign in530_1 = {s506[0],s507[1]};
    assign in530_2 = {s507[0],s508[1]};
    CLA_2_c KS_530(s530, c530, in530_1, in530_2, s505[0]);
    wire[3:0] s531, in531_1, in531_2;
    wire c531;
    assign in531_1 = {s137[1],pp61[7],pp55[14],s177[0]};
    assign in531_2 = {s138[1],pp62[6],pp56[13],s178[0]};
    CLA_4 KS_531(s531, c531, in531_1, in531_2);
    wire[3:0] s532, in532_1, in532_2;
    wire c532;
    assign in532_1 = {s139[1],pp63[5],pp57[12],s179[0]};
    assign in532_2 = {s140[1],c129,pp58[11],s180[0]};
    CLA_4 KS_532(s532, c532, in532_1, in532_2);
    wire[3:0] s533, in533_1, in533_2;
    wire c533;
    assign in533_1 = {s141[1],s130[3],pp59[10],s181[0]};
    assign in533_2 = {s142[1],s131[3],pp60[9],s182[0]};
    CLA_4 KS_533(s533, c533, in533_1, in533_2);
    wire[3:0] s534, in534_1, in534_2;
    wire c534;
    assign in534_1 = {s143[1],s132[3],pp61[8],s183[0]};
    assign in534_2 = {s144[1],s133[3],pp62[7],s184[0]};
    CLA_4 KS_534(s534, c534, in534_1, in534_2);
    wire[3:0] s535, in535_1, in535_2;
    wire c535;
    assign in535_1 = {s145[1],s134[3],pp63[6],s185[0]};
    assign in535_2 = {s146[1],s135[2],c130,s186[0]};
    CLA_4 KS_535(s535, c535, in535_1, in535_2);
    wire[3:0] s536, in536_1, in536_2;
    wire c536;
    assign in536_1 = {s147[1],s136[2],c131,s187[0]};
    assign in536_2 = {s148[1],s137[2],c132,s188[0]};
    CLA_4 KS_536(s536, c536, in536_1, in536_2);
    wire[3:0] s537, in537_1, in537_2;
    wire c537;
    assign in537_1 = {s149[1],s138[2],c133,s189[0]};
    assign in537_2 = {s150[1],s139[2],c134,s190[0]};
    CLA_4 KS_537(s537, c537, in537_1, in537_2);
    wire[3:0] s538, in538_1, in538_2;
    wire c538;
    assign in538_1 = {s151[1],s140[2],s135[3],s191[0]};
    assign in538_2 = {c152,s141[2],s136[3],s192[0]};
    CLA_4 KS_538(s538, c538, in538_1, in538_2);
    wire[3:0] s539, in539_1, in539_2;
    wire c539;
    assign in539_1 = {s153[1],s142[2],s137[3],s193[0]};
    assign in539_2 = {c154,s143[2],s138[3],s194[0]};
    CLA_4 KS_539(s539, c539, in539_1, in539_2);
    wire[3:0] s540, in540_1, in540_2;
    wire c540;
    assign in540_1 = {s155[1],s144[2],s139[3],s195[0]};
    assign in540_2 = {c156,s145[2],s140[3],s196[0]};
    CLA_4 KS_540(s540, c540, in540_1, in540_2);
    wire[3:0] s541, in541_1, in541_2;
    wire c541;
    assign in541_1 = {s157[1],s146[2],s141[3],s197[0]};
    assign in541_2 = {c158,s147[2],s142[3],s198[0]};
    CLA_4 KS_541(s541, c541, in541_1, in541_2);
    wire[3:0] s542, in542_1, in542_2;
    wire c542;
    assign in542_1 = {s159[1],s148[2],s143[3],s199[0]};
    assign in542_2 = {c160,s149[2],s144[3],s200[0]};
    CLA_4 KS_542(s542, c542, in542_1, in542_2);
    wire[3:0] s543, in543_1, in543_2;
    wire c543;
    assign in543_1 = {s161[1],s150[2],s145[3],s201[0]};
    assign in543_2 = {c162,s151[2],s146[3],s202[0]};
    CLA_4 KS_543(s543, c543, in543_1, in543_2);
    wire[3:0] s544, in544_1, in544_2;
    wire c544;
    assign in544_1 = {s163[1],s153[2],s147[3],s203[0]};
    assign in544_2 = {c164,c155,s148[3],s204[0]};
    CLA_4 KS_544(s544, c544, in544_1, in544_2);
    wire[3:0] s545, in545_1, in545_2;
    wire c545;
    assign in545_1 = {s165[1],s157[2],s149[3],s205[0]};
    assign in545_2 = {c166,c159,s150[3],s206[0]};
    CLA_4 KS_545(s545, c545, in545_1, in545_2);
    wire[0:0] s546, in546_1, in546_2;
    wire c546;
    assign in546_1 = {s167[1]};
    assign in546_2 = {c168};
    Half_Adder KS_546(s546, c546, in546_1, in546_2);
    wire[3:0] s547, in547_1, in547_2;
    wire c547;
    assign in547_1 = {s169[1],s161[2],s151[3],s207[0]};
    assign in547_2 = {c170,c163,s153[3],s208[0]};
    CLA_4 KS_547(s547, c547, in547_1, in547_2);
    wire[0:0] s548, in548_1, in548_2;
    wire c548;
    assign in548_1 = {s171[1]};
    assign in548_2 = {c172};
    Half_Adder KS_548(s548, c548, in548_1, in548_2);
    wire[1:0] s549, in549_1, in549_2;
    wire c549;
    assign in549_1 = {s173[1],s165[2]};
    assign in549_2 = {c501,c167};
    CLA_2 KS_549(s549, c549, in549_1, in549_2);
    wire[0:0] s550, in550_1, in550_2;
    wire c550;
    assign in550_1 = {c502};
    assign in550_2 = {c503};
    Half_Adder KS_550(s550, c550, in550_1, in550_2);
    wire[2:0] s551, in551_1, in551_2;
    wire c551;
    assign in551_1 = {c504,s169[2],s157[3]};
    assign in551_2 = {c505,c171,s161[3]};
    CLA_3 KS_551(s551, c551, in551_1, in551_2);
    wire[0:0] s552, in552_1, in552_2;
    wire c552;
    assign in552_1 = {c506};
    assign in552_2 = {c507};
    Half_Adder KS_552(s552, c552, in552_1, in552_2);
    wire[1:0] s553, in553_1, in553_2;
    wire c553;
    assign in553_1 = {c508,s173[2]};
    assign in553_2 = {c509,s531[1]};
    CLA_2 KS_553(s553, c553, in553_1, in553_2);
    wire[0:0] s554, in554_1, in554_2;
    wire c554;
    assign in554_1 = {c510};
    assign in554_2 = {c511};
    Half_Adder KS_554(s554, c554, in554_1, in554_2);
    wire[3:0] s555, in555_1, in555_2;
    wire c555;
    assign in555_1 = {c512,s532[1],s165[3],s209[0]};
    assign in555_2 = {c513,s533[1],s169[3],s210[0]};
    CLA_4 KS_555(s555, c555, in555_1, in555_2);
    wire[0:0] s556, in556_1, in556_2;
    wire c556;
    assign in556_1 = {c514};
    assign in556_2 = {c515};
    Half_Adder KS_556(s556, c556, in556_1, in556_2);
    wire[1:0] s557, in557_1, in557_2;
    wire c557;
    assign in557_1 = {c516,s534[1]};
    assign in557_2 = {c524,s535[1]};
    CLA_2 KS_557(s557, c557, in557_1, in557_2);
    wire[0:0] s558, in558_1, in558_2;
    wire c558;
    assign in558_1 = {s531[0]};
    assign in558_2 = {s532[0]};
    Half_Adder KS_558(s558, c558, in558_1, in558_2);
    wire[2:0] s559, in559_1, in559_2;
    wire c559;
    assign in559_1 = {s533[0],s536[1],s173[3]};
    assign in559_2 = {s534[0],s537[1],s174[0]};
    CLA_3 KS_559(s559, c559, in559_1, in559_2);
    wire[0:0] s560, in560_1, in560_2;
    wire c560;
    assign in560_1 = {s536[0]};
    assign in560_2 = {s537[0]};
    Full_Adder KS_560(s560, c560, in560_1, in560_2, s535[0]);
    wire[3:0] s561, in561_1, in561_2;
    wire c561;
    assign in561_1 = {s178[1],pp57[15],pp50[23],c191};
    assign in561_2 = {s179[1],pp58[14],pp51[22],c194};
    CLA_4 KS_561(s561, c561, in561_1, in561_2);
    wire[3:0] s562, in562_1, in562_2;
    wire c562;
    assign in562_1 = {s180[1],pp59[13],pp52[21],c202};
    assign in562_2 = {s181[1],pp60[12],pp53[20],c210};
    CLA_4 KS_562(s562, c562, in562_1, in562_2);
    wire[3:0] s563, in563_1, in563_2;
    wire c563;
    assign in563_1 = {s182[1],pp61[11],pp54[19],s215[0]};
    assign in563_2 = {s183[1],pp62[10],pp55[18],s216[0]};
    CLA_4 KS_563(s563, c563, in563_1, in563_2);
    wire[3:0] s564, in564_1, in564_2;
    wire c564;
    assign in564_1 = {s184[1],pp63[9],pp56[17],s217[0]};
    assign in564_2 = {s185[1],s174[3],pp57[16],s218[0]};
    CLA_4 KS_564(s564, c564, in564_1, in564_2);
    wire[3:0] s565, in565_1, in565_2;
    wire c565;
    assign in565_1 = {s186[1],s175[2],pp58[15],s219[0]};
    assign in565_2 = {s187[1],s176[2],pp59[14],s220[0]};
    CLA_4 KS_565(s565, c565, in565_1, in565_2);
    wire[3:0] s566, in566_1, in566_2;
    wire c566;
    assign in566_1 = {s188[1],s177[2],pp60[13],s221[0]};
    assign in566_2 = {s189[1],s178[2],pp61[12],s222[0]};
    CLA_4 KS_566(s566, c566, in566_1, in566_2);
    wire[3:0] s567, in567_1, in567_2;
    wire c567;
    assign in567_1 = {s190[1],s179[2],pp62[11],s223[0]};
    assign in567_2 = {s191[1],s180[2],pp63[10],s224[0]};
    CLA_4 KS_567(s567, c567, in567_1, in567_2);
    wire[3:0] s568, in568_1, in568_2;
    wire c568;
    assign in568_1 = {s192[1],s181[2],c174,s225[0]};
    assign in568_2 = {c193,s182[2],s175[3],s226[0]};
    CLA_4 KS_568(s568, c568, in568_1, in568_2);
    wire[3:0] s569, in569_1, in569_2;
    wire c569;
    assign in569_1 = {s194[1],s183[2],s176[3],s227[0]};
    assign in569_2 = {c195,s184[2],s177[3],s228[0]};
    CLA_4 KS_569(s569, c569, in569_1, in569_2);
    wire[3:0] s570, in570_1, in570_2;
    wire c570;
    assign in570_1 = {s196[1],s185[2],s178[3],s229[0]};
    assign in570_2 = {c197,s186[2],s179[3],s230[0]};
    CLA_4 KS_570(s570, c570, in570_1, in570_2);
    wire[3:0] s571, in571_1, in571_2;
    wire c571;
    assign in571_1 = {s198[1],s187[2],s180[3],s231[0]};
    assign in571_2 = {c199,s188[2],s181[3],s232[0]};
    CLA_4 KS_571(s571, c571, in571_1, in571_2);
    wire[3:0] s572, in572_1, in572_2;
    wire c572;
    assign in572_1 = {s200[1],s189[2],s182[3],s233[0]};
    assign in572_2 = {c201,s190[2],s183[3],s234[0]};
    CLA_4 KS_572(s572, c572, in572_1, in572_2);
    wire[3:0] s573, in573_1, in573_2;
    wire c573;
    assign in573_1 = {s202[1],s191[2],s184[3],s235[0]};
    assign in573_2 = {c203,c192,s185[3],s236[0]};
    CLA_4 KS_573(s573, c573, in573_1, in573_2);
    wire[3:0] s574, in574_1, in574_2;
    wire c574;
    assign in574_1 = {s204[1],s194[2],s186[3],s237[0]};
    assign in574_2 = {c205,c196,s187[3],s238[0]};
    CLA_4 KS_574(s574, c574, in574_1, in574_2);
    wire[3:0] s575, in575_1, in575_2;
    wire c575;
    assign in575_1 = {s206[1],s198[2],s188[3],s239[0]};
    assign in575_2 = {c207,c200,s189[3],s240[0]};
    CLA_4 KS_575(s575, c575, in575_1, in575_2);
    wire[0:0] s576, in576_1, in576_2;
    wire c576;
    assign in576_1 = {s208[1]};
    assign in576_2 = {c209};
    Half_Adder KS_576(s576, c576, in576_1, in576_2);
    wire[3:0] s577, in577_1, in577_2;
    wire c577;
    assign in577_1 = {s210[1],s202[2],s190[3],s241[0]};
    assign in577_2 = {c211,c204,s191[3],s242[0]};
    CLA_4 KS_577(s577, c577, in577_1, in577_2);
    wire[0:0] s578, in578_1, in578_2;
    wire c578;
    assign in578_1 = {s212[1]};
    assign in578_2 = {c213};
    Half_Adder KS_578(s578, c578, in578_1, in578_2);
    wire[1:0] s579, in579_1, in579_2;
    wire c579;
    assign in579_1 = {s214[1],s206[2]};
    assign in579_2 = {c531,c208};
    CLA_2 KS_579(s579, c579, in579_1, in579_2);
    wire[0:0] s580, in580_1, in580_2;
    wire c580;
    assign in580_1 = {c532};
    assign in580_2 = {c533};
    Half_Adder KS_580(s580, c580, in580_1, in580_2);
    wire[2:0] s581, in581_1, in581_2;
    wire c581;
    assign in581_1 = {c534,s210[2],s194[3]};
    assign in581_2 = {c535,c212,c198};
    CLA_3 KS_581(s581, c581, in581_1, in581_2);
    wire[0:0] s582, in582_1, in582_2;
    wire c582;
    assign in582_1 = {c536};
    assign in582_2 = {c537};
    Half_Adder KS_582(s582, c582, in582_1, in582_2);
    wire[1:0] s583, in583_1, in583_2;
    wire c583;
    assign in583_1 = {c538,s214[2]};
    assign in583_2 = {c539,s561[1]};
    CLA_2 KS_583(s583, c583, in583_1, in583_2);
    wire[0:0] s584, in584_1, in584_2;
    wire c584;
    assign in584_1 = {c540};
    assign in584_2 = {c541};
    Half_Adder KS_584(s584, c584, in584_1, in584_2);
    wire[3:0] s585, in585_1, in585_2;
    wire c585;
    assign in585_1 = {c542,s562[1],s202[3],s243[0]};
    assign in585_2 = {c543,s563[1],c206,s244[0]};
    CLA_4 KS_585(s585, c585, in585_1, in585_2);
    wire[0:0] s586, in586_1, in586_2;
    wire c586;
    assign in586_1 = {c544};
    assign in586_2 = {c545};
    Half_Adder KS_586(s586, c586, in586_1, in586_2);
    wire[1:0] s587, in587_1, in587_2;
    wire c587;
    assign in587_1 = {c547,s564[1]};
    assign in587_2 = {c555,s565[1]};
    CLA_2 KS_587(s587, c587, in587_1, in587_2);
    wire[0:0] s588, in588_1, in588_2;
    wire c588;
    assign in588_1 = {s561[0]};
    assign in588_2 = {s562[0]};
    Half_Adder KS_588(s588, c588, in588_1, in588_2);
    wire[2:0] s589, in589_1, in589_2;
    wire c589;
    assign in589_1 = {s563[0],s566[1],s210[3]};
    assign in589_2 = {s564[0],s567[1],c214};
    CLA_3 KS_589(s589, c589, in589_1, in589_2);
    wire[0:0] s590, in590_1, in590_2;
    wire c590;
    assign in590_1 = {s566[0]};
    assign in590_2 = {s567[0]};
    Full_Adder KS_590(s590, c590, in590_1, in590_2, s565[0]);
    wire[3:0] s591, in591_1, in591_2;
    wire c591;
    assign in591_1 = {pp60[15],pp51[25],pp46[31],c219};
    assign in591_2 = {pp61[14],pp52[24],pp47[30],c220};
    CLA_4 KS_591(s591, c591, in591_1, in591_2);
    wire[3:0] s592, in592_1, in592_2;
    wire c592;
    assign in592_1 = {pp62[13],pp53[23],pp48[29],c221};
    assign in592_2 = {pp63[12],pp54[22],pp49[28],c222};
    CLA_4 KS_592(s592, c592, in592_1, in592_2);
    wire[3:0] s593, in593_1, in593_2;
    wire c593;
    assign in593_1 = {s215[1],pp55[21],pp50[27],c223};
    assign in593_2 = {s216[1],pp56[20],pp51[26],c224};
    CLA_4 KS_593(s593, c593, in593_1, in593_2);
    wire[3:0] s594, in594_1, in594_2;
    wire c594;
    assign in594_1 = {s217[1],pp57[19],pp52[25],c225};
    assign in594_2 = {s218[1],pp58[18],pp53[24],c226};
    CLA_4 KS_594(s594, c594, in594_1, in594_2);
    wire[3:0] s595, in595_1, in595_2;
    wire c595;
    assign in595_1 = {s219[1],pp59[17],pp54[23],c227};
    assign in595_2 = {s220[1],pp60[16],pp55[22],c231};
    CLA_4 KS_595(s595, c595, in595_1, in595_2);
    wire[3:0] s596, in596_1, in596_2;
    wire c596;
    assign in596_1 = {s221[1],pp61[15],pp56[21],c239};
    assign in596_2 = {s222[1],pp62[14],pp57[20],c247};
    CLA_4 KS_596(s596, c596, in596_1, in596_2);
    wire[3:0] s597, in597_1, in597_2;
    wire c597;
    assign in597_1 = {s223[1],pp63[13],pp58[19],s249[0]};
    assign in597_2 = {s224[1],s215[2],pp59[18],s250[0]};
    CLA_4 KS_597(s597, c597, in597_1, in597_2);
    wire[3:0] s598, in598_1, in598_2;
    wire c598;
    assign in598_1 = {s225[1],s216[2],pp60[17],s251[0]};
    assign in598_2 = {s226[1],s217[2],pp61[16],s252[0]};
    CLA_4 KS_598(s598, c598, in598_1, in598_2);
    wire[3:0] s599, in599_1, in599_2;
    wire c599;
    assign in599_1 = {s227[1],s218[2],pp62[15],s253[0]};
    assign in599_2 = {s228[1],s219[2],pp63[14],s254[0]};
    CLA_4 KS_599(s599, c599, in599_1, in599_2);
    wire[3:0] s600, in600_1, in600_2;
    wire c600;
    assign in600_1 = {s229[1],s220[2],s215[3],s255[0]};
    assign in600_2 = {c230,s221[2],s216[3],s256[0]};
    CLA_4 KS_600(s600, c600, in600_1, in600_2);
    wire[3:0] s601, in601_1, in601_2;
    wire c601;
    assign in601_1 = {s231[1],s222[2],s217[3],s257[0]};
    assign in601_2 = {c232,s223[2],s218[3],s258[0]};
    CLA_4 KS_601(s601, c601, in601_1, in601_2);
    wire[3:0] s602, in602_1, in602_2;
    wire c602;
    assign in602_1 = {s233[1],s224[2],s219[3],s259[0]};
    assign in602_2 = {c234,s225[2],s220[3],s260[0]};
    CLA_4 KS_602(s602, c602, in602_1, in602_2);
    wire[3:0] s603, in603_1, in603_2;
    wire c603;
    assign in603_1 = {s235[1],s226[2],s221[3],s261[0]};
    assign in603_2 = {c236,s227[2],s222[3],s262[0]};
    CLA_4 KS_603(s603, c603, in603_1, in603_2);
    wire[3:0] s604, in604_1, in604_2;
    wire c604;
    assign in604_1 = {s237[1],s228[2],s223[3],s263[0]};
    assign in604_2 = {c238,c229,s224[3],s264[0]};
    CLA_4 KS_604(s604, c604, in604_1, in604_2);
    wire[3:0] s605, in605_1, in605_2;
    wire c605;
    assign in605_1 = {s239[1],s231[2],s225[3],s265[0]};
    assign in605_2 = {c240,c233,s226[3],s266[0]};
    CLA_4 KS_605(s605, c605, in605_1, in605_2);
    wire[0:0] s606, in606_1, in606_2;
    wire c606;
    assign in606_1 = {s241[1]};
    assign in606_2 = {c242};
    Half_Adder KS_606(s606, c606, in606_1, in606_2);
    wire[1:0] s607, in607_1, in607_2;
    wire c607;
    assign in607_1 = {s243[1],s235[2]};
    assign in607_2 = {c244,c237};
    CLA_2 KS_607(s607, c607, in607_1, in607_2);
    wire[0:0] s608, in608_1, in608_2;
    wire c608;
    assign in608_1 = {s245[1]};
    assign in608_2 = {c246};
    Half_Adder KS_608(s608, c608, in608_1, in608_2);
    wire[3:0] s609, in609_1, in609_2;
    wire c609;
    assign in609_1 = {s247[1],s239[2],s227[3],s267[0]};
    assign in609_2 = {c248,c241,c228,s268[0]};
    CLA_4 KS_609(s609, c609, in609_1, in609_2);
    wire[0:0] s610, in610_1, in610_2;
    wire c610;
    assign in610_1 = {c561};
    assign in610_2 = {c562};
    Half_Adder KS_610(s610, c610, in610_1, in610_2);
    wire[1:0] s611, in611_1, in611_2;
    wire c611;
    assign in611_1 = {c563,s243[2]};
    assign in611_2 = {c564,c245};
    CLA_2 KS_611(s611, c611, in611_1, in611_2);
    wire[0:0] s612, in612_1, in612_2;
    wire c612;
    assign in612_1 = {c565};
    assign in612_2 = {c566};
    Half_Adder KS_612(s612, c612, in612_1, in612_2);
    wire[2:0] s613, in613_1, in613_2;
    wire c613;
    assign in613_1 = {c567,s247[2],s231[3]};
    assign in613_2 = {c568,s591[1],c235};
    CLA_3 KS_613(s613, c613, in613_1, in613_2);
    wire[0:0] s614, in614_1, in614_2;
    wire c614;
    assign in614_1 = {c569};
    assign in614_2 = {c570};
    Half_Adder KS_614(s614, c614, in614_1, in614_2);
    wire[1:0] s615, in615_1, in615_2;
    wire c615;
    assign in615_1 = {c571,s592[1]};
    assign in615_2 = {c572,s593[1]};
    CLA_2 KS_615(s615, c615, in615_1, in615_2);
    wire[0:0] s616, in616_1, in616_2;
    wire c616;
    assign in616_1 = {c573};
    assign in616_2 = {c574};
    Half_Adder KS_616(s616, c616, in616_1, in616_2);
    wire[3:0] s617, in617_1, in617_2;
    wire c617;
    assign in617_1 = {c575,s594[1],s239[3],s269[0]};
    assign in617_2 = {c577,s595[1],c243,s270[0]};
    CLA_4 KS_617(s617, c617, in617_1, in617_2);
    wire[0:0] s618, in618_1, in618_2;
    wire c618;
    assign in618_1 = {c585};
    assign in618_2 = {s591[0]};
    Half_Adder KS_618(s618, c618, in618_1, in618_2);
    wire[1:0] s619, in619_1, in619_2;
    wire c619;
    assign in619_1 = {s592[0],s596[1]};
    assign in619_2 = {s593[0],s597[1]};
    CLA_2 KS_619(s619, c619, in619_1, in619_2);
    wire[0:0] s620, in620_1, in620_2;
    wire c620;
    assign in620_1 = {s594[0]};
    assign in620_2 = {s595[0]};
    Half_Adder KS_620(s620, c620, in620_1, in620_2);
    wire[2:0] s621, in621_1, in621_2;
    wire c621;
    assign in621_1 = {s597[0],s598[1],s247[3]};
    assign in621_2 = {s598[0],s599[1],s591[2]};
    CLA_3_c KS_621(s621, c621, in621_1, in621_2, s596[0]);
    wire[3:0] s622, in622_1, in622_2;
    wire c622;
    assign in622_1 = {pp52[27],pp45[35],pp40[41],pp54[28]};
    assign in622_2 = {pp53[26],pp46[34],pp41[40],pp55[27]};
    CLA_4 KS_622(s622, c622, in622_1, in622_2);
    wire[3:0] s623, in623_1, in623_2;
    wire c623;
    assign in623_1 = {pp54[25],pp47[33],pp42[39],pp56[26]};
    assign in623_2 = {pp55[24],pp48[32],pp43[38],pp57[25]};
    CLA_4 KS_623(s623, c623, in623_1, in623_2);
    wire[3:0] s624, in624_1, in624_2;
    wire c624;
    assign in624_1 = {pp56[23],pp49[31],pp44[37],pp58[24]};
    assign in624_2 = {pp57[22],pp50[30],pp45[36],pp59[23]};
    CLA_4 KS_624(s624, c624, in624_1, in624_2);
    wire[3:0] s625, in625_1, in625_2;
    wire c625;
    assign in625_1 = {pp58[21],pp51[29],pp46[35],pp60[22]};
    assign in625_2 = {pp59[20],pp52[28],pp47[34],pp61[21]};
    CLA_4 KS_625(s625, c625, in625_1, in625_2);
    wire[3:0] s626, in626_1, in626_2;
    wire c626;
    assign in626_1 = {pp60[19],pp53[27],pp48[33],pp62[20]};
    assign in626_2 = {pp61[18],pp54[26],pp49[32],pp63[19]};
    CLA_4 KS_626(s626, c626, in626_1, in626_2);
    wire[3:0] s627, in627_1, in627_2;
    wire c627;
    assign in627_1 = {pp62[17],pp55[25],pp50[31],c249};
    assign in627_2 = {pp63[16],pp56[24],pp51[30],c250};
    CLA_4 KS_627(s627, c627, in627_1, in627_2);
    wire[3:0] s628, in628_1, in628_2;
    wire c628;
    assign in628_1 = {s249[1],pp57[23],pp52[29],c251};
    assign in628_2 = {s250[1],pp58[22],pp53[28],c252};
    CLA_4 KS_628(s628, c628, in628_1, in628_2);
    wire[3:0] s629, in629_1, in629_2;
    wire c629;
    assign in629_1 = {s251[1],pp59[21],pp54[27],c253};
    assign in629_2 = {s252[1],pp60[20],pp55[26],c254};
    CLA_4 KS_629(s629, c629, in629_1, in629_2);
    wire[3:0] s630, in630_1, in630_2;
    wire c630;
    assign in630_1 = {s253[1],pp61[19],pp56[25],c255};
    assign in630_2 = {s254[1],pp62[18],pp57[24],c256};
    CLA_4 KS_630(s630, c630, in630_1, in630_2);
    wire[3:0] s631, in631_1, in631_2;
    wire c631;
    assign in631_1 = {s255[1],pp63[17],pp58[23],c257};
    assign in631_2 = {s256[1],s249[2],pp59[22],c261};
    CLA_4 KS_631(s631, c631, in631_1, in631_2);
    wire[3:0] s632, in632_1, in632_2;
    wire c632;
    assign in632_1 = {s257[1],s250[2],pp60[21],c269};
    assign in632_2 = {s258[1],s251[2],pp61[20],s275[0]};
    CLA_4 KS_632(s632, c632, in632_1, in632_2);
    wire[3:0] s633, in633_1, in633_2;
    wire c633;
    assign in633_1 = {s259[1],s252[2],pp62[19],s276[0]};
    assign in633_2 = {c260,s253[2],pp63[18],s277[0]};
    CLA_4 KS_633(s633, c633, in633_1, in633_2);
    wire[3:0] s634, in634_1, in634_2;
    wire c634;
    assign in634_1 = {s261[1],s254[2],s249[3],s278[0]};
    assign in634_2 = {c262,s255[2],s250[3],s279[0]};
    CLA_4 KS_634(s634, c634, in634_1, in634_2);
    wire[3:0] s635, in635_1, in635_2;
    wire c635;
    assign in635_1 = {s263[1],s256[2],s251[3],s280[0]};
    assign in635_2 = {c264,s257[2],s252[3],s281[0]};
    CLA_4 KS_635(s635, c635, in635_1, in635_2);
    wire[3:0] s636, in636_1, in636_2;
    wire c636;
    assign in636_1 = {s265[1],s258[2],s253[3],s282[0]};
    assign in636_2 = {c266,c259,s254[3],s283[0]};
    CLA_4 KS_636(s636, c636, in636_1, in636_2);
    wire[0:0] s637, in637_1, in637_2;
    wire c637;
    assign in637_1 = {s267[1]};
    assign in637_2 = {c268};
    Half_Adder KS_637(s637, c637, in637_1, in637_2);
    wire[3:0] s638, in638_1, in638_2;
    wire c638;
    assign in638_1 = {s269[1],s261[2],s255[3],s284[0]};
    assign in638_2 = {c270,c263,s256[3],s285[0]};
    CLA_4 KS_638(s638, c638, in638_1, in638_2);
    wire[0:0] s639, in639_1, in639_2;
    wire c639;
    assign in639_1 = {s271[1]};
    assign in639_2 = {c272};
    Half_Adder KS_639(s639, c639, in639_1, in639_2);
    wire[1:0] s640, in640_1, in640_2;
    wire c640;
    assign in640_1 = {s273[1],s265[2]};
    assign in640_2 = {c274,c267};
    CLA_2 KS_640(s640, c640, in640_1, in640_2);
    wire[0:0] s641, in641_1, in641_2;
    wire c641;
    assign in641_1 = {c591};
    assign in641_2 = {c592};
    Half_Adder KS_641(s641, c641, in641_1, in641_2);
    wire[2:0] s642, in642_1, in642_2;
    wire c642;
    assign in642_1 = {c593,s269[2],s257[3]};
    assign in642_2 = {c594,c271,c258};
    CLA_3 KS_642(s642, c642, in642_1, in642_2);
    wire[0:0] s643, in643_1, in643_2;
    wire c643;
    assign in643_1 = {c595};
    assign in643_2 = {c596};
    Half_Adder KS_643(s643, c643, in643_1, in643_2);
    wire[1:0] s644, in644_1, in644_2;
    wire c644;
    assign in644_1 = {c597,s273[2]};
    assign in644_2 = {c598,s622[1]};
    CLA_2 KS_644(s644, c644, in644_1, in644_2);
    wire[0:0] s645, in645_1, in645_2;
    wire c645;
    assign in645_1 = {c599};
    assign in645_2 = {c600};
    Half_Adder KS_645(s645, c645, in645_1, in645_2);
    wire[3:0] s646, in646_1, in646_2;
    wire c646;
    assign in646_1 = {c601,s623[1],s261[3],s286[0]};
    assign in646_2 = {c602,s624[1],c265,s287[0]};
    CLA_4 KS_646(s646, c646, in646_1, in646_2);
    wire[0:0] s647, in647_1, in647_2;
    wire c647;
    assign in647_1 = {c603};
    assign in647_2 = {c604};
    Half_Adder KS_647(s647, c647, in647_1, in647_2);
    wire[1:0] s648, in648_1, in648_2;
    wire c648;
    assign in648_1 = {c605,s625[1]};
    assign in648_2 = {c609,s626[1]};
    CLA_2 KS_648(s648, c648, in648_1, in648_2);
    wire[0:0] s649, in649_1, in649_2;
    wire c649;
    assign in649_1 = {c617};
    assign in649_2 = {s622[0]};
    Half_Adder KS_649(s649, c649, in649_1, in649_2);
    wire[2:0] s650, in650_1, in650_2;
    wire c650;
    assign in650_1 = {s623[0],s627[1],s269[3]};
    assign in650_2 = {s624[0],s628[1],c273};
    CLA_3 KS_650(s650, c650, in650_1, in650_2);
    wire[0:0] s651, in651_1, in651_2;
    wire c651;
    assign in651_1 = {s625[0]};
    assign in651_2 = {s626[0]};
    Half_Adder KS_651(s651, c651, in651_1, in651_2);
    wire[1:0] s652, in652_1, in652_2;
    wire c652;
    assign in652_1 = {s628[0],s629[1]};
    assign in652_2 = {s629[0],s630[1]};
    CLA_2_c KS_652(s652, c652, in652_1, in652_2, s627[0]);
    wire[3:0] s653, in653_1, in653_2;
    wire c653;
    assign in653_1 = {pp44[39],pp39[45],pp36[49],pp42[44]};
    assign in653_2 = {pp45[38],pp40[44],pp37[48],pp43[43]};
    CLA_4 KS_653(s653, c653, in653_1, in653_2);
    wire[3:0] s654, in654_1, in654_2;
    wire c654;
    assign in654_1 = {pp46[37],pp41[43],pp38[47],pp44[42]};
    assign in654_2 = {pp47[36],pp42[42],pp39[46],pp45[41]};
    CLA_4 KS_654(s654, c654, in654_1, in654_2);
    wire[3:0] s655, in655_1, in655_2;
    wire c655;
    assign in655_1 = {pp48[35],pp43[41],pp40[45],pp46[40]};
    assign in655_2 = {pp49[34],pp44[40],pp41[44],pp47[39]};
    CLA_4 KS_655(s655, c655, in655_1, in655_2);
    wire[3:0] s656, in656_1, in656_2;
    wire c656;
    assign in656_1 = {pp50[33],pp45[39],pp42[43],pp48[38]};
    assign in656_2 = {pp51[32],pp46[38],pp43[42],pp49[37]};
    CLA_4 KS_656(s656, c656, in656_1, in656_2);
    wire[3:0] s657, in657_1, in657_2;
    wire c657;
    assign in657_1 = {pp52[31],pp47[37],pp44[41],pp50[36]};
    assign in657_2 = {pp53[30],pp48[36],pp45[40],pp51[35]};
    CLA_4 KS_657(s657, c657, in657_1, in657_2);
    wire[3:0] s658, in658_1, in658_2;
    wire c658;
    assign in658_1 = {pp54[29],pp49[35],pp46[39],pp52[34]};
    assign in658_2 = {pp55[28],pp50[34],pp47[38],pp53[33]};
    CLA_4 KS_658(s658, c658, in658_1, in658_2);
    wire[3:0] s659, in659_1, in659_2;
    wire c659;
    assign in659_1 = {pp56[27],pp51[33],pp48[37],pp54[32]};
    assign in659_2 = {pp57[26],pp52[32],pp49[36],pp55[31]};
    CLA_4 KS_659(s659, c659, in659_1, in659_2);
    wire[3:0] s660, in660_1, in660_2;
    wire c660;
    assign in660_1 = {pp58[25],pp53[31],pp50[35],pp56[30]};
    assign in660_2 = {pp59[24],pp54[30],pp51[34],pp57[29]};
    CLA_4 KS_660(s660, c660, in660_1, in660_2);
    wire[3:0] s661, in661_1, in661_2;
    wire c661;
    assign in661_1 = {pp60[23],pp55[29],pp52[33],pp58[28]};
    assign in661_2 = {pp61[22],pp56[28],pp53[32],pp59[27]};
    CLA_4 KS_661(s661, c661, in661_1, in661_2);
    wire[3:0] s662, in662_1, in662_2;
    wire c662;
    assign in662_1 = {pp62[21],pp57[27],pp54[31],pp60[26]};
    assign in662_2 = {pp63[20],pp58[26],pp55[30],pp61[25]};
    CLA_4 KS_662(s662, c662, in662_1, in662_2);
    wire[3:0] s663, in663_1, in663_2;
    wire c663;
    assign in663_1 = {s275[1],pp59[25],pp56[29],pp62[24]};
    assign in663_2 = {s276[1],pp60[24],pp57[28],pp63[23]};
    CLA_4 KS_663(s663, c663, in663_1, in663_2);
    wire[3:0] s664, in664_1, in664_2;
    wire c664;
    assign in664_1 = {s277[1],pp61[23],pp58[27],c275};
    assign in664_2 = {s278[1],pp62[22],pp59[26],c276};
    CLA_4 KS_664(s664, c664, in664_1, in664_2);
    wire[3:0] s665, in665_1, in665_2;
    wire c665;
    assign in665_1 = {s279[1],pp63[21],pp60[25],c277};
    assign in665_2 = {s280[1],s275[2],pp61[24],c278};
    CLA_4 KS_665(s665, c665, in665_1, in665_2);
    wire[3:0] s666, in666_1, in666_2;
    wire c666;
    assign in666_1 = {s281[1],s276[2],pp62[23],c279};
    assign in666_2 = {c282,s277[2],pp63[22],c283};
    CLA_4 KS_666(s666, c666, in666_1, in666_2);
    wire[3:0] s667, in667_1, in667_2;
    wire c667;
    assign in667_1 = {s283[1],s278[2],s275[3],c291};
    assign in667_2 = {c284,s279[2],s276[3],s292[0]};
    CLA_4 KS_667(s667, c667, in667_1, in667_2);
    wire[0:0] s668, in668_1, in668_2;
    wire c668;
    assign in668_1 = {s285[1]};
    assign in668_2 = {c286};
    Half_Adder KS_668(s668, c668, in668_1, in668_2);
    wire[1:0] s669, in669_1, in669_2;
    wire c669;
    assign in669_1 = {s287[1],s280[2]};
    assign in669_2 = {c288,c281};
    CLA_2 KS_669(s669, c669, in669_1, in669_2);
    wire[0:0] s670, in670_1, in670_2;
    wire c670;
    assign in670_1 = {s289[1]};
    assign in670_2 = {c290};
    Half_Adder KS_670(s670, c670, in670_1, in670_2);
    wire[3:0] s671, in671_1, in671_2;
    wire c671;
    assign in671_1 = {s291[1],s283[2],s277[3],s293[0]};
    assign in671_2 = {c622,c285,s278[3],s294[0]};
    CLA_4 KS_671(s671, c671, in671_1, in671_2);
    wire[0:0] s672, in672_1, in672_2;
    wire c672;
    assign in672_1 = {c623};
    assign in672_2 = {c624};
    Half_Adder KS_672(s672, c672, in672_1, in672_2);
    wire[1:0] s673, in673_1, in673_2;
    wire c673;
    assign in673_1 = {c625,s287[2]};
    assign in673_2 = {c626,c289};
    CLA_2 KS_673(s673, c673, in673_1, in673_2);
    wire[0:0] s674, in674_1, in674_2;
    wire c674;
    assign in674_1 = {c627};
    assign in674_2 = {c628};
    Half_Adder KS_674(s674, c674, in674_1, in674_2);
    wire[2:0] s675, in675_1, in675_2;
    wire c675;
    assign in675_1 = {c629,s291[2],s279[3]};
    assign in675_2 = {c630,s653[1],c280};
    CLA_3 KS_675(s675, c675, in675_1, in675_2);
    wire[0:0] s676, in676_1, in676_2;
    wire c676;
    assign in676_1 = {c631};
    assign in676_2 = {c632};
    Half_Adder KS_676(s676, c676, in676_1, in676_2);
    wire[1:0] s677, in677_1, in677_2;
    wire c677;
    assign in677_1 = {c633,s654[1]};
    assign in677_2 = {c634,s655[1]};
    CLA_2 KS_677(s677, c677, in677_1, in677_2);
    wire[0:0] s678, in678_1, in678_2;
    wire c678;
    assign in678_1 = {c635};
    assign in678_2 = {c636};
    Half_Adder KS_678(s678, c678, in678_1, in678_2);
    wire[3:0] s679, in679_1, in679_2;
    wire c679;
    assign in679_1 = {c638,s656[1],s283[3],s295[0]};
    assign in679_2 = {c646,s657[1],c287,s296[0]};
    CLA_4 KS_679(s679, c679, in679_1, in679_2);
    wire[0:0] s680, in680_1, in680_2;
    wire c680;
    assign in680_1 = {s653[0]};
    assign in680_2 = {s654[0]};
    Half_Adder KS_680(s680, c680, in680_1, in680_2);
    wire[1:0] s681, in681_1, in681_2;
    wire c681;
    assign in681_1 = {s655[0],s658[1]};
    assign in681_2 = {s656[0],s659[1]};
    CLA_2 KS_681(s681, c681, in681_1, in681_2);
    wire[0:0] s682, in682_1, in682_2;
    wire c682;
    assign in682_1 = {s658[0]};
    assign in682_2 = {s659[0]};
    Full_Adder KS_682(s682, c682, in682_1, in682_2, s657[0]);
    wire[3:0] s683, in683_1, in683_2;
    wire c683;
    assign in683_1 = {pp36[51],pp33[55],pp30[59],pp29[61]};
    assign in683_2 = {pp37[50],pp34[54],pp31[58],pp30[60]};
    CLA_4 KS_683(s683, c683, in683_1, in683_2);
    wire[3:0] s684, in684_1, in684_2;
    wire c684;
    assign in684_1 = {pp38[49],pp35[53],pp32[57],pp31[59]};
    assign in684_2 = {pp39[48],pp36[52],pp33[56],pp32[58]};
    CLA_4 KS_684(s684, c684, in684_1, in684_2);
    wire[3:0] s685, in685_1, in685_2;
    wire c685;
    assign in685_1 = {pp40[47],pp37[51],pp34[55],pp33[57]};
    assign in685_2 = {pp41[46],pp38[50],pp35[54],pp34[56]};
    CLA_4 KS_685(s685, c685, in685_1, in685_2);
    wire[3:0] s686, in686_1, in686_2;
    wire c686;
    assign in686_1 = {pp42[45],pp39[49],pp36[53],pp35[55]};
    assign in686_2 = {pp43[44],pp40[48],pp37[52],pp36[54]};
    CLA_4 KS_686(s686, c686, in686_1, in686_2);
    wire[3:0] s687, in687_1, in687_2;
    wire c687;
    assign in687_1 = {pp44[43],pp41[47],pp38[51],pp37[53]};
    assign in687_2 = {pp45[42],pp42[46],pp39[50],pp38[52]};
    CLA_4 KS_687(s687, c687, in687_1, in687_2);
    wire[3:0] s688, in688_1, in688_2;
    wire c688;
    assign in688_1 = {pp46[41],pp43[45],pp40[49],pp39[51]};
    assign in688_2 = {pp47[40],pp44[44],pp41[48],pp40[50]};
    CLA_4 KS_688(s688, c688, in688_1, in688_2);
    wire[3:0] s689, in689_1, in689_2;
    wire c689;
    assign in689_1 = {pp48[39],pp45[43],pp42[47],pp41[49]};
    assign in689_2 = {pp49[38],pp46[42],pp43[46],pp42[48]};
    CLA_4 KS_689(s689, c689, in689_1, in689_2);
    wire[3:0] s690, in690_1, in690_2;
    wire c690;
    assign in690_1 = {pp50[37],pp47[41],pp44[45],pp43[47]};
    assign in690_2 = {pp51[36],pp48[40],pp45[44],pp44[46]};
    CLA_4 KS_690(s690, c690, in690_1, in690_2);
    wire[3:0] s691, in691_1, in691_2;
    wire c691;
    assign in691_1 = {pp52[35],pp49[39],pp46[43],pp45[45]};
    assign in691_2 = {pp53[34],pp50[38],pp47[42],pp46[44]};
    CLA_4 KS_691(s691, c691, in691_1, in691_2);
    wire[3:0] s692, in692_1, in692_2;
    wire c692;
    assign in692_1 = {pp54[33],pp51[37],pp48[41],pp47[43]};
    assign in692_2 = {pp55[32],pp52[36],pp49[40],pp48[42]};
    CLA_4 KS_692(s692, c692, in692_1, in692_2);
    wire[3:0] s693, in693_1, in693_2;
    wire c693;
    assign in693_1 = {pp56[31],pp53[35],pp50[39],pp49[41]};
    assign in693_2 = {pp57[30],pp54[34],pp51[38],pp50[40]};
    CLA_4 KS_693(s693, c693, in693_1, in693_2);
    wire[3:0] s694, in694_1, in694_2;
    wire c694;
    assign in694_1 = {pp58[29],pp55[33],pp52[37],pp51[39]};
    assign in694_2 = {pp59[28],pp56[32],pp53[36],pp52[38]};
    CLA_4 KS_694(s694, c694, in694_1, in694_2);
    wire[3:0] s695, in695_1, in695_2;
    wire c695;
    assign in695_1 = {pp60[27],pp57[31],pp54[35],pp53[37]};
    assign in695_2 = {pp61[26],pp58[30],pp55[34],pp54[36]};
    CLA_4 KS_695(s695, c695, in695_1, in695_2);
    wire[3:0] s696, in696_1, in696_2;
    wire c696;
    assign in696_1 = {pp62[25],pp59[29],pp56[33],pp55[35]};
    assign in696_2 = {pp63[24],pp60[28],pp57[32],pp56[34]};
    CLA_4 KS_696(s696, c696, in696_1, in696_2);
    wire[3:0] s697, in697_1, in697_2;
    wire c697;
    assign in697_1 = {s292[1],pp61[27],pp58[31],pp57[33]};
    assign in697_2 = {s293[1],pp62[26],pp59[30],pp58[32]};
    CLA_4 KS_697(s697, c697, in697_1, in697_2);
    wire[0:0] s698, in698_1, in698_2;
    wire c698;
    assign in698_1 = {s294[1]};
    assign in698_2 = {c295};
    Half_Adder KS_698(s698, c698, in698_1, in698_2);
    wire[3:0] s699, in699_1, in699_2;
    wire c699;
    assign in699_1 = {s296[1],pp63[25],pp60[29],pp59[31]};
    assign in699_2 = {c297,s292[2],pp61[28],pp60[30]};
    CLA_4 KS_699(s699, c699, in699_1, in699_2);
    wire[0:0] s700, in700_1, in700_2;
    wire c700;
    assign in700_1 = {s298[1]};
    assign in700_2 = {c299};
    Half_Adder KS_700(s700, c700, in700_1, in700_2);
    wire[1:0] s701, in701_1, in701_2;
    wire c701;
    assign in701_1 = {s300[1],s293[2]};
    assign in701_2 = {c653,c294};
    CLA_2 KS_701(s701, c701, in701_1, in701_2);
    wire[0:0] s702, in702_1, in702_2;
    wire c702;
    assign in702_1 = {c654};
    assign in702_2 = {c655};
    Half_Adder KS_702(s702, c702, in702_1, in702_2);
    wire[2:0] s703, in703_1, in703_2;
    wire c703;
    assign in703_1 = {c656,s296[2],pp62[27]};
    assign in703_2 = {c657,c298,pp63[26]};
    CLA_3 KS_703(s703, c703, in703_1, in703_2);
    wire[0:0] s704, in704_1, in704_2;
    wire c704;
    assign in704_1 = {c658};
    assign in704_2 = {c659};
    Half_Adder KS_704(s704, c704, in704_1, in704_2);
    wire[1:0] s705, in705_1, in705_2;
    wire c705;
    assign in705_1 = {c660,s300[2]};
    assign in705_2 = {c661,s683[1]};
    CLA_2 KS_705(s705, c705, in705_1, in705_2);
    wire[0:0] s706, in706_1, in706_2;
    wire c706;
    assign in706_1 = {c662};
    assign in706_2 = {c663};
    Half_Adder KS_706(s706, c706, in706_1, in706_2);
    wire[3:0] s707, in707_1, in707_2;
    wire c707;
    assign in707_1 = {c664,s684[1],s292[3],pp61[29]};
    assign in707_2 = {c665,s685[1],c293,pp62[28]};
    CLA_4 KS_707(s707, c707, in707_1, in707_2);
    wire[0:0] s708, in708_1, in708_2;
    wire c708;
    assign in708_1 = {c666};
    assign in708_2 = {c667};
    Half_Adder KS_708(s708, c708, in708_1, in708_2);
    wire[1:0] s709, in709_1, in709_2;
    wire c709;
    assign in709_1 = {c671,s686[1]};
    assign in709_2 = {c679,s687[1]};
    CLA_2 KS_709(s709, c709, in709_1, in709_2);
    wire[0:0] s710, in710_1, in710_2;
    wire c710;
    assign in710_1 = {s683[0]};
    assign in710_2 = {s684[0]};
    Half_Adder KS_710(s710, c710, in710_1, in710_2);
    wire[2:0] s711, in711_1, in711_2;
    wire c711;
    assign in711_1 = {s685[0],s688[1],s296[3]};
    assign in711_2 = {s686[0],s689[1],c300};
    CLA_3 KS_711(s711, c711, in711_1, in711_2);
    wire[0:0] s712, in712_1, in712_2;
    wire c712;
    assign in712_1 = {s688[0]};
    assign in712_2 = {s689[0]};
    Full_Adder KS_712(s712, c712, in712_1, in712_2, s687[0]);
    wire[3:0] s713, in713_1, in713_2;
    wire c713;
    assign in713_1 = {pp28[63],pp29[63],pp30[63],pp31[63]};
    assign in713_2 = {pp29[62],pp30[62],pp31[62],pp32[62]};
    CLA_4 KS_713(s713, c713, in713_1, in713_2);
    wire[3:0] s714, in714_1, in714_2;
    wire c714;
    assign in714_1 = {pp30[61],pp31[61],pp32[61],pp33[61]};
    assign in714_2 = {pp31[60],pp32[60],pp33[60],pp34[60]};
    CLA_4 KS_714(s714, c714, in714_1, in714_2);
    wire[3:0] s715, in715_1, in715_2;
    wire c715;
    assign in715_1 = {pp32[59],pp33[59],pp34[59],pp35[59]};
    assign in715_2 = {pp33[58],pp34[58],pp35[58],pp36[58]};
    CLA_4 KS_715(s715, c715, in715_1, in715_2);
    wire[3:0] s716, in716_1, in716_2;
    wire c716;
    assign in716_1 = {pp34[57],pp35[57],pp36[57],pp37[57]};
    assign in716_2 = {pp35[56],pp36[56],pp37[56],pp38[56]};
    CLA_4 KS_716(s716, c716, in716_1, in716_2);
    wire[3:0] s717, in717_1, in717_2;
    wire c717;
    assign in717_1 = {pp36[55],pp37[55],pp38[55],pp39[55]};
    assign in717_2 = {pp37[54],pp38[54],pp39[54],pp40[54]};
    CLA_4 KS_717(s717, c717, in717_1, in717_2);
    wire[3:0] s718, in718_1, in718_2;
    wire c718;
    assign in718_1 = {pp38[53],pp39[53],pp40[53],pp41[53]};
    assign in718_2 = {pp39[52],pp40[52],pp41[52],pp42[52]};
    CLA_4 KS_718(s718, c718, in718_1, in718_2);
    wire[3:0] s719, in719_1, in719_2;
    wire c719;
    assign in719_1 = {pp40[51],pp41[51],pp42[51],pp43[51]};
    assign in719_2 = {pp41[50],pp42[50],pp43[50],pp44[50]};
    CLA_4 KS_719(s719, c719, in719_1, in719_2);
    wire[3:0] s720, in720_1, in720_2;
    wire c720;
    assign in720_1 = {pp42[49],pp43[49],pp44[49],pp45[49]};
    assign in720_2 = {pp43[48],pp44[48],pp45[48],pp46[48]};
    CLA_4 KS_720(s720, c720, in720_1, in720_2);
    wire[3:0] s721, in721_1, in721_2;
    wire c721;
    assign in721_1 = {pp44[47],pp45[47],pp46[47],pp47[47]};
    assign in721_2 = {pp45[46],pp46[46],pp47[46],pp48[46]};
    CLA_4 KS_721(s721, c721, in721_1, in721_2);
    wire[3:0] s722, in722_1, in722_2;
    wire c722;
    assign in722_1 = {pp46[45],pp47[45],pp48[45],pp49[45]};
    assign in722_2 = {pp47[44],pp48[44],pp49[44],pp50[44]};
    CLA_4 KS_722(s722, c722, in722_1, in722_2);
    wire[3:0] s723, in723_1, in723_2;
    wire c723;
    assign in723_1 = {pp48[43],pp49[43],pp50[43],pp51[43]};
    assign in723_2 = {pp49[42],pp50[42],pp51[42],pp52[42]};
    CLA_4 KS_723(s723, c723, in723_1, in723_2);
    wire[2:0] s724, in724_1, in724_2;
    wire c724;
    assign in724_1 = {pp50[41],pp51[41],pp52[41]};
    assign in724_2 = {pp51[40],pp52[40],pp53[40]};
    CLA_3 KS_724(s724, c724, in724_1, in724_2);
    wire[1:0] s725, in725_1, in725_2;
    wire c725;
    assign in725_1 = {pp52[39],pp53[39]};
    assign in725_2 = {pp53[38],pp54[38]};
    CLA_2 KS_725(s725, c725, in725_1, in725_2);
    wire[0:0] s726, in726_1, in726_2;
    wire c726;
    assign in726_1 = {pp54[37]};
    assign in726_2 = {pp55[36]};
    Half_Adder KS_726(s726, c726, in726_1, in726_2);
    wire[3:0] s727, in727_1, in727_2;
    wire c727;
    assign in727_1 = {pp56[35],pp55[37],pp54[39],pp53[41]};
    assign in727_2 = {pp57[34],pp56[36],pp55[38],pp54[40]};
    CLA_4 KS_727(s727, c727, in727_1, in727_2);
    wire[0:0] s728, in728_1, in728_2;
    wire c728;
    assign in728_1 = {pp58[33]};
    assign in728_2 = {pp59[32]};
    Half_Adder KS_728(s728, c728, in728_1, in728_2);
    wire[1:0] s729, in729_1, in729_2;
    wire c729;
    assign in729_1 = {pp60[31],pp57[35]};
    assign in729_2 = {pp61[30],pp58[34]};
    CLA_2 KS_729(s729, c729, in729_1, in729_2);
    wire[0:0] s730, in730_1, in730_2;
    wire c730;
    assign in730_1 = {pp62[29]};
    assign in730_2 = {pp63[28]};
    Half_Adder KS_730(s730, c730, in730_1, in730_2);
    wire[2:0] s731, in731_1, in731_2;
    wire c731;
    assign in731_1 = {c301,pp59[33],pp56[37]};
    assign in731_2 = {c683,pp60[32],pp57[36]};
    CLA_3 KS_731(s731, c731, in731_1, in731_2);
    wire[0:0] s732, in732_1, in732_2;
    wire c732;
    assign in732_1 = {c684};
    assign in732_2 = {c685};
    Half_Adder KS_732(s732, c732, in732_1, in732_2);
    wire[1:0] s733, in733_1, in733_2;
    wire c733;
    assign in733_1 = {c686,pp61[31]};
    assign in733_2 = {c687,pp62[30]};
    CLA_2 KS_733(s733, c733, in733_1, in733_2);
    wire[0:0] s734, in734_1, in734_2;
    wire c734;
    assign in734_1 = {c688};
    assign in734_2 = {c689};
    Half_Adder KS_734(s734, c734, in734_1, in734_2);
    wire[3:0] s735, in735_1, in735_2;
    wire c735;
    assign in735_1 = {c690,pp63[29],pp58[35],pp55[39]};
    assign in735_2 = {c691,s713[1],pp59[34],pp56[38]};
    CLA_4 KS_735(s735, c735, in735_1, in735_2);
    wire[0:0] s736, in736_1, in736_2;
    wire c736;
    assign in736_1 = {c692};
    assign in736_2 = {c693};
    Half_Adder KS_736(s736, c736, in736_1, in736_2);
    wire[1:0] s737, in737_1, in737_2;
    wire c737;
    assign in737_1 = {c694,s714[1]};
    assign in737_2 = {c695,s715[1]};
    CLA_2 KS_737(s737, c737, in737_1, in737_2);
    wire[0:0] s738, in738_1, in738_2;
    wire c738;
    assign in738_1 = {c696};
    assign in738_2 = {c697};
    Half_Adder KS_738(s738, c738, in738_1, in738_2);
    wire[2:0] s739, in739_1, in739_2;
    wire c739;
    assign in739_1 = {c699,s716[1],pp60[33]};
    assign in739_2 = {c707,s717[1],pp61[32]};
    CLA_3 KS_739(s739, c739, in739_1, in739_2);
    wire[0:0] s740, in740_1, in740_2;
    wire c740;
    assign in740_1 = {s713[0]};
    assign in740_2 = {s714[0]};
    Half_Adder KS_740(s740, c740, in740_1, in740_2);
    wire[1:0] s741, in741_1, in741_2;
    wire c741;
    assign in741_1 = {s715[0],s718[1]};
    assign in741_2 = {s716[0],s719[1]};
    CLA_2 KS_741(s741, c741, in741_1, in741_2);
    wire[0:0] s742, in742_1, in742_2;
    wire c742;
    assign in742_1 = {s718[0]};
    assign in742_2 = {s719[0]};
    Full_Adder KS_742(s742, c742, in742_1, in742_2, s717[0]);
    wire[3:0] s743, in743_1, in743_2;
    wire c743;
    assign in743_1 = {pp32[63],pp33[63],pp34[63],pp35[63]};
    assign in743_2 = {pp33[62],pp34[62],pp35[62],pp36[62]};
    CLA_4 KS_743(s743, c743, in743_1, in743_2);
    wire[3:0] s744, in744_1, in744_2;
    wire c744;
    assign in744_1 = {pp34[61],pp35[61],pp36[61],pp37[61]};
    assign in744_2 = {pp35[60],pp36[60],pp37[60],pp38[60]};
    CLA_4 KS_744(s744, c744, in744_1, in744_2);
    wire[3:0] s745, in745_1, in745_2;
    wire c745;
    assign in745_1 = {pp36[59],pp37[59],pp38[59],pp39[59]};
    assign in745_2 = {pp37[58],pp38[58],pp39[58],pp40[58]};
    CLA_4 KS_745(s745, c745, in745_1, in745_2);
    wire[3:0] s746, in746_1, in746_2;
    wire c746;
    assign in746_1 = {pp38[57],pp39[57],pp40[57],pp41[57]};
    assign in746_2 = {pp39[56],pp40[56],pp41[56],pp42[56]};
    CLA_4 KS_746(s746, c746, in746_1, in746_2);
    wire[3:0] s747, in747_1, in747_2;
    wire c747;
    assign in747_1 = {pp40[55],pp41[55],pp42[55],pp43[55]};
    assign in747_2 = {pp41[54],pp42[54],pp43[54],pp44[54]};
    CLA_4 KS_747(s747, c747, in747_1, in747_2);
    wire[3:0] s748, in748_1, in748_2;
    wire c748;
    assign in748_1 = {pp42[53],pp43[53],pp44[53],pp45[53]};
    assign in748_2 = {pp43[52],pp44[52],pp45[52],pp46[52]};
    CLA_4 KS_748(s748, c748, in748_1, in748_2);
    wire[3:0] s749, in749_1, in749_2;
    wire c749;
    assign in749_1 = {pp44[51],pp45[51],pp46[51],pp47[51]};
    assign in749_2 = {pp45[50],pp46[50],pp47[50],pp48[50]};
    CLA_4 KS_749(s749, c749, in749_1, in749_2);
    wire[2:0] s750, in750_1, in750_2;
    wire c750;
    assign in750_1 = {pp46[49],pp47[49],pp48[49]};
    assign in750_2 = {pp47[48],pp48[48],pp49[48]};
    CLA_3 KS_750(s750, c750, in750_1, in750_2);
    wire[1:0] s751, in751_1, in751_2;
    wire c751;
    assign in751_1 = {pp48[47],pp49[47]};
    assign in751_2 = {pp49[46],pp50[46]};
    CLA_2 KS_751(s751, c751, in751_1, in751_2);
    wire[0:0] s752, in752_1, in752_2;
    wire c752;
    assign in752_1 = {pp50[45]};
    assign in752_2 = {pp51[44]};
    Half_Adder KS_752(s752, c752, in752_1, in752_2);
    wire[3:0] s753, in753_1, in753_2;
    wire c753;
    assign in753_1 = {pp52[43],pp51[45],pp50[47],pp49[49]};
    assign in753_2 = {pp53[42],pp52[44],pp51[46],pp50[48]};
    CLA_4 KS_753(s753, c753, in753_1, in753_2);
    wire[0:0] s754, in754_1, in754_2;
    wire c754;
    assign in754_1 = {pp54[41]};
    assign in754_2 = {pp55[40]};
    Half_Adder KS_754(s754, c754, in754_1, in754_2);
    wire[1:0] s755, in755_1, in755_2;
    wire c755;
    assign in755_1 = {pp56[39],pp53[43]};
    assign in755_2 = {pp57[38],pp54[42]};
    CLA_2 KS_755(s755, c755, in755_1, in755_2);
    wire[0:0] s756, in756_1, in756_2;
    wire c756;
    assign in756_1 = {pp58[37]};
    assign in756_2 = {pp59[36]};
    Half_Adder KS_756(s756, c756, in756_1, in756_2);
    wire[2:0] s757, in757_1, in757_2;
    wire c757;
    assign in757_1 = {pp60[35],pp55[41],pp52[45]};
    assign in757_2 = {pp61[34],pp56[40],pp53[44]};
    CLA_3 KS_757(s757, c757, in757_1, in757_2);
    wire[0:0] s758, in758_1, in758_2;
    wire c758;
    assign in758_1 = {pp62[33]};
    assign in758_2 = {pp63[32]};
    Half_Adder KS_758(s758, c758, in758_1, in758_2);
    wire[1:0] s759, in759_1, in759_2;
    wire c759;
    assign in759_1 = {c713,pp57[39]};
    assign in759_2 = {c714,pp58[38]};
    CLA_2 KS_759(s759, c759, in759_1, in759_2);
    wire[0:0] s760, in760_1, in760_2;
    wire c760;
    assign in760_1 = {c715};
    assign in760_2 = {c716};
    Half_Adder KS_760(s760, c760, in760_1, in760_2);
    wire[3:0] s761, in761_1, in761_2;
    wire c761;
    assign in761_1 = {c717,pp59[37],pp54[43],pp51[47]};
    assign in761_2 = {c718,pp60[36],pp55[42],pp52[46]};
    CLA_4 KS_761(s761, c761, in761_1, in761_2);
    wire[0:0] s762, in762_1, in762_2;
    wire c762;
    assign in762_1 = {c719};
    assign in762_2 = {c720};
    Half_Adder KS_762(s762, c762, in762_1, in762_2);
    wire[1:0] s763, in763_1, in763_2;
    wire c763;
    assign in763_1 = {c722,pp61[35]};
    assign in763_2 = {c723,pp62[34]};
    CLA_2_c KS_763(s763, c763, in763_1, in763_2, c721);
    wire[3:0] s764, in764_1, in764_2;
    wire c764;
    assign in764_1 = {pp36[63],pp37[63],pp38[63],pp39[63]};
    assign in764_2 = {pp37[62],pp38[62],pp39[62],pp40[62]};
    CLA_4 KS_764(s764, c764, in764_1, in764_2);
    wire[3:0] s765, in765_1, in765_2;
    wire c765;
    assign in765_1 = {pp38[61],pp39[61],pp40[61],pp41[61]};
    assign in765_2 = {pp39[60],pp40[60],pp41[60],pp42[60]};
    CLA_4 KS_765(s765, c765, in765_1, in765_2);
    wire[3:0] s766, in766_1, in766_2;
    wire c766;
    assign in766_1 = {pp40[59],pp41[59],pp42[59],pp43[59]};
    assign in766_2 = {pp41[58],pp42[58],pp43[58],pp44[58]};
    CLA_4 KS_766(s766, c766, in766_1, in766_2);
    wire[2:0] s767, in767_1, in767_2;
    wire c767;
    assign in767_1 = {pp42[57],pp43[57],pp44[57]};
    assign in767_2 = {pp43[56],pp44[56],pp45[56]};
    CLA_3 KS_767(s767, c767, in767_1, in767_2);
    wire[1:0] s768, in768_1, in768_2;
    wire c768;
    assign in768_1 = {pp44[55],pp45[55]};
    assign in768_2 = {pp45[54],pp46[54]};
    CLA_2 KS_768(s768, c768, in768_1, in768_2);
    wire[0:0] s769, in769_1, in769_2;
    wire c769;
    assign in769_1 = {pp46[53]};
    assign in769_2 = {pp47[52]};
    Half_Adder KS_769(s769, c769, in769_1, in769_2);
    wire[3:0] s770, in770_1, in770_2;
    wire c770;
    assign in770_1 = {pp48[51],pp47[53],pp46[55],pp45[57]};
    assign in770_2 = {pp49[50],pp48[52],pp47[54],pp46[56]};
    CLA_4 KS_770(s770, c770, in770_1, in770_2);
    wire[0:0] s771, in771_1, in771_2;
    wire c771;
    assign in771_1 = {pp50[49]};
    assign in771_2 = {pp51[48]};
    Half_Adder KS_771(s771, c771, in771_1, in771_2);
    wire[1:0] s772, in772_1, in772_2;
    wire c772;
    assign in772_1 = {pp52[47],pp49[51]};
    assign in772_2 = {pp53[46],pp50[50]};
    CLA_2 KS_772(s772, c772, in772_1, in772_2);
    wire[0:0] s773, in773_1, in773_2;
    wire c773;
    assign in773_1 = {pp54[45]};
    assign in773_2 = {pp55[44]};
    Half_Adder KS_773(s773, c773, in773_1, in773_2);
    wire[2:0] s774, in774_1, in774_2;
    wire c774;
    assign in774_1 = {pp56[43],pp51[49],pp48[53]};
    assign in774_2 = {pp57[42],pp52[48],pp49[52]};
    CLA_3 KS_774(s774, c774, in774_1, in774_2);
    wire[0:0] s775, in775_1, in775_2;
    wire c775;
    assign in775_1 = {pp58[41]};
    assign in775_2 = {pp59[40]};
    Half_Adder KS_775(s775, c775, in775_1, in775_2);
    wire[1:0] s776, in776_1, in776_2;
    wire c776;
    assign in776_1 = {pp61[38],pp53[47]};
    assign in776_2 = {pp62[37],pp54[46]};
    CLA_2_c KS_776(s776, c776, in776_1, in776_2, pp60[39]);
    wire[1:0] s777, in777_1, in777_2;
    wire c777;
    assign in777_1 = {pp40[63],pp41[63]};
    assign in777_2 = {pp41[62],pp42[62]};
    CLA_2 KS_777(s777, c777, in777_1, in777_2);
    wire[0:0] s778, in778_1, in778_2;
    wire c778;
    assign in778_1 = {pp42[61]};
    assign in778_2 = {pp43[60]};
    Half_Adder KS_778(s778, c778, in778_1, in778_2);
    wire[2:0] s779, in779_1, in779_2;
    wire c779;
    assign in779_1 = {pp44[59],pp43[61],pp42[63]};
    assign in779_2 = {pp45[58],pp44[60],pp43[62]};
    CLA_3 KS_779(s779, c779, in779_1, in779_2);
    wire[0:0] s780, in780_1, in780_2;
    wire c780;
    assign in780_1 = {pp47[56]};
    assign in780_2 = {pp48[55]};
    Full_Adder KS_780(s780, c780, in780_1, in780_2, pp46[57]);

    /*Stage 3*/
    wire[3:0] s781, in781_1, in781_2;
    wire c781;
    assign in781_1 = {pp0[14],pp0[15],pp0[16],pp0[17]};
    assign in781_2 = {pp1[13],pp1[14],pp1[15],pp1[16]};
    CLA_4 KS_781(s781, c781, in781_1, in781_2);
    wire[3:0] s782, in782_1, in782_2;
    wire c782;
    assign in782_1 = {pp2[13],pp2[14],pp2[15],pp0[18]};
    assign in782_2 = {pp3[12],pp3[13],pp3[14],pp1[17]};
    CLA_4 KS_782(s782, c782, in782_1, in782_2);
    wire[3:0] s783, in783_1, in783_2;
    wire c783;
    assign in783_1 = {pp4[12],pp4[13],pp2[16],pp0[19]};
    assign in783_2 = {pp5[11],pp5[12],pp3[15],pp1[18]};
    CLA_4 KS_783(s783, c783, in783_1, in783_2);
    wire[3:0] s784, in784_1, in784_2;
    wire c784;
    assign in784_1 = {pp6[11],pp4[14],pp2[17],pp0[20]};
    assign in784_2 = {pp7[10],pp5[13],pp3[16],pp1[19]};
    CLA_4 KS_784(s784, c784, in784_1, in784_2);
    wire[3:0] s785, in785_1, in785_2;
    wire c785;
    assign in785_1 = {pp6[12],pp4[15],pp2[18],pp0[21]};
    assign in785_2 = {pp7[11],pp5[14],pp3[17],pp1[20]};
    CLA_4 KS_785(s785, c785, in785_1, in785_2);
    wire[3:0] s786, in786_1, in786_2;
    wire c786;
    assign in786_1 = {pp9[9],pp6[13],pp4[16],pp2[19]};
    assign in786_2 = {pp10[8],pp7[12],pp5[15],pp3[18]};
    CLA_4_c KS_786(s786, c786, in786_1, in786_2, pp8[10]);
    wire[3:0] s787, in787_1, in787_2;
    wire c787;
    assign in787_1 = {pp8[11],pp6[14],pp4[17],pp0[22]};
    assign in787_2 = {pp9[10],pp7[13],pp5[16],pp1[21]};
    CLA_4 KS_787(s787, c787, in787_1, in787_2);
    wire[3:0] s788, in788_1, in788_2;
    wire c788;
    assign in788_1 = {pp11[8],pp8[12],pp6[15],pp2[20]};
    assign in788_2 = {pp12[7],pp9[11],pp7[14],pp3[19]};
    CLA_4_c KS_788(s788, c788, in788_1, in788_2, pp10[9]);
    wire[3:0] s789, in789_1, in789_2;
    wire c789;
    assign in789_1 = {pp10[10],pp8[13],pp4[18],pp2[21]};
    assign in789_2 = {pp11[9],pp9[12],pp5[17],pp3[20]};
    CLA_4 KS_789(s789, c789, in789_1, in789_2);
    wire[3:0] s790, in790_1, in790_2;
    wire c790;
    assign in790_1 = {pp13[7],pp10[11],pp6[16],pp4[19]};
    assign in790_2 = {pp14[6],pp11[10],pp7[15],pp5[18]};
    CLA_4_c KS_790(s790, c790, in790_1, in790_2, pp12[8]);
    wire[3:0] s791, in791_1, in791_2;
    wire c791;
    assign in791_1 = {pp12[9],pp8[14],pp6[17],pp4[20]};
    assign in791_2 = {pp13[8],pp9[13],pp7[16],pp5[19]};
    CLA_4 KS_791(s791, c791, in791_1, in791_2);
    wire[3:0] s792, in792_1, in792_2;
    wire c792;
    assign in792_1 = {pp15[6],pp10[12],pp8[15],pp6[18]};
    assign in792_2 = {pp16[5],pp11[11],pp9[14],pp7[17]};
    CLA_4_c KS_792(s792, c792, in792_1, in792_2, pp14[7]);
    wire[3:0] s793, in793_1, in793_2;
    wire c793;
    assign in793_1 = {pp12[10],pp10[13],pp8[16],pp6[19]};
    assign in793_2 = {pp13[9],pp11[12],pp9[15],pp7[18]};
    CLA_4 KS_793(s793, c793, in793_1, in793_2);
    wire[3:0] s794, in794_1, in794_2;
    wire c794;
    assign in794_1 = {pp14[8],pp12[11],pp10[14],pp8[17]};
    assign in794_2 = {pp15[7],pp13[10],pp11[13],pp9[16]};
    CLA_4 KS_794(s794, c794, in794_1, in794_2);
    wire[3:0] s795, in795_1, in795_2;
    wire c795;
    assign in795_1 = {pp16[6],pp14[9],pp12[12],pp10[15]};
    assign in795_2 = {pp17[5],pp15[8],pp13[11],pp11[14]};
    CLA_4 KS_795(s795, c795, in795_1, in795_2);
    wire[3:0] s796, in796_1, in796_2;
    wire c796;
    assign in796_1 = {pp19[3],pp16[7],pp14[10],pp12[13]};
    assign in796_2 = {pp20[2],pp17[6],pp15[9],pp13[12]};
    CLA_4_c KS_796(s796, c796, in796_1, in796_2, pp18[4]);
    wire[3:0] s797, in797_1, in797_2;
    wire c797;
    assign in797_1 = {pp18[5],pp16[8],pp14[11],pp8[18]};
    assign in797_2 = {pp19[4],pp17[7],pp15[10],pp9[17]};
    CLA_4 KS_797(s797, c797, in797_1, in797_2);
    wire[3:0] s798, in798_1, in798_2;
    wire c798;
    assign in798_1 = {pp21[2],pp18[6],pp16[9],pp10[16]};
    assign in798_2 = {pp22[1],pp19[5],pp17[8],pp11[15]};
    CLA_4_c KS_798(s798, c798, in798_1, in798_2, pp20[3]);
    wire[3:0] s799, in799_1, in799_2;
    wire c799;
    assign in799_1 = {pp20[4],pp18[7],pp12[14],pp11[16]};
    assign in799_2 = {pp21[3],pp19[6],pp13[13],pp12[15]};
    CLA_4 KS_799(s799, c799, in799_1, in799_2);
    wire[3:0] s800, in800_1, in800_2;
    wire c800;
    assign in800_1 = {pp23[1],pp20[5],pp14[12],pp13[14]};
    assign in800_2 = {pp24[0],pp21[4],pp15[11],pp14[13]};
    CLA_4_c KS_800(s800, c800, in800_1, in800_2, pp22[2]);
    wire[3:0] s801, in801_1, in801_2;
    wire c801;
    assign in801_1 = {pp22[3],pp16[10],pp15[12],pp13[15]};
    assign in801_2 = {pp23[2],pp17[9],pp16[11],pp14[14]};
    CLA_4 KS_801(s801, c801, in801_1, in801_2);
    wire[3:0] s802, in802_1, in802_2;
    wire c802;
    assign in802_1 = {pp25[0],pp18[8],pp17[10],pp15[13]};
    assign in802_2 = {s302[2],pp19[7],pp18[9],pp16[12]};
    CLA_4_c KS_802(s802, c802, in802_1, in802_2, pp24[1]);
    wire[3:0] s803, in803_1, in803_2;
    wire c803;
    assign in803_1 = {pp20[6],pp19[8],pp17[11],pp15[14]};
    assign in803_2 = {pp21[5],pp20[7],pp18[10],pp16[13]};
    CLA_4 KS_803(s803, c803, in803_1, in803_2);
    wire[3:0] s804, in804_1, in804_2;
    wire c804;
    assign in804_1 = {pp22[4],pp21[6],pp19[9],pp17[12]};
    assign in804_2 = {pp23[3],pp22[5],pp20[8],pp18[11]};
    CLA_4 KS_804(s804, c804, in804_1, in804_2);
    wire[3:0] s805, in805_1, in805_2;
    wire c805;
    assign in805_1 = {pp24[2],pp23[4],pp21[7],pp19[10]};
    assign in805_2 = {pp25[1],pp24[3],pp22[6],pp20[9]};
    CLA_4 KS_805(s805, c805, in805_1, in805_2);
    wire[3:0] s806, in806_1, in806_2;
    wire c806;
    assign in806_1 = {pp26[0],pp25[2],pp23[5],pp21[8]};
    assign in806_2 = {s302[3],pp26[1],pp24[4],pp22[7]};
    CLA_4 KS_806(s806, c806, in806_1, in806_2);
    wire[3:0] s807, in807_1, in807_2;
    wire c807;
    assign in807_1 = {s303[2],pp27[0],pp25[3],pp23[6]};
    assign in807_2 = {s304[1],c302,pp26[2],pp24[5]};
    CLA_4 KS_807(s807, c807, in807_1, in807_2);
    wire[3:0] s808, in808_1, in808_2;
    wire c808;
    assign in808_1 = {c793,s303[3],pp27[1],pp25[4]};
    assign in808_2 = {c794,s304[2],pp28[0],pp26[3]};
    CLA_4_c KS_808(s808, c808, in808_1, in808_2, s305[0]);
    wire[3:0] s809, in809_1, in809_2;
    wire c809;
    assign in809_1 = {s305[1],c303,pp27[2],pp17[13]};
    assign in809_2 = {s306[0],s304[3],pp28[1],pp18[12]};
    CLA_4 KS_809(s809, c809, in809_1, in809_2);
    wire[3:0] s810, in810_1, in810_2;
    wire c810;
    assign in810_1 = {s306[1],pp29[0],pp19[11],pp21[10]};
    assign in810_2 = {s307[1],c304,pp20[10],pp22[9]};
    CLA_4_c KS_810(s810, c810, in810_1, in810_2, s305[2]);
    wire[3:0] s811, in811_1, in811_2;
    wire c811;
    assign in811_1 = {s305[3],pp21[9],pp23[8],pp23[9]};
    assign in811_2 = {s306[2],pp22[8],pp24[7],pp24[8]};
    CLA_4 KS_811(s811, c811, in811_1, in811_2);
    wire[3:0] s812, in812_1, in812_2;
    wire c812;
    assign in812_1 = {s308[1],pp23[7],pp25[6],pp25[7]};
    assign in812_2 = {s309[1],pp24[6],pp26[5],pp26[6]};
    CLA_4_c KS_812(s812, c812, in812_1, in812_2, s307[2]);
    wire[3:0] s813, in813_1, in813_2;
    wire c813;
    assign in813_1 = {pp25[5],pp27[4],pp27[5],pp25[8]};
    assign in813_2 = {pp26[4],pp28[3],pp28[4],pp26[7]};
    CLA_4 KS_813(s813, c813, in813_1, in813_2);
    wire[3:0] s814, in814_1, in814_2;
    wire c814;
    assign in814_1 = {pp27[3],pp29[2],pp29[3],pp27[6]};
    assign in814_2 = {pp28[2],pp30[1],pp30[2],pp28[5]};
    CLA_4 KS_814(s814, c814, in814_1, in814_2);
    wire[3:0] s815, in815_1, in815_2;
    wire c815;
    assign in815_1 = {pp29[1],pp31[0],pp31[1],pp29[4]};
    assign in815_2 = {pp30[0],c306,pp32[0],pp30[3]};
    CLA_4 KS_815(s815, c815, in815_1, in815_2);
    wire[3:0] s816, in816_1, in816_2;
    wire c816;
    assign in816_1 = {c305,c307,c308,pp31[2]};
    assign in816_2 = {s306[3],s308[3],c309,pp32[1]};
    CLA_4 KS_816(s816, c816, in816_1, in816_2);
    wire[3:0] s817, in817_1, in817_2;
    wire c817;
    assign in817_1 = {s307[3],s309[3],s310[3],pp33[0]};
    assign in817_2 = {s308[2],s310[2],s311[3],c310};
    CLA_4 KS_817(s817, c817, in817_1, in817_2);
    wire[3:0] s818, in818_1, in818_2;
    wire c818;
    assign in818_1 = {s309[2],s311[2],s312[2],c311};
    assign in818_2 = {s310[1],s312[1],s313[2],s312[3]};
    CLA_4 KS_818(s818, c818, in818_1, in818_2);
    wire[3:0] s819, in819_1, in819_2;
    wire c819;
    assign in819_1 = {s311[1],s313[1],s314[1],s313[3]};
    assign in819_2 = {s312[0],s314[0],s315[1],s314[2]};
    CLA_4 KS_819(s819, c819, in819_1, in819_2);
    wire[3:0] s820, in820_1, in820_2;
    wire c820;
    assign in820_1 = {s313[0],s315[0],s316[1],s315[2]};
    assign in820_2 = {c803,s316[0],s317[1],s316[2]};
    CLA_4 KS_820(s820, c820, in820_1, in820_2);
    wire[0:0] s821, in821_1, in821_2;
    wire c821;
    assign in821_1 = {c804};
    assign in821_2 = {c805};
    Half_Adder KS_821(s821, c821, in821_1, in821_2);
    wire[3:0] s822, in822_1, in822_2;
    wire c822;
    assign in822_1 = {c807,s317[0],s318[0],s317[2]};
    assign in822_2 = {c808,c809,s319[0],s318[1]};
    CLA_4_c KS_822(s822, c822, in822_1, in822_2, c806);
    wire[3:0] s823, in823_1, in823_2;
    wire c823;
    assign in823_1 = {s320[1],pp27[7],pp33[2],pp33[3]};
    assign in823_2 = {s321[0],pp28[6],pp34[1],pp34[2]};
    CLA_4_c KS_823(s823, c823, in823_1, in823_2, s319[1]);
    wire[3:0] s824, in824_1, in824_2;
    wire c824;
    assign in824_1 = {pp29[5],pp35[0],pp35[1],pp35[2]};
    assign in824_2 = {pp30[4],c314,pp36[0],pp36[1]};
    CLA_4 KS_824(s824, c824, in824_1, in824_2);
    wire[3:0] s825, in825_1, in825_2;
    wire c825;
    assign in825_1 = {pp31[3],c315,c318,pp37[0]};
    assign in825_2 = {pp32[2],c316,c319,c321};
    CLA_4 KS_825(s825, c825, in825_1, in825_2);
    wire[3:0] s826, in826_1, in826_2;
    wire c826;
    assign in826_1 = {pp33[1],c317,c320,c322};
    assign in826_2 = {pp34[0],s318[3],s321[3],c323};
    CLA_4 KS_826(s826, c826, in826_1, in826_2);
    wire[3:0] s827, in827_1, in827_2;
    wire c827;
    assign in827_1 = {c312,s319[3],s322[3],s324[3]};
    assign in827_2 = {c313,s320[3],s323[3],s325[3]};
    CLA_4 KS_827(s827, c827, in827_1, in827_2);
    wire[3:0] s828, in828_1, in828_2;
    wire c828;
    assign in828_1 = {s314[3],s321[2],s324[2],s326[3]};
    assign in828_2 = {s315[3],s322[2],s325[2],s327[2]};
    CLA_4 KS_828(s828, c828, in828_1, in828_2);
    wire[3:0] s829, in829_1, in829_2;
    wire c829;
    assign in829_1 = {s316[3],s323[2],s326[2],s328[2]};
    assign in829_2 = {s317[3],s324[1],s327[1],s329[2]};
    CLA_4 KS_829(s829, c829, in829_1, in829_2);
    wire[3:0] s830, in830_1, in830_2;
    wire c830;
    assign in830_1 = {s318[2],s325[1],s328[1],s330[2]};
    assign in830_2 = {s319[2],s326[1],s329[1],s331[2]};
    CLA_4 KS_830(s830, c830, in830_1, in830_2);
    wire[3:0] s831, in831_1, in831_2;
    wire c831;
    assign in831_1 = {s320[2],s327[0],s330[1],s332[2]};
    assign in831_2 = {s321[1],s328[0],s331[1],s333[2]};
    CLA_4 KS_831(s831, c831, in831_1, in831_2);
    wire[3:0] s832, in832_1, in832_2;
    wire c832;
    assign in832_1 = {s322[1],s329[0],s332[1],s334[1]};
    assign in832_2 = {s323[1],s330[0],s333[1],s335[1]};
    CLA_4 KS_832(s832, c832, in832_1, in832_2);
    wire[0:0] s833, in833_1, in833_2;
    wire c833;
    assign in833_1 = {s324[0]};
    assign in833_2 = {s325[0]};
    Half_Adder KS_833(s833, c833, in833_1, in833_2);
    wire[1:0] s834, in834_1, in834_2;
    wire c834;
    assign in834_1 = {s326[0],s331[0]};
    assign in834_2 = {c813,s332[0]};
    CLA_2 KS_834(s834, c834, in834_1, in834_2);
    wire[0:0] s835, in835_1, in835_2;
    wire c835;
    assign in835_1 = {c814};
    assign in835_2 = {c815};
    Half_Adder KS_835(s835, c835, in835_1, in835_2);
    wire[3:0] s836, in836_1, in836_2;
    wire c836;
    assign in836_1 = {c816,s333[0],s334[0],s336[1]};
    assign in836_2 = {c817,s823[2],s335[0],s337[0]};
    CLA_4 KS_836(s836, c836, in836_1, in836_2);
    wire[0:0] s837, in837_1, in837_2;
    wire c837;
    assign in837_1 = {c818};
    assign in837_2 = {c819};
    Half_Adder KS_837(s837, c837, in837_1, in837_2);
    wire[1:0] s838, in838_1, in838_2;
    wire c838;
    assign in838_1 = {c820,s824[1]};
    assign in838_2 = {c822,s825[1]};
    CLA_2 KS_838(s838, c838, in838_1, in838_2);
    wire[0:0] s839, in839_1, in839_2;
    wire c839;
    assign in839_1 = {s824[0]};
    assign in839_2 = {s825[0]};
    Full_Adder KS_839(s839, c839, in839_1, in839_2, s823[1]);
    wire[3:0] s840, in840_1, in840_2;
    wire c840;
    assign in840_1 = {pp37[1],c332,s2[1],s4[0]};
    assign in840_2 = {pp38[0],c333,s3[0],c337};
    CLA_4 KS_840(s840, c840, in840_1, in840_2);
    wire[3:0] s841, in841_1, in841_2;
    wire c841;
    assign in841_1 = {s1[0],s334[3],c334,c338};
    assign in841_2 = {c324,s335[3],c335,c339};
    CLA_4 KS_841(s841, c841, in841_1, in841_2);
    wire[3:0] s842, in842_1, in842_2;
    wire c842;
    assign in842_1 = {c325,s336[3],c336,c340};
    assign in842_2 = {c326,s337[2],s337[3],s341[3]};
    CLA_4 KS_842(s842, c842, in842_1, in842_2);
    wire[3:0] s843, in843_1, in843_2;
    wire c843;
    assign in843_1 = {s327[3],s338[2],s338[3],s342[3]};
    assign in843_2 = {s328[3],s339[2],s339[3],s343[3]};
    CLA_4 KS_843(s843, c843, in843_1, in843_2);
    wire[3:0] s844, in844_1, in844_2;
    wire c844;
    assign in844_1 = {s329[3],s340[2],s340[3],s344[2]};
    assign in844_2 = {s330[3],s341[1],s341[2],s345[2]};
    CLA_4 KS_844(s844, c844, in844_1, in844_2);
    wire[3:0] s845, in845_1, in845_2;
    wire c845;
    assign in845_1 = {s331[3],s342[1],s342[2],s346[2]};
    assign in845_2 = {s332[3],s343[1],s343[2],s347[2]};
    CLA_4 KS_845(s845, c845, in845_1, in845_2);
    wire[3:0] s846, in846_1, in846_2;
    wire c846;
    assign in846_1 = {s333[3],s344[0],s344[1],s348[2]};
    assign in846_2 = {s334[2],s345[0],s345[1],s349[2]};
    CLA_4 KS_846(s846, c846, in846_1, in846_2);
    wire[3:0] s847, in847_1, in847_2;
    wire c847;
    assign in847_1 = {s335[2],s346[0],s346[1],s350[2]};
    assign in847_2 = {s336[2],s347[0],s347[1],s351[2]};
    CLA_4 KS_847(s847, c847, in847_1, in847_2);
    wire[3:0] s848, in848_1, in848_2;
    wire c848;
    assign in848_1 = {s337[1],s348[0],s348[1],s352[2]};
    assign in848_2 = {s338[1],s349[0],s349[1],s353[2]};
    CLA_4 KS_848(s848, c848, in848_1, in848_2);
    wire[3:0] s849, in849_1, in849_2;
    wire c849;
    assign in849_1 = {s339[1],s350[0],s350[1],s354[2]};
    assign in849_2 = {s340[1],s351[0],s351[1],s355[0]};
    CLA_4 KS_849(s849, c849, in849_1, in849_2);
    wire[0:0] s850, in850_1, in850_2;
    wire c850;
    assign in850_1 = {s341[0]};
    assign in850_2 = {s342[0]};
    Half_Adder KS_850(s850, c850, in850_1, in850_2);
    wire[1:0] s851, in851_1, in851_2;
    wire c851;
    assign in851_1 = {s343[0],s352[0]};
    assign in851_2 = {c824,s353[0]};
    CLA_2 KS_851(s851, c851, in851_1, in851_2);
    wire[0:0] s852, in852_1, in852_2;
    wire c852;
    assign in852_1 = {c825};
    assign in852_2 = {c826};
    Half_Adder KS_852(s852, c852, in852_1, in852_2);
    wire[2:0] s853, in853_1, in853_2;
    wire c853;
    assign in853_1 = {c827,s354[0],s352[1]};
    assign in853_2 = {c828,s840[1],s353[1]};
    CLA_3 KS_853(s853, c853, in853_1, in853_2);
    wire[0:0] s854, in854_1, in854_2;
    wire c854;
    assign in854_1 = {c829};
    assign in854_2 = {c830};
    Half_Adder KS_854(s854, c854, in854_1, in854_2);
    wire[1:0] s855, in855_1, in855_2;
    wire c855;
    assign in855_1 = {c831,s841[1]};
    assign in855_2 = {c832,s842[1]};
    CLA_2 KS_855(s855, c855, in855_1, in855_2);
    wire[0:0] s856, in856_1, in856_2;
    wire c856;
    assign in856_1 = {c836};
    assign in856_2 = {s840[0]};
    Half_Adder KS_856(s856, c856, in856_1, in856_2);
    wire[3:0] s857, in857_1, in857_2;
    wire c857;
    assign in857_1 = {s842[0],s843[1],s354[1],s356[0]};
    assign in857_2 = {s843[0],s844[1],s840[2],s357[0]};
    CLA_4_c KS_857(s857, c857, in857_1, in857_2, s841[0]);
    wire[3:0] s858, in858_1, in858_2;
    wire c858;
    assign in858_1 = {s4[1],s357[2],s357[3],s12[0]};
    assign in858_2 = {s5[0],s358[2],s358[3],c355};
    CLA_4 KS_858(s858, c858, in858_1, in858_2);
    wire[3:0] s859, in859_1, in859_2;
    wire c859;
    assign in859_1 = {s6[0],s359[1],s359[2],c356};
    assign in859_2 = {c341,s360[1],s360[2],c357};
    CLA_4 KS_859(s859, c859, in859_1, in859_2);
    wire[3:0] s860, in860_1, in860_2;
    wire c860;
    assign in860_1 = {c342,s361[0],s361[1],c358};
    assign in860_2 = {c343,s362[0],s362[1],s359[3]};
    CLA_4 KS_860(s860, c860, in860_1, in860_2);
    wire[3:0] s861, in861_1, in861_2;
    wire c861;
    assign in861_1 = {s344[3],s363[0],s363[1],s360[3]};
    assign in861_2 = {s345[3],s364[0],s364[1],s361[2]};
    CLA_4 KS_861(s861, c861, in861_1, in861_2);
    wire[3:0] s862, in862_1, in862_2;
    wire c862;
    assign in862_1 = {s346[3],s365[0],s365[1],s362[2]};
    assign in862_2 = {s347[3],s366[0],s366[1],s363[2]};
    CLA_4 KS_862(s862, c862, in862_1, in862_2);
    wire[3:0] s863, in863_1, in863_2;
    wire c863;
    assign in863_1 = {s348[3],s367[0],s367[1],s364[2]};
    assign in863_2 = {s349[3],s368[0],s368[1],s365[2]};
    CLA_4 KS_863(s863, c863, in863_1, in863_2);
    wire[3:0] s864, in864_1, in864_2;
    wire c864;
    assign in864_1 = {s350[3],s369[0],s369[1],s366[2]};
    assign in864_2 = {s351[3],s370[0],s370[1],s367[2]};
    CLA_4 KS_864(s864, c864, in864_1, in864_2);
    wire[3:0] s865, in865_1, in865_2;
    wire c865;
    assign in865_1 = {s352[3],s371[0],c371,s368[2]};
    assign in865_2 = {s353[3],s372[0],s372[1],s369[2]};
    CLA_4 KS_865(s865, c865, in865_1, in865_2);
    wire[3:0] s866, in866_1, in866_2;
    wire c866;
    assign in866_1 = {s354[3],s373[0],c373,s370[2]};
    assign in866_2 = {s355[1],s374[0],s374[1],s372[2]};
    CLA_4 KS_866(s866, c866, in866_1, in866_2);
    wire[3:0] s867, in867_1, in867_2;
    wire c867;
    assign in867_1 = {s356[1],s375[0],c375,s374[2]};
    assign in867_2 = {s357[1],s376[0],s376[1],s376[2]};
    CLA_4 KS_867(s867, c867, in867_1, in867_2);
    wire[0:0] s868, in868_1, in868_2;
    wire c868;
    assign in868_1 = {s358[1]};
    assign in868_2 = {s359[0]};
    Half_Adder KS_868(s868, c868, in868_1, in868_2);
    wire[1:0] s869, in869_1, in869_2;
    wire c869;
    assign in869_1 = {s360[0],s377[0]};
    assign in869_2 = {c840,s378[0]};
    CLA_2 KS_869(s869, c869, in869_1, in869_2);
    wire[0:0] s870, in870_1, in870_2;
    wire c870;
    assign in870_1 = {c841};
    assign in870_2 = {c842};
    Half_Adder KS_870(s870, c870, in870_1, in870_2);
    wire[2:0] s871, in871_1, in871_2;
    wire c871;
    assign in871_1 = {c843,s379[0],c377};
    assign in871_2 = {c844,s858[1],s378[1]};
    CLA_3 KS_871(s871, c871, in871_1, in871_2);
    wire[0:0] s872, in872_1, in872_2;
    wire c872;
    assign in872_1 = {c845};
    assign in872_2 = {c846};
    Half_Adder KS_872(s872, c872, in872_1, in872_2);
    wire[1:0] s873, in873_1, in873_2;
    wire c873;
    assign in873_1 = {c847,s859[1]};
    assign in873_2 = {c848,s860[1]};
    CLA_2 KS_873(s873, c873, in873_1, in873_2);
    wire[0:0] s874, in874_1, in874_2;
    wire c874;
    assign in874_1 = {c849};
    assign in874_2 = {c857};
    Half_Adder KS_874(s874, c874, in874_1, in874_2);
    wire[3:0] s875, in875_1, in875_2;
    wire c875;
    assign in875_1 = {s858[0],s861[1],c379,s378[2]};
    assign in875_2 = {s859[0],s862[1],s858[2],s380[0]};
    CLA_4 KS_875(s875, c875, in875_1, in875_2);
    wire[0:0] s876, in876_1, in876_2;
    wire c876;
    assign in876_1 = {s861[0]};
    assign in876_2 = {s862[0]};
    Full_Adder KS_876(s876, c876, in876_1, in876_2, s860[0]);
    wire[3:0] s877, in877_1, in877_2;
    wire c877;
    assign in877_1 = {s13[0],s385[0],s386[1],c380};
    assign in877_2 = {s14[0],s386[0],s387[1],c381};
    CLA_4 KS_877(s877, c877, in877_1, in877_2);
    wire[3:0] s878, in878_1, in878_2;
    wire c878;
    assign in878_1 = {s15[0],s387[0],s388[1],s382[3]};
    assign in878_2 = {s16[0],s388[0],s389[1],s383[2]};
    CLA_4 KS_878(s878, c878, in878_1, in878_2);
    wire[3:0] s879, in879_1, in879_2;
    wire c879;
    assign in879_1 = {c359,s389[0],s390[1],s384[2]};
    assign in879_2 = {c360,s390[0],s391[1],s385[2]};
    CLA_4 KS_879(s879, c879, in879_1, in879_2);
    wire[3:0] s880, in880_1, in880_2;
    wire c880;
    assign in880_1 = {s361[3],s391[0],s392[1],s386[2]};
    assign in880_2 = {s362[3],s392[0],s393[1],s387[2]};
    CLA_4 KS_880(s880, c880, in880_1, in880_2);
    wire[3:0] s881, in881_1, in881_2;
    wire c881;
    assign in881_1 = {s363[3],s393[0],s394[1],s388[2]};
    assign in881_2 = {s364[3],s394[0],s395[1],s389[2]};
    CLA_4 KS_881(s881, c881, in881_1, in881_2);
    wire[3:0] s882, in882_1, in882_2;
    wire c882;
    assign in882_1 = {s365[3],s395[0],c396,s390[2]};
    assign in882_2 = {s366[3],s396[0],s397[1],s391[2]};
    CLA_4 KS_882(s882, c882, in882_1, in882_2);
    wire[3:0] s883, in883_1, in883_2;
    wire c883;
    assign in883_1 = {s367[3],s397[0],c398,s392[2]};
    assign in883_2 = {s368[3],s398[0],s399[1],s393[2]};
    CLA_4 KS_883(s883, c883, in883_1, in883_2);
    wire[3:0] s884, in884_1, in884_2;
    wire c884;
    assign in884_1 = {s369[3],s399[0],c400,s394[2]};
    assign in884_2 = {s370[3],s400[0],s401[1],s395[2]};
    CLA_4 KS_884(s884, c884, in884_1, in884_2);
    wire[3:0] s885, in885_1, in885_2;
    wire c885;
    assign in885_1 = {s372[3],s401[0],c402,s397[2]};
    assign in885_2 = {s374[3],s402[0],s403[1],s399[2]};
    CLA_4 KS_885(s885, c885, in885_1, in885_2);
    wire[1:0] s886, in886_1, in886_2;
    wire c886;
    assign in886_1 = {s376[3],s403[0]};
    assign in886_2 = {s378[3],s404[0]};
    CLA_2 KS_886(s886, c886, in886_1, in886_2);
    wire[0:0] s887, in887_1, in887_2;
    wire c887;
    assign in887_1 = {s380[1]};
    assign in887_2 = {s381[1]};
    Half_Adder KS_887(s887, c887, in887_1, in887_2);
    wire[2:0] s888, in888_1, in888_2;
    wire c888;
    assign in888_1 = {s382[0],s405[0],c404};
    assign in888_2 = {c858,s406[0],s405[1]};
    CLA_3 KS_888(s888, c888, in888_1, in888_2);
    wire[0:0] s889, in889_1, in889_2;
    wire c889;
    assign in889_1 = {c859};
    assign in889_2 = {c860};
    Half_Adder KS_889(s889, c889, in889_1, in889_2);
    wire[1:0] s890, in890_1, in890_2;
    wire c890;
    assign in890_1 = {c861,s407[0]};
    assign in890_2 = {c862,s877[1]};
    CLA_2 KS_890(s890, c890, in890_1, in890_2);
    wire[0:0] s891, in891_1, in891_2;
    wire c891;
    assign in891_1 = {c863};
    assign in891_2 = {c864};
    Half_Adder KS_891(s891, c891, in891_1, in891_2);
    wire[3:0] s892, in892_1, in892_2;
    wire c892;
    assign in892_1 = {c865,s878[1],c406,s401[2]};
    assign in892_2 = {c866,s879[1],s407[1],s403[2]};
    CLA_4 KS_892(s892, c892, in892_1, in892_2);
    wire[0:0] s893, in893_1, in893_2;
    wire c893;
    assign in893_1 = {c867};
    assign in893_2 = {c875};
    Half_Adder KS_893(s893, c893, in893_1, in893_2);
    wire[1:0] s894, in894_1, in894_2;
    wire c894;
    assign in894_1 = {s877[0],s880[1]};
    assign in894_2 = {s878[0],s881[1]};
    CLA_2 KS_894(s894, c894, in894_1, in894_2);
    wire[0:0] s895, in895_1, in895_2;
    wire c895;
    assign in895_1 = {s880[0]};
    assign in895_2 = {s881[0]};
    Full_Adder KS_895(s895, c895, in895_1, in895_2, s879[0]);
    wire[3:0] s896, in896_1, in896_2;
    wire c896;
    assign in896_1 = {s29[0],s416[0],s416[1],s408[2]};
    assign in896_2 = {s30[0],s417[0],s417[1],s409[2]};
    CLA_4 KS_896(s896, c896, in896_1, in896_2);
    wire[3:0] s897, in897_1, in897_2;
    wire c897;
    assign in897_1 = {s31[0],s418[0],s418[1],s410[2]};
    assign in897_2 = {s32[0],s419[0],s419[1],s411[2]};
    CLA_4 KS_897(s897, c897, in897_1, in897_2);
    wire[3:0] s898, in898_1, in898_2;
    wire c898;
    assign in898_1 = {c382,s420[0],s420[1],s412[2]};
    assign in898_2 = {s383[3],s421[0],s421[1],s413[2]};
    CLA_4 KS_898(s898, c898, in898_1, in898_2);
    wire[3:0] s899, in899_1, in899_2;
    wire c899;
    assign in899_1 = {s384[3],s422[0],s422[1],s414[2]};
    assign in899_2 = {s385[3],s423[0],s423[1],s415[2]};
    CLA_4 KS_899(s899, c899, in899_1, in899_2);
    wire[3:0] s900, in900_1, in900_2;
    wire c900;
    assign in900_1 = {s386[3],s424[0],c424,s416[2]};
    assign in900_2 = {s387[3],s425[0],s425[1],s417[2]};
    CLA_4 KS_900(s900, c900, in900_1, in900_2);
    wire[3:0] s901, in901_1, in901_2;
    wire c901;
    assign in901_1 = {s388[3],s426[0],c426,s418[2]};
    assign in901_2 = {s389[3],s427[0],s427[1],s419[2]};
    CLA_4 KS_901(s901, c901, in901_1, in901_2);
    wire[3:0] s902, in902_1, in902_2;
    wire c902;
    assign in902_1 = {s390[3],s428[0],c428,s420[2]};
    assign in902_2 = {s391[3],s429[0],s429[1],s421[2]};
    CLA_4 KS_902(s902, c902, in902_1, in902_2);
    wire[3:0] s903, in903_1, in903_2;
    wire c903;
    assign in903_1 = {s392[3],s430[0],c430,s422[2]};
    assign in903_2 = {s393[3],s431[0],s431[1],s423[2]};
    CLA_4 KS_903(s903, c903, in903_1, in903_2);
    wire[3:0] s904, in904_1, in904_2;
    wire c904;
    assign in904_1 = {s394[3],s432[0],c432,c425};
    assign in904_2 = {s395[3],s433[0],s433[1],s427[2]};
    CLA_4 KS_904(s904, c904, in904_1, in904_2);
    wire[3:0] s905, in905_1, in905_2;
    wire c905;
    assign in905_1 = {s397[3],s434[0],c434,c429};
    assign in905_2 = {s399[3],s435[0],s435[1],s431[2]};
    CLA_4 KS_905(s905, c905, in905_1, in905_2);
    wire[0:0] s906, in906_1, in906_2;
    wire c906;
    assign in906_1 = {s401[3]};
    assign in906_2 = {s403[3]};
    Half_Adder KS_906(s906, c906, in906_1, in906_2);
    wire[1:0] s907, in907_1, in907_2;
    wire c907;
    assign in907_1 = {c407,s436[0]};
    assign in907_2 = {c877,s437[0]};
    CLA_2 KS_907(s907, c907, in907_1, in907_2);
    wire[0:0] s908, in908_1, in908_2;
    wire c908;
    assign in908_1 = {c878};
    assign in908_2 = {c879};
    Half_Adder KS_908(s908, c908, in908_1, in908_2);
    wire[2:0] s909, in909_1, in909_2;
    wire c909;
    assign in909_1 = {c880,s438[0],c436};
    assign in909_2 = {c881,s896[1],s437[1]};
    CLA_3 KS_909(s909, c909, in909_1, in909_2);
    wire[0:0] s910, in910_1, in910_2;
    wire c910;
    assign in910_1 = {c882};
    assign in910_2 = {c883};
    Half_Adder KS_910(s910, c910, in910_1, in910_2);
    wire[1:0] s911, in911_1, in911_2;
    wire c911;
    assign in911_1 = {c884,s897[1]};
    assign in911_2 = {c885,s898[1]};
    CLA_2 KS_911(s911, c911, in911_1, in911_2);
    wire[0:0] s912, in912_1, in912_2;
    wire c912;
    assign in912_1 = {c892};
    assign in912_2 = {s896[0]};
    Half_Adder KS_912(s912, c912, in912_1, in912_2);
    wire[3:0] s913, in913_1, in913_2;
    wire c913;
    assign in913_1 = {s898[0],s899[1],c438,c433};
    assign in913_2 = {s899[0],s900[1],s896[2],s435[2]};
    CLA_4_c KS_913(s913, c913, in913_1, in913_2, s897[0]);
    wire[3:0] s914, in914_1, in914_2;
    wire c914;
    assign in914_1 = {s52[0],s447[0],s447[1],s439[2]};
    assign in914_2 = {s53[0],s448[0],s448[1],s440[2]};
    CLA_4 KS_914(s914, c914, in914_1, in914_2);
    wire[3:0] s915, in915_1, in915_2;
    wire c915;
    assign in915_1 = {s54[0],s449[0],s449[1],s441[2]};
    assign in915_2 = {s55[0],s450[0],s450[1],s442[2]};
    CLA_4 KS_915(s915, c915, in915_1, in915_2);
    wire[3:0] s916, in916_1, in916_2;
    wire c916;
    assign in916_1 = {s408[3],s451[0],s451[1],s443[2]};
    assign in916_2 = {s409[3],s452[0],s452[1],s444[2]};
    CLA_4 KS_916(s916, c916, in916_1, in916_2);
    wire[3:0] s917, in917_1, in917_2;
    wire c917;
    assign in917_1 = {s410[3],s453[0],s453[1],s445[2]};
    assign in917_2 = {s411[3],s454[0],s454[1],s446[2]};
    CLA_4 KS_917(s917, c917, in917_1, in917_2);
    wire[3:0] s918, in918_1, in918_2;
    wire c918;
    assign in918_1 = {s412[3],s455[0],c455,s447[2]};
    assign in918_2 = {s413[3],s456[0],s456[1],s448[2]};
    CLA_4 KS_918(s918, c918, in918_1, in918_2);
    wire[3:0] s919, in919_1, in919_2;
    wire c919;
    assign in919_1 = {s414[3],s457[0],c457,s449[2]};
    assign in919_2 = {s415[3],s458[0],s458[1],s450[2]};
    CLA_4 KS_919(s919, c919, in919_1, in919_2);
    wire[3:0] s920, in920_1, in920_2;
    wire c920;
    assign in920_1 = {s416[3],s459[0],c459,s451[2]};
    assign in920_2 = {s417[3],s460[0],s460[1],s452[2]};
    CLA_4 KS_920(s920, c920, in920_1, in920_2);
    wire[3:0] s921, in921_1, in921_2;
    wire c921;
    assign in921_1 = {s418[3],s461[0],c461,s453[2]};
    assign in921_2 = {s419[3],s462[0],s462[1],s454[2]};
    CLA_4 KS_921(s921, c921, in921_1, in921_2);
    wire[3:0] s922, in922_1, in922_2;
    wire c922;
    assign in922_1 = {s420[3],s463[0],c463,c456};
    assign in922_2 = {s421[3],s464[0],s464[1],s458[2]};
    CLA_4 KS_922(s922, c922, in922_1, in922_2);
    wire[3:0] s923, in923_1, in923_2;
    wire c923;
    assign in923_1 = {s422[3],s465[0],c465,c460};
    assign in923_2 = {s423[3],s466[0],s466[1],s462[2]};
    CLA_4 KS_923(s923, c923, in923_1, in923_2);
    wire[0:0] s924, in924_1, in924_2;
    wire c924;
    assign in924_1 = {c427};
    assign in924_2 = {s431[3]};
    Half_Adder KS_924(s924, c924, in924_1, in924_2);
    wire[1:0] s925, in925_1, in925_2;
    wire c925;
    assign in925_1 = {c435,s467[0]};
    assign in925_2 = {c896,s468[0]};
    CLA_2 KS_925(s925, c925, in925_1, in925_2);
    wire[0:0] s926, in926_1, in926_2;
    wire c926;
    assign in926_1 = {c897};
    assign in926_2 = {c898};
    Half_Adder KS_926(s926, c926, in926_1, in926_2);
    wire[2:0] s927, in927_1, in927_2;
    wire c927;
    assign in927_1 = {c899,s469[0],c467};
    assign in927_2 = {c900,s914[1],s468[1]};
    CLA_3 KS_927(s927, c927, in927_1, in927_2);
    wire[0:0] s928, in928_1, in928_2;
    wire c928;
    assign in928_1 = {c901};
    assign in928_2 = {c902};
    Half_Adder KS_928(s928, c928, in928_1, in928_2);
    wire[1:0] s929, in929_1, in929_2;
    wire c929;
    assign in929_1 = {c903,s915[1]};
    assign in929_2 = {c904,s916[1]};
    CLA_2 KS_929(s929, c929, in929_1, in929_2);
    wire[0:0] s930, in930_1, in930_2;
    wire c930;
    assign in930_1 = {c905};
    assign in930_2 = {c913};
    Half_Adder KS_930(s930, c930, in930_1, in930_2);
    wire[3:0] s931, in931_1, in931_2;
    wire c931;
    assign in931_1 = {s914[0],s917[1],c469,c464};
    assign in931_2 = {s915[0],s918[1],s914[2],s466[2]};
    CLA_4 KS_931(s931, c931, in931_1, in931_2);
    wire[0:0] s932, in932_1, in932_2;
    wire c932;
    assign in932_1 = {s917[0]};
    assign in932_2 = {s918[0]};
    Full_Adder KS_932(s932, c932, in932_1, in932_2, s916[0]);
    wire[3:0] s933, in933_1, in933_2;
    wire c933;
    assign in933_1 = {s84[0],s478[0],s478[1],s470[2]};
    assign in933_2 = {s85[0],s479[0],s479[1],s471[2]};
    CLA_4 KS_933(s933, c933, in933_1, in933_2);
    wire[3:0] s934, in934_1, in934_2;
    wire c934;
    assign in934_1 = {s86[0],s480[0],s480[1],s472[2]};
    assign in934_2 = {s87[0],s481[0],s481[1],s473[2]};
    CLA_4 KS_934(s934, c934, in934_1, in934_2);
    wire[3:0] s935, in935_1, in935_2;
    wire c935;
    assign in935_1 = {s439[3],s482[0],s482[1],s474[2]};
    assign in935_2 = {s440[3],s483[0],s483[1],s475[2]};
    CLA_4 KS_935(s935, c935, in935_1, in935_2);
    wire[3:0] s936, in936_1, in936_2;
    wire c936;
    assign in936_1 = {s441[3],s484[0],s484[1],s476[2]};
    assign in936_2 = {s442[3],s485[0],s485[1],s477[2]};
    CLA_4 KS_936(s936, c936, in936_1, in936_2);
    wire[3:0] s937, in937_1, in937_2;
    wire c937;
    assign in937_1 = {s443[3],s486[0],c486,s478[2]};
    assign in937_2 = {s444[3],s487[0],s487[1],s479[2]};
    CLA_4 KS_937(s937, c937, in937_1, in937_2);
    wire[3:0] s938, in938_1, in938_2;
    wire c938;
    assign in938_1 = {s445[3],s488[0],c488,s480[2]};
    assign in938_2 = {s446[3],s489[0],s489[1],s481[2]};
    CLA_4 KS_938(s938, c938, in938_1, in938_2);
    wire[3:0] s939, in939_1, in939_2;
    wire c939;
    assign in939_1 = {s447[3],s490[0],c490,s482[2]};
    assign in939_2 = {s448[3],s491[0],s491[1],s483[2]};
    CLA_4 KS_939(s939, c939, in939_1, in939_2);
    wire[3:0] s940, in940_1, in940_2;
    wire c940;
    assign in940_1 = {s449[3],s492[0],c492,s484[2]};
    assign in940_2 = {s450[3],s493[0],s493[1],s485[2]};
    CLA_4 KS_940(s940, c940, in940_1, in940_2);
    wire[3:0] s941, in941_1, in941_2;
    wire c941;
    assign in941_1 = {s451[3],s494[0],c494,c487};
    assign in941_2 = {s452[3],s495[0],s495[1],s489[2]};
    CLA_4 KS_941(s941, c941, in941_1, in941_2);
    wire[3:0] s942, in942_1, in942_2;
    wire c942;
    assign in942_1 = {s453[3],s496[0],c496,c491};
    assign in942_2 = {s454[3],s497[0],s497[1],s493[2]};
    CLA_4 KS_942(s942, c942, in942_1, in942_2);
    wire[0:0] s943, in943_1, in943_2;
    wire c943;
    assign in943_1 = {c458};
    assign in943_2 = {s462[3]};
    Half_Adder KS_943(s943, c943, in943_1, in943_2);
    wire[1:0] s944, in944_1, in944_2;
    wire c944;
    assign in944_1 = {c466,s498[0]};
    assign in944_2 = {c914,s499[0]};
    CLA_2 KS_944(s944, c944, in944_1, in944_2);
    wire[0:0] s945, in945_1, in945_2;
    wire c945;
    assign in945_1 = {c915};
    assign in945_2 = {c916};
    Half_Adder KS_945(s945, c945, in945_1, in945_2);
    wire[2:0] s946, in946_1, in946_2;
    wire c946;
    assign in946_1 = {c917,s500[0],c498};
    assign in946_2 = {c918,s933[1],s499[1]};
    CLA_3 KS_946(s946, c946, in946_1, in946_2);
    wire[0:0] s947, in947_1, in947_2;
    wire c947;
    assign in947_1 = {c919};
    assign in947_2 = {c920};
    Half_Adder KS_947(s947, c947, in947_1, in947_2);
    wire[1:0] s948, in948_1, in948_2;
    wire c948;
    assign in948_1 = {c921,s934[1]};
    assign in948_2 = {c922,s935[1]};
    CLA_2 KS_948(s948, c948, in948_1, in948_2);
    wire[0:0] s949, in949_1, in949_2;
    wire c949;
    assign in949_1 = {c923};
    assign in949_2 = {c931};
    Half_Adder KS_949(s949, c949, in949_1, in949_2);
    wire[3:0] s950, in950_1, in950_2;
    wire c950;
    assign in950_1 = {s933[0],s936[1],c500,c495};
    assign in950_2 = {s934[0],s937[1],s933[2],s497[2]};
    CLA_4 KS_950(s950, c950, in950_1, in950_2);
    wire[0:0] s951, in951_1, in951_2;
    wire c951;
    assign in951_1 = {s936[0]};
    assign in951_2 = {s937[0]};
    Full_Adder KS_951(s951, c951, in951_1, in951_2, s935[0]);
    wire[3:0] s952, in952_1, in952_2;
    wire c952;
    assign in952_1 = {s125[0],s508[0],s509[1],s501[2]};
    assign in952_2 = {s126[0],s509[0],s510[1],s502[2]};
    CLA_4 KS_952(s952, c952, in952_1, in952_2);
    wire[3:0] s953, in953_1, in953_2;
    wire c953;
    assign in953_1 = {s127[0],s510[0],s511[1],s503[2]};
    assign in953_2 = {s128[0],s511[0],s512[1],s504[2]};
    CLA_4 KS_953(s953, c953, in953_1, in953_2);
    wire[3:0] s954, in954_1, in954_2;
    wire c954;
    assign in954_1 = {s470[3],s512[0],s513[1],s505[2]};
    assign in954_2 = {s471[3],s513[0],s514[1],s506[2]};
    CLA_4 KS_954(s954, c954, in954_1, in954_2);
    wire[3:0] s955, in955_1, in955_2;
    wire c955;
    assign in955_1 = {s472[3],s514[0],s515[1],s507[2]};
    assign in955_2 = {s473[3],s515[0],s516[1],s508[2]};
    CLA_4 KS_955(s955, c955, in955_1, in955_2);
    wire[3:0] s956, in956_1, in956_2;
    wire c956;
    assign in956_1 = {s474[3],s516[0],c517,s509[2]};
    assign in956_2 = {s475[3],s517[0],s518[1],s510[2]};
    CLA_4 KS_956(s956, c956, in956_1, in956_2);
    wire[3:0] s957, in957_1, in957_2;
    wire c957;
    assign in957_1 = {s476[3],s518[0],c519,s511[2]};
    assign in957_2 = {s477[3],s519[0],s520[1],s512[2]};
    CLA_4 KS_957(s957, c957, in957_1, in957_2);
    wire[3:0] s958, in958_1, in958_2;
    wire c958;
    assign in958_1 = {s478[3],s520[0],c521,s513[2]};
    assign in958_2 = {s479[3],s521[0],s522[1],s514[2]};
    CLA_4 KS_958(s958, c958, in958_1, in958_2);
    wire[3:0] s959, in959_1, in959_2;
    wire c959;
    assign in959_1 = {s480[3],s522[0],c523,s515[2]};
    assign in959_2 = {s481[3],s523[0],s524[1],s516[2]};
    CLA_4 KS_959(s959, c959, in959_1, in959_2);
    wire[3:0] s960, in960_1, in960_2;
    wire c960;
    assign in960_1 = {s482[3],s524[0],c525,c518};
    assign in960_2 = {s483[3],s525[0],s526[1],s520[2]};
    CLA_4 KS_960(s960, c960, in960_1, in960_2);
    wire[1:0] s961, in961_1, in961_2;
    wire c961;
    assign in961_1 = {s484[3],s526[0]};
    assign in961_2 = {s485[3],s527[0]};
    CLA_2 KS_961(s961, c961, in961_1, in961_2);
    wire[0:0] s962, in962_1, in962_2;
    wire c962;
    assign in962_1 = {c489};
    assign in962_2 = {s493[3]};
    Half_Adder KS_962(s962, c962, in962_1, in962_2);
    wire[3:0] s963, in963_1, in963_2;
    wire c963;
    assign in963_1 = {c497,s528[0],c527,c522};
    assign in963_2 = {c933,s529[0],s528[1],s524[2]};
    CLA_4 KS_963(s963, c963, in963_1, in963_2);
    wire[0:0] s964, in964_1, in964_2;
    wire c964;
    assign in964_1 = {c934};
    assign in964_2 = {c935};
    Half_Adder KS_964(s964, c964, in964_1, in964_2);
    wire[1:0] s965, in965_1, in965_2;
    wire c965;
    assign in965_1 = {c936,s530[0]};
    assign in965_2 = {c937,s952[1]};
    CLA_2 KS_965(s965, c965, in965_1, in965_2);
    wire[0:0] s966, in966_1, in966_2;
    wire c966;
    assign in966_1 = {c938};
    assign in966_2 = {c939};
    Half_Adder KS_966(s966, c966, in966_1, in966_2);
    wire[2:0] s967, in967_1, in967_2;
    wire c967;
    assign in967_1 = {c940,s953[1],c529};
    assign in967_2 = {c941,s954[1],s530[1]};
    CLA_3 KS_967(s967, c967, in967_1, in967_2);
    wire[0:0] s968, in968_1, in968_2;
    wire c968;
    assign in968_1 = {c942};
    assign in968_2 = {c950};
    Half_Adder KS_968(s968, c968, in968_1, in968_2);
    wire[1:0] s969, in969_1, in969_2;
    wire c969;
    assign in969_1 = {s952[0],s955[1]};
    assign in969_2 = {s953[0],s956[1]};
    CLA_2 KS_969(s969, c969, in969_1, in969_2);
    wire[0:0] s970, in970_1, in970_2;
    wire c970;
    assign in970_1 = {s955[0]};
    assign in970_2 = {s956[0]};
    Full_Adder KS_970(s970, c970, in970_1, in970_2, s954[0]);
    wire[3:0] s971, in971_1, in971_2;
    wire c971;
    assign in971_1 = {s170[0],s538[0],s538[1],s531[2]};
    assign in971_2 = {s171[0],s539[0],s539[1],s532[2]};
    CLA_4 KS_971(s971, c971, in971_1, in971_2);
    wire[3:0] s972, in972_1, in972_2;
    wire c972;
    assign in972_1 = {s172[0],s540[0],s540[1],s533[2]};
    assign in972_2 = {s173[0],s541[0],s541[1],s534[2]};
    CLA_4 KS_972(s972, c972, in972_1, in972_2);
    wire[3:0] s973, in973_1, in973_2;
    wire c973;
    assign in973_1 = {s501[3],s542[0],s542[1],s535[2]};
    assign in973_2 = {s502[3],s543[0],s543[1],s536[2]};
    CLA_4 KS_973(s973, c973, in973_1, in973_2);
    wire[3:0] s974, in974_1, in974_2;
    wire c974;
    assign in974_1 = {s503[3],s544[0],s544[1],s537[2]};
    assign in974_2 = {s504[3],s545[0],s545[1],s538[2]};
    CLA_4 KS_974(s974, c974, in974_1, in974_2);
    wire[3:0] s975, in975_1, in975_2;
    wire c975;
    assign in975_1 = {s505[3],s546[0],c546,s539[2]};
    assign in975_2 = {s506[3],s547[0],s547[1],s540[2]};
    CLA_4 KS_975(s975, c975, in975_1, in975_2);
    wire[3:0] s976, in976_1, in976_2;
    wire c976;
    assign in976_1 = {s507[3],s548[0],c548,s541[2]};
    assign in976_2 = {s508[3],s549[0],s549[1],s542[2]};
    CLA_4 KS_976(s976, c976, in976_1, in976_2);
    wire[3:0] s977, in977_1, in977_2;
    wire c977;
    assign in977_1 = {s509[3],s550[0],c550,s543[2]};
    assign in977_2 = {s510[3],s551[0],s551[1],s544[2]};
    CLA_4 KS_977(s977, c977, in977_1, in977_2);
    wire[3:0] s978, in978_1, in978_2;
    wire c978;
    assign in978_1 = {s511[3],s552[0],c552,s545[2]};
    assign in978_2 = {s512[3],s553[0],s553[1],s547[2]};
    CLA_4 KS_978(s978, c978, in978_1, in978_2);
    wire[3:0] s979, in979_1, in979_2;
    wire c979;
    assign in979_1 = {s513[3],s554[0],c554,c549};
    assign in979_2 = {s514[3],s555[0],s555[1],s551[2]};
    CLA_4 KS_979(s979, c979, in979_1, in979_2);
    wire[2:0] s980, in980_1, in980_2;
    wire c980;
    assign in980_1 = {s515[3],s556[0],c556};
    assign in980_2 = {s516[3],s557[0],s557[1]};
    CLA_3 KS_980(s980, c980, in980_1, in980_2);
    wire[0:0] s981, in981_1, in981_2;
    wire c981;
    assign in981_1 = {c520};
    assign in981_2 = {s524[3]};
    Half_Adder KS_981(s981, c981, in981_1, in981_2);
    wire[1:0] s982, in982_1, in982_2;
    wire c982;
    assign in982_1 = {c528,s558[0]};
    assign in982_2 = {c952,s559[0]};
    CLA_2 KS_982(s982, c982, in982_1, in982_2);
    wire[0:0] s983, in983_1, in983_2;
    wire c983;
    assign in983_1 = {c953};
    assign in983_2 = {c954};
    Half_Adder KS_983(s983, c983, in983_1, in983_2);
    wire[3:0] s984, in984_1, in984_2;
    wire c984;
    assign in984_1 = {c955,s560[0],c558,c553};
    assign in984_2 = {c956,s971[1],s559[1],s555[2]};
    CLA_4 KS_984(s984, c984, in984_1, in984_2);
    wire[0:0] s985, in985_1, in985_2;
    wire c985;
    assign in985_1 = {c957};
    assign in985_2 = {c958};
    Half_Adder KS_985(s985, c985, in985_1, in985_2);
    wire[1:0] s986, in986_1, in986_2;
    wire c986;
    assign in986_1 = {c959,s972[1]};
    assign in986_2 = {c960,s973[1]};
    CLA_2 KS_986(s986, c986, in986_1, in986_2);
    wire[0:0] s987, in987_1, in987_2;
    wire c987;
    assign in987_1 = {c963};
    assign in987_2 = {s971[0]};
    Half_Adder KS_987(s987, c987, in987_1, in987_2);
    wire[2:0] s988, in988_1, in988_2;
    wire c988;
    assign in988_1 = {s973[0],s974[1],c560};
    assign in988_2 = {s974[0],s975[1],s971[2]};
    CLA_3_c KS_988(s988, c988, in988_1, in988_2, s972[0]);
    wire[3:0] s989, in989_1, in989_2;
    wire c989;
    assign in989_1 = {s211[0],s568[0],s568[1],s561[2]};
    assign in989_2 = {s212[0],s569[0],s569[1],s562[2]};
    CLA_4 KS_989(s989, c989, in989_1, in989_2);
    wire[3:0] s990, in990_1, in990_2;
    wire c990;
    assign in990_1 = {s213[0],s570[0],s570[1],s563[2]};
    assign in990_2 = {s214[0],s571[0],s571[1],s564[2]};
    CLA_4 KS_990(s990, c990, in990_1, in990_2);
    wire[3:0] s991, in991_1, in991_2;
    wire c991;
    assign in991_1 = {s531[3],s572[0],s572[1],s565[2]};
    assign in991_2 = {s532[3],s573[0],s573[1],s566[2]};
    CLA_4 KS_991(s991, c991, in991_1, in991_2);
    wire[3:0] s992, in992_1, in992_2;
    wire c992;
    assign in992_1 = {s533[3],s574[0],s574[1],s567[2]};
    assign in992_2 = {s534[3],s575[0],s575[1],s568[2]};
    CLA_4 KS_992(s992, c992, in992_1, in992_2);
    wire[3:0] s993, in993_1, in993_2;
    wire c993;
    assign in993_1 = {s535[3],s576[0],c576,s569[2]};
    assign in993_2 = {s536[3],s577[0],s577[1],s570[2]};
    CLA_4 KS_993(s993, c993, in993_1, in993_2);
    wire[3:0] s994, in994_1, in994_2;
    wire c994;
    assign in994_1 = {s537[3],s578[0],c578,s571[2]};
    assign in994_2 = {s538[3],s579[0],s579[1],s572[2]};
    CLA_4 KS_994(s994, c994, in994_1, in994_2);
    wire[3:0] s995, in995_1, in995_2;
    wire c995;
    assign in995_1 = {s539[3],s580[0],c580,s573[2]};
    assign in995_2 = {s540[3],s581[0],s581[1],s574[2]};
    CLA_4 KS_995(s995, c995, in995_1, in995_2);
    wire[3:0] s996, in996_1, in996_2;
    wire c996;
    assign in996_1 = {s541[3],s582[0],c582,s575[2]};
    assign in996_2 = {s542[3],s583[0],s583[1],s577[2]};
    CLA_4 KS_996(s996, c996, in996_1, in996_2);
    wire[3:0] s997, in997_1, in997_2;
    wire c997;
    assign in997_1 = {s543[3],s584[0],c584,c579};
    assign in997_2 = {s544[3],s585[0],s585[1],s581[2]};
    CLA_4 KS_997(s997, c997, in997_1, in997_2);
    wire[2:0] s998, in998_1, in998_2;
    wire c998;
    assign in998_1 = {s545[3],s586[0],c586};
    assign in998_2 = {s547[3],s587[0],s587[1]};
    CLA_3 KS_998(s998, c998, in998_1, in998_2);
    wire[0:0] s999, in999_1, in999_2;
    wire c999;
    assign in999_1 = {c551};
    assign in999_2 = {s555[3]};
    Half_Adder KS_999(s999, c999, in999_1, in999_2);
    wire[1:0] s1000, in1000_1, in1000_2;
    wire c1000;
    assign in1000_1 = {c559,s588[0]};
    assign in1000_2 = {c971,s589[0]};
    CLA_2 KS_1000(s1000, c1000, in1000_1, in1000_2);
    wire[0:0] s1001, in1001_1, in1001_2;
    wire c1001;
    assign in1001_1 = {c972};
    assign in1001_2 = {c973};
    Half_Adder KS_1001(s1001, c1001, in1001_1, in1001_2);
    wire[3:0] s1002, in1002_1, in1002_2;
    wire c1002;
    assign in1002_1 = {c974,s590[0],c588,c583};
    assign in1002_2 = {c975,s989[1],s589[1],s585[2]};
    CLA_4 KS_1002(s1002, c1002, in1002_1, in1002_2);
    wire[0:0] s1003, in1003_1, in1003_2;
    wire c1003;
    assign in1003_1 = {c976};
    assign in1003_2 = {c977};
    Half_Adder KS_1003(s1003, c1003, in1003_1, in1003_2);
    wire[1:0] s1004, in1004_1, in1004_2;
    wire c1004;
    assign in1004_1 = {c978,s990[1]};
    assign in1004_2 = {c979,s991[1]};
    CLA_2 KS_1004(s1004, c1004, in1004_1, in1004_2);
    wire[0:0] s1005, in1005_1, in1005_2;
    wire c1005;
    assign in1005_1 = {c984};
    assign in1005_2 = {s989[0]};
    Half_Adder KS_1005(s1005, c1005, in1005_1, in1005_2);
    wire[2:0] s1006, in1006_1, in1006_2;
    wire c1006;
    assign in1006_1 = {s991[0],s992[1],c590};
    assign in1006_2 = {s992[0],s993[1],s989[2]};
    CLA_3_c KS_1006(s1006, c1006, in1006_1, in1006_2, s990[0]);
    wire[3:0] s1007, in1007_1, in1007_2;
    wire c1007;
    assign in1007_1 = {s245[0],s599[0],s600[1],s592[2]};
    assign in1007_2 = {s246[0],s600[0],s601[1],s593[2]};
    CLA_4 KS_1007(s1007, c1007, in1007_1, in1007_2);
    wire[3:0] s1008, in1008_1, in1008_2;
    wire c1008;
    assign in1008_1 = {s247[0],s601[0],s602[1],s594[2]};
    assign in1008_2 = {s248[0],s602[0],s603[1],s595[2]};
    CLA_4 KS_1008(s1008, c1008, in1008_1, in1008_2);
    wire[3:0] s1009, in1009_1, in1009_2;
    wire c1009;
    assign in1009_1 = {s561[3],s603[0],s604[1],s596[2]};
    assign in1009_2 = {s562[3],s604[0],s605[1],s597[2]};
    CLA_4 KS_1009(s1009, c1009, in1009_1, in1009_2);
    wire[3:0] s1010, in1010_1, in1010_2;
    wire c1010;
    assign in1010_1 = {s563[3],s605[0],c606,s598[2]};
    assign in1010_2 = {s564[3],s606[0],s607[1],s599[2]};
    CLA_4 KS_1010(s1010, c1010, in1010_1, in1010_2);
    wire[3:0] s1011, in1011_1, in1011_2;
    wire c1011;
    assign in1011_1 = {s565[3],s607[0],c608,s600[2]};
    assign in1011_2 = {s566[3],s608[0],s609[1],s601[2]};
    CLA_4 KS_1011(s1011, c1011, in1011_1, in1011_2);
    wire[3:0] s1012, in1012_1, in1012_2;
    wire c1012;
    assign in1012_1 = {s567[3],s609[0],c610,s602[2]};
    assign in1012_2 = {s568[3],s610[0],s611[1],s603[2]};
    CLA_4 KS_1012(s1012, c1012, in1012_1, in1012_2);
    wire[3:0] s1013, in1013_1, in1013_2;
    wire c1013;
    assign in1013_1 = {s569[3],s611[0],c612,s604[2]};
    assign in1013_2 = {s570[3],s612[0],s613[1],s605[2]};
    CLA_4 KS_1013(s1013, c1013, in1013_1, in1013_2);
    wire[3:0] s1014, in1014_1, in1014_2;
    wire c1014;
    assign in1014_1 = {s571[3],s613[0],c614,c607};
    assign in1014_2 = {s572[3],s614[0],s615[1],s609[2]};
    CLA_4 KS_1014(s1014, c1014, in1014_1, in1014_2);
    wire[3:0] s1015, in1015_1, in1015_2;
    wire c1015;
    assign in1015_1 = {s573[3],s615[0],c616,c611};
    assign in1015_2 = {s574[3],s616[0],s617[1],s613[2]};
    CLA_4 KS_1015(s1015, c1015, in1015_1, in1015_2);
    wire[1:0] s1016, in1016_1, in1016_2;
    wire c1016;
    assign in1016_1 = {s575[3],s617[0]};
    assign in1016_2 = {s577[3],s618[0]};
    CLA_2 KS_1016(s1016, c1016, in1016_1, in1016_2);
    wire[0:0] s1017, in1017_1, in1017_2;
    wire c1017;
    assign in1017_1 = {c581};
    assign in1017_2 = {s585[3]};
    Half_Adder KS_1017(s1017, c1017, in1017_1, in1017_2);
    wire[2:0] s1018, in1018_1, in1018_2;
    wire c1018;
    assign in1018_1 = {c589,s619[0],c618};
    assign in1018_2 = {c989,s620[0],s619[1]};
    CLA_3 KS_1018(s1018, c1018, in1018_1, in1018_2);
    wire[0:0] s1019, in1019_1, in1019_2;
    wire c1019;
    assign in1019_1 = {c990};
    assign in1019_2 = {c991};
    Half_Adder KS_1019(s1019, c1019, in1019_1, in1019_2);
    wire[1:0] s1020, in1020_1, in1020_2;
    wire c1020;
    assign in1020_1 = {c992,s621[0]};
    assign in1020_2 = {c993,s1007[1]};
    CLA_2 KS_1020(s1020, c1020, in1020_1, in1020_2);
    wire[0:0] s1021, in1021_1, in1021_2;
    wire c1021;
    assign in1021_1 = {c994};
    assign in1021_2 = {c995};
    Half_Adder KS_1021(s1021, c1021, in1021_1, in1021_2);
    wire[3:0] s1022, in1022_1, in1022_2;
    wire c1022;
    assign in1022_1 = {c996,s1008[1],c620,c615};
    assign in1022_2 = {c997,s1009[1],s621[1],s617[2]};
    CLA_4 KS_1022(s1022, c1022, in1022_1, in1022_2);
    wire[0:0] s1023, in1023_1, in1023_2;
    wire c1023;
    assign in1023_1 = {c1002};
    assign in1023_2 = {s1007[0]};
    Half_Adder KS_1023(s1023, c1023, in1023_1, in1023_2);
    wire[1:0] s1024, in1024_1, in1024_2;
    wire c1024;
    assign in1024_1 = {s1009[0],s1010[1]};
    assign in1024_2 = {s1010[0],s1011[1]};
    CLA_2_c KS_1024(s1024, c1024, in1024_1, in1024_2, s1008[0]);
    wire[3:0] s1025, in1025_1, in1025_2;
    wire c1025;
    assign in1025_1 = {s271[0],s630[0],s631[1],s622[2]};
    assign in1025_2 = {s272[0],s631[0],s632[1],s623[2]};
    CLA_4 KS_1025(s1025, c1025, in1025_1, in1025_2);
    wire[3:0] s1026, in1026_1, in1026_2;
    wire c1026;
    assign in1026_1 = {s273[0],s632[0],s633[1],s624[2]};
    assign in1026_2 = {s274[0],s633[0],s634[1],s625[2]};
    CLA_4 KS_1026(s1026, c1026, in1026_1, in1026_2);
    wire[3:0] s1027, in1027_1, in1027_2;
    wire c1027;
    assign in1027_1 = {s591[3],s634[0],s635[1],s626[2]};
    assign in1027_2 = {s592[3],s635[0],s636[1],s627[2]};
    CLA_4 KS_1027(s1027, c1027, in1027_1, in1027_2);
    wire[3:0] s1028, in1028_1, in1028_2;
    wire c1028;
    assign in1028_1 = {s593[3],s636[0],c637,s628[2]};
    assign in1028_2 = {s594[3],s637[0],s638[1],s629[2]};
    CLA_4 KS_1028(s1028, c1028, in1028_1, in1028_2);
    wire[3:0] s1029, in1029_1, in1029_2;
    wire c1029;
    assign in1029_1 = {s595[3],s638[0],c639,s630[2]};
    assign in1029_2 = {s596[3],s639[0],s640[1],s631[2]};
    CLA_4 KS_1029(s1029, c1029, in1029_1, in1029_2);
    wire[3:0] s1030, in1030_1, in1030_2;
    wire c1030;
    assign in1030_1 = {s597[3],s640[0],c641,s632[2]};
    assign in1030_2 = {s598[3],s641[0],s642[1],s633[2]};
    CLA_4 KS_1030(s1030, c1030, in1030_1, in1030_2);
    wire[3:0] s1031, in1031_1, in1031_2;
    wire c1031;
    assign in1031_1 = {s599[3],s642[0],c643,s634[2]};
    assign in1031_2 = {s600[3],s643[0],s644[1],s635[2]};
    CLA_4 KS_1031(s1031, c1031, in1031_1, in1031_2);
    wire[3:0] s1032, in1032_1, in1032_2;
    wire c1032;
    assign in1032_1 = {s601[3],s644[0],c645,s636[2]};
    assign in1032_2 = {s602[3],s645[0],s646[1],s638[2]};
    CLA_4 KS_1032(s1032, c1032, in1032_1, in1032_2);
    wire[3:0] s1033, in1033_1, in1033_2;
    wire c1033;
    assign in1033_1 = {s603[3],s646[0],c647,c640};
    assign in1033_2 = {s604[3],s647[0],s648[1],s642[2]};
    CLA_4 KS_1033(s1033, c1033, in1033_1, in1033_2);
    wire[1:0] s1034, in1034_1, in1034_2;
    wire c1034;
    assign in1034_1 = {s605[3],s648[0]};
    assign in1034_2 = {s609[3],s649[0]};
    CLA_2 KS_1034(s1034, c1034, in1034_1, in1034_2);
    wire[0:0] s1035, in1035_1, in1035_2;
    wire c1035;
    assign in1035_1 = {c613};
    assign in1035_2 = {s617[3]};
    Half_Adder KS_1035(s1035, c1035, in1035_1, in1035_2);
    wire[3:0] s1036, in1036_1, in1036_2;
    wire c1036;
    assign in1036_1 = {c621,s650[0],c649,c644};
    assign in1036_2 = {c1007,s651[0],s650[1],s646[2]};
    CLA_4 KS_1036(s1036, c1036, in1036_1, in1036_2);
    wire[0:0] s1037, in1037_1, in1037_2;
    wire c1037;
    assign in1037_1 = {c1008};
    assign in1037_2 = {c1009};
    Half_Adder KS_1037(s1037, c1037, in1037_1, in1037_2);
    wire[1:0] s1038, in1038_1, in1038_2;
    wire c1038;
    assign in1038_1 = {c1010,s652[0]};
    assign in1038_2 = {c1011,s1025[1]};
    CLA_2 KS_1038(s1038, c1038, in1038_1, in1038_2);
    wire[0:0] s1039, in1039_1, in1039_2;
    wire c1039;
    assign in1039_1 = {c1012};
    assign in1039_2 = {c1013};
    Half_Adder KS_1039(s1039, c1039, in1039_1, in1039_2);
    wire[2:0] s1040, in1040_1, in1040_2;
    wire c1040;
    assign in1040_1 = {c1014,s1026[1],c651};
    assign in1040_2 = {c1015,s1027[1],s652[1]};
    CLA_3 KS_1040(s1040, c1040, in1040_1, in1040_2);
    wire[0:0] s1041, in1041_1, in1041_2;
    wire c1041;
    assign in1041_1 = {c1022};
    assign in1041_2 = {s1025[0]};
    Half_Adder KS_1041(s1041, c1041, in1041_1, in1041_2);
    wire[1:0] s1042, in1042_1, in1042_2;
    wire c1042;
    assign in1042_1 = {s1027[0],s1028[1]};
    assign in1042_2 = {s1028[0],s1029[1]};
    CLA_2_c KS_1042(s1042, c1042, in1042_1, in1042_2, s1026[0]);
    wire[3:0] s1043, in1043_1, in1043_2;
    wire c1043;
    assign in1043_1 = {s288[0],s660[0],s660[1],s291[3]};
    assign in1043_2 = {s289[0],s661[0],s661[1],s653[2]};
    CLA_4 KS_1043(s1043, c1043, in1043_1, in1043_2);
    wire[3:0] s1044, in1044_1, in1044_2;
    wire c1044;
    assign in1044_1 = {s290[0],s662[0],s662[1],s654[2]};
    assign in1044_2 = {s291[0],s663[0],s663[1],s655[2]};
    CLA_4 KS_1044(s1044, c1044, in1044_1, in1044_2);
    wire[3:0] s1045, in1045_1, in1045_2;
    wire c1045;
    assign in1045_1 = {s622[3],s664[0],s664[1],s656[2]};
    assign in1045_2 = {s623[3],s665[0],s665[1],s657[2]};
    CLA_4 KS_1045(s1045, c1045, in1045_1, in1045_2);
    wire[3:0] s1046, in1046_1, in1046_2;
    wire c1046;
    assign in1046_1 = {s624[3],s666[0],s666[1],s658[2]};
    assign in1046_2 = {s625[3],s667[0],s667[1],s659[2]};
    CLA_4 KS_1046(s1046, c1046, in1046_1, in1046_2);
    wire[3:0] s1047, in1047_1, in1047_2;
    wire c1047;
    assign in1047_1 = {s626[3],s668[0],c668,s660[2]};
    assign in1047_2 = {s627[3],s669[0],s669[1],s661[2]};
    CLA_4 KS_1047(s1047, c1047, in1047_1, in1047_2);
    wire[3:0] s1048, in1048_1, in1048_2;
    wire c1048;
    assign in1048_1 = {s628[3],s670[0],c670,s662[2]};
    assign in1048_2 = {s629[3],s671[0],s671[1],s663[2]};
    CLA_4 KS_1048(s1048, c1048, in1048_1, in1048_2);
    wire[3:0] s1049, in1049_1, in1049_2;
    wire c1049;
    assign in1049_1 = {s630[3],s672[0],c672,s664[2]};
    assign in1049_2 = {s631[3],s673[0],s673[1],s665[2]};
    CLA_4 KS_1049(s1049, c1049, in1049_1, in1049_2);
    wire[3:0] s1050, in1050_1, in1050_2;
    wire c1050;
    assign in1050_1 = {s632[3],s674[0],c674,s666[2]};
    assign in1050_2 = {s633[3],s675[0],s675[1],s667[2]};
    CLA_4 KS_1050(s1050, c1050, in1050_1, in1050_2);
    wire[3:0] s1051, in1051_1, in1051_2;
    wire c1051;
    assign in1051_1 = {s634[3],s676[0],c676,c669};
    assign in1051_2 = {s635[3],s677[0],s677[1],s671[2]};
    CLA_4 KS_1051(s1051, c1051, in1051_1, in1051_2);
    wire[3:0] s1052, in1052_1, in1052_2;
    wire c1052;
    assign in1052_1 = {s636[3],s678[0],c678,c673};
    assign in1052_2 = {s638[3],s679[0],s679[1],s675[2]};
    CLA_4 KS_1052(s1052, c1052, in1052_1, in1052_2);
    wire[0:0] s1053, in1053_1, in1053_2;
    wire c1053;
    assign in1053_1 = {c642};
    assign in1053_2 = {s646[3]};
    Half_Adder KS_1053(s1053, c1053, in1053_1, in1053_2);
    wire[1:0] s1054, in1054_1, in1054_2;
    wire c1054;
    assign in1054_1 = {c650,s680[0]};
    assign in1054_2 = {c1025,s681[0]};
    CLA_2 KS_1054(s1054, c1054, in1054_1, in1054_2);
    wire[0:0] s1055, in1055_1, in1055_2;
    wire c1055;
    assign in1055_1 = {c1026};
    assign in1055_2 = {c1027};
    Half_Adder KS_1055(s1055, c1055, in1055_1, in1055_2);
    wire[2:0] s1056, in1056_1, in1056_2;
    wire c1056;
    assign in1056_1 = {c1028,s682[0],c680};
    assign in1056_2 = {c1029,s1043[1],s681[1]};
    CLA_3 KS_1056(s1056, c1056, in1056_1, in1056_2);
    wire[0:0] s1057, in1057_1, in1057_2;
    wire c1057;
    assign in1057_1 = {c1030};
    assign in1057_2 = {c1031};
    Half_Adder KS_1057(s1057, c1057, in1057_1, in1057_2);
    wire[1:0] s1058, in1058_1, in1058_2;
    wire c1058;
    assign in1058_1 = {c1032,s1044[1]};
    assign in1058_2 = {c1033,s1045[1]};
    CLA_2 KS_1058(s1058, c1058, in1058_1, in1058_2);
    wire[0:0] s1059, in1059_1, in1059_2;
    wire c1059;
    assign in1059_1 = {c1036};
    assign in1059_2 = {s1043[0]};
    Half_Adder KS_1059(s1059, c1059, in1059_1, in1059_2);
    wire[3:0] s1060, in1060_1, in1060_2;
    wire c1060;
    assign in1060_1 = {s1045[0],s1046[1],c682,c677};
    assign in1060_2 = {s1046[0],s1047[1],s1043[2],s679[2]};
    CLA_4_c KS_1060(s1060, c1060, in1060_1, in1060_2, s1044[0]);
    wire[3:0] s1061, in1061_1, in1061_2;
    wire c1061;
    assign in1061_1 = {s297[0],s690[0],s690[1],s683[2]};
    assign in1061_2 = {s298[0],s691[0],s691[1],s684[2]};
    CLA_4 KS_1061(s1061, c1061, in1061_1, in1061_2);
    wire[3:0] s1062, in1062_1, in1062_2;
    wire c1062;
    assign in1062_1 = {s299[0],s692[0],s692[1],s685[2]};
    assign in1062_2 = {s300[0],s693[0],s693[1],s686[2]};
    CLA_4 KS_1062(s1062, c1062, in1062_1, in1062_2);
    wire[3:0] s1063, in1063_1, in1063_2;
    wire c1063;
    assign in1063_1 = {s653[3],s694[0],s694[1],s687[2]};
    assign in1063_2 = {s654[3],s695[0],s695[1],s688[2]};
    CLA_4 KS_1063(s1063, c1063, in1063_1, in1063_2);
    wire[3:0] s1064, in1064_1, in1064_2;
    wire c1064;
    assign in1064_1 = {s655[3],s696[0],s696[1],s689[2]};
    assign in1064_2 = {s656[3],s697[0],s697[1],s690[2]};
    CLA_4 KS_1064(s1064, c1064, in1064_1, in1064_2);
    wire[3:0] s1065, in1065_1, in1065_2;
    wire c1065;
    assign in1065_1 = {s657[3],s698[0],c698,s691[2]};
    assign in1065_2 = {s658[3],s699[0],s699[1],s692[2]};
    CLA_4 KS_1065(s1065, c1065, in1065_1, in1065_2);
    wire[3:0] s1066, in1066_1, in1066_2;
    wire c1066;
    assign in1066_1 = {s659[3],s700[0],c700,s693[2]};
    assign in1066_2 = {s660[3],s701[0],s701[1],s694[2]};
    CLA_4 KS_1066(s1066, c1066, in1066_1, in1066_2);
    wire[3:0] s1067, in1067_1, in1067_2;
    wire c1067;
    assign in1067_1 = {s661[3],s702[0],c702,s695[2]};
    assign in1067_2 = {s662[3],s703[0],s703[1],s696[2]};
    CLA_4 KS_1067(s1067, c1067, in1067_1, in1067_2);
    wire[3:0] s1068, in1068_1, in1068_2;
    wire c1068;
    assign in1068_1 = {s663[3],s704[0],c704,s697[2]};
    assign in1068_2 = {s664[3],s705[0],s705[1],s699[2]};
    CLA_4 KS_1068(s1068, c1068, in1068_1, in1068_2);
    wire[3:0] s1069, in1069_1, in1069_2;
    wire c1069;
    assign in1069_1 = {s665[3],s706[0],c706,c701};
    assign in1069_2 = {s666[3],s707[0],s707[1],s703[2]};
    CLA_4 KS_1069(s1069, c1069, in1069_1, in1069_2);
    wire[2:0] s1070, in1070_1, in1070_2;
    wire c1070;
    assign in1070_1 = {s667[3],s708[0],c708};
    assign in1070_2 = {s671[3],s709[0],s709[1]};
    CLA_3 KS_1070(s1070, c1070, in1070_1, in1070_2);
    wire[0:0] s1071, in1071_1, in1071_2;
    wire c1071;
    assign in1071_1 = {c675};
    assign in1071_2 = {s679[3]};
    Half_Adder KS_1071(s1071, c1071, in1071_1, in1071_2);
    wire[1:0] s1072, in1072_1, in1072_2;
    wire c1072;
    assign in1072_1 = {c1043,s710[0]};
    assign in1072_2 = {c1044,s711[0]};
    CLA_2 KS_1072(s1072, c1072, in1072_1, in1072_2);
    wire[0:0] s1073, in1073_1, in1073_2;
    wire c1073;
    assign in1073_1 = {c1045};
    assign in1073_2 = {c1046};
    Half_Adder KS_1073(s1073, c1073, in1073_1, in1073_2);
    wire[3:0] s1074, in1074_1, in1074_2;
    wire c1074;
    assign in1074_1 = {c1047,s712[0],c710,c705};
    assign in1074_2 = {c1048,s1061[1],s711[1],s707[2]};
    CLA_4 KS_1074(s1074, c1074, in1074_1, in1074_2);
    wire[0:0] s1075, in1075_1, in1075_2;
    wire c1075;
    assign in1075_1 = {c1049};
    assign in1075_2 = {c1050};
    Half_Adder KS_1075(s1075, c1075, in1075_1, in1075_2);
    wire[1:0] s1076, in1076_1, in1076_2;
    wire c1076;
    assign in1076_1 = {c1051,s1062[1]};
    assign in1076_2 = {c1052,s1063[1]};
    CLA_2 KS_1076(s1076, c1076, in1076_1, in1076_2);
    wire[0:0] s1077, in1077_1, in1077_2;
    wire c1077;
    assign in1077_1 = {c1060};
    assign in1077_2 = {s1061[0]};
    Half_Adder KS_1077(s1077, c1077, in1077_1, in1077_2);
    wire[2:0] s1078, in1078_1, in1078_2;
    wire c1078;
    assign in1078_1 = {s1063[0],s1064[1],c712};
    assign in1078_2 = {s1064[0],s1065[1],s1061[2]};
    CLA_3_c KS_1078(s1078, c1078, in1078_1, in1078_2, s1062[0]);
    wire[3:0] s1079, in1079_1, in1079_2;
    wire c1079;
    assign in1079_1 = {pp63[27],s720[0],s720[1],pp62[31]};
    assign in1079_2 = {c292,s721[0],s721[1],pp63[30]};
    CLA_4 KS_1079(s1079, c1079, in1079_1, in1079_2);
    wire[3:0] s1080, in1080_1, in1080_2;
    wire c1080;
    assign in1080_1 = {c296,s722[0],s722[1],s713[2]};
    assign in1080_2 = {s301[0],s723[0],s723[1],s714[2]};
    CLA_4 KS_1080(s1080, c1080, in1080_1, in1080_2);
    wire[3:0] s1081, in1081_1, in1081_2;
    wire c1081;
    assign in1081_1 = {s683[3],s724[0],s724[1],s715[2]};
    assign in1081_2 = {s684[3],s725[0],s725[1],s716[2]};
    CLA_4 KS_1081(s1081, c1081, in1081_1, in1081_2);
    wire[3:0] s1082, in1082_1, in1082_2;
    wire c1082;
    assign in1082_1 = {s685[3],s726[0],c726,s717[2]};
    assign in1082_2 = {s686[3],s727[0],s727[1],s718[2]};
    CLA_4 KS_1082(s1082, c1082, in1082_1, in1082_2);
    wire[3:0] s1083, in1083_1, in1083_2;
    wire c1083;
    assign in1083_1 = {s687[3],s728[0],c728,s719[2]};
    assign in1083_2 = {s688[3],s729[0],s729[1],s720[2]};
    CLA_4 KS_1083(s1083, c1083, in1083_1, in1083_2);
    wire[3:0] s1084, in1084_1, in1084_2;
    wire c1084;
    assign in1084_1 = {s689[3],s730[0],c730,s721[2]};
    assign in1084_2 = {s690[3],s731[0],s731[1],s722[2]};
    CLA_4 KS_1084(s1084, c1084, in1084_1, in1084_2);
    wire[3:0] s1085, in1085_1, in1085_2;
    wire c1085;
    assign in1085_1 = {s691[3],s732[0],c732,s723[2]};
    assign in1085_2 = {s692[3],s733[0],s733[1],s724[2]};
    CLA_4 KS_1085(s1085, c1085, in1085_1, in1085_2);
    wire[3:0] s1086, in1086_1, in1086_2;
    wire c1086;
    assign in1086_1 = {s693[3],s734[0],c734,c725};
    assign in1086_2 = {s694[3],s735[0],s735[1],s727[2]};
    CLA_4 KS_1086(s1086, c1086, in1086_1, in1086_2);
    wire[3:0] s1087, in1087_1, in1087_2;
    wire c1087;
    assign in1087_1 = {s695[3],s736[0],c736,c729};
    assign in1087_2 = {s696[3],s737[0],s737[1],s731[2]};
    CLA_4 KS_1087(s1087, c1087, in1087_1, in1087_2);
    wire[3:0] s1088, in1088_1, in1088_2;
    wire c1088;
    assign in1088_1 = {s697[3],s738[0],c738,c733};
    assign in1088_2 = {s699[3],s739[0],s739[1],s735[2]};
    CLA_4 KS_1088(s1088, c1088, in1088_1, in1088_2);
    wire[0:0] s1089, in1089_1, in1089_2;
    wire c1089;
    assign in1089_1 = {c703};
    assign in1089_2 = {s707[3]};
    Half_Adder KS_1089(s1089, c1089, in1089_1, in1089_2);
    wire[1:0] s1090, in1090_1, in1090_2;
    wire c1090;
    assign in1090_1 = {c711,s740[0]};
    assign in1090_2 = {c1061,s741[0]};
    CLA_2 KS_1090(s1090, c1090, in1090_1, in1090_2);
    wire[0:0] s1091, in1091_1, in1091_2;
    wire c1091;
    assign in1091_1 = {c1062};
    assign in1091_2 = {c1063};
    Half_Adder KS_1091(s1091, c1091, in1091_1, in1091_2);
    wire[2:0] s1092, in1092_1, in1092_2;
    wire c1092;
    assign in1092_1 = {c1064,s742[0],c740};
    assign in1092_2 = {c1065,s1079[1],s741[1]};
    CLA_3 KS_1092(s1092, c1092, in1092_1, in1092_2);
    wire[0:0] s1093, in1093_1, in1093_2;
    wire c1093;
    assign in1093_1 = {c1066};
    assign in1093_2 = {c1067};
    Half_Adder KS_1093(s1093, c1093, in1093_1, in1093_2);
    wire[1:0] s1094, in1094_1, in1094_2;
    wire c1094;
    assign in1094_1 = {c1068,s1080[1]};
    assign in1094_2 = {c1069,s1081[1]};
    CLA_2 KS_1094(s1094, c1094, in1094_1, in1094_2);
    wire[0:0] s1095, in1095_1, in1095_2;
    wire c1095;
    assign in1095_1 = {c1074};
    assign in1095_2 = {s1079[0]};
    Half_Adder KS_1095(s1095, c1095, in1095_1, in1095_2);
    wire[3:0] s1096, in1096_1, in1096_2;
    wire c1096;
    assign in1096_1 = {s1081[0],s1082[1],c742,c737};
    assign in1096_2 = {s1082[0],s1083[1],s1079[2],s739[2]};
    CLA_4_c KS_1096(s1096, c1096, in1096_1, in1096_2, s1080[0]);
    wire[3:0] s1097, in1097_1, in1097_2;
    wire c1097;
    assign in1097_1 = {pp57[37],c727,pp63[33],pp56[41]};
    assign in1097_2 = {pp58[36],c735,s743[1],pp57[40]};
    CLA_4 KS_1097(s1097, c1097, in1097_1, in1097_2);
    wire[3:0] s1098, in1098_1, in1098_2;
    wire c1098;
    assign in1098_1 = {pp59[35],s743[0],s744[1],pp58[39]};
    assign in1098_2 = {pp60[34],s744[0],s745[1],pp59[38]};
    CLA_4 KS_1098(s1098, c1098, in1098_1, in1098_2);
    wire[3:0] s1099, in1099_1, in1099_2;
    wire c1099;
    assign in1099_1 = {pp61[33],s745[0],s746[1],pp60[37]};
    assign in1099_2 = {pp62[32],s746[0],s747[1],pp61[36]};
    CLA_4 KS_1099(s1099, c1099, in1099_1, in1099_2);
    wire[3:0] s1100, in1100_1, in1100_2;
    wire c1100;
    assign in1100_1 = {pp63[31],s747[0],s748[1],pp62[35]};
    assign in1100_2 = {s713[3],s748[0],s749[1],pp63[34]};
    CLA_4 KS_1100(s1100, c1100, in1100_1, in1100_2);
    wire[3:0] s1101, in1101_1, in1101_2;
    wire c1101;
    assign in1101_1 = {s714[3],s749[0],s750[1],s743[2]};
    assign in1101_2 = {s715[3],s750[0],s751[1],s744[2]};
    CLA_4 KS_1101(s1101, c1101, in1101_1, in1101_2);
    wire[3:0] s1102, in1102_1, in1102_2;
    wire c1102;
    assign in1102_1 = {s716[3],s751[0],c752,s745[2]};
    assign in1102_2 = {s717[3],s752[0],s753[1],s746[2]};
    CLA_4 KS_1102(s1102, c1102, in1102_1, in1102_2);
    wire[3:0] s1103, in1103_1, in1103_2;
    wire c1103;
    assign in1103_1 = {s718[3],s753[0],c754,s747[2]};
    assign in1103_2 = {s719[3],s754[0],s755[1],s748[2]};
    CLA_4 KS_1103(s1103, c1103, in1103_1, in1103_2);
    wire[3:0] s1104, in1104_1, in1104_2;
    wire c1104;
    assign in1104_1 = {s720[3],s755[0],c756,s749[2]};
    assign in1104_2 = {s721[3],s756[0],s757[1],s750[2]};
    CLA_4 KS_1104(s1104, c1104, in1104_1, in1104_2);
    wire[3:0] s1105, in1105_1, in1105_2;
    wire c1105;
    assign in1105_1 = {s722[3],s757[0],c758,c751};
    assign in1105_2 = {s723[3],s758[0],s759[1],s753[2]};
    CLA_4 KS_1105(s1105, c1105, in1105_1, in1105_2);
    wire[1:0] s1106, in1106_1, in1106_2;
    wire c1106;
    assign in1106_1 = {c724,s759[0]};
    assign in1106_2 = {s727[3],s760[0]};
    CLA_2 KS_1106(s1106, c1106, in1106_1, in1106_2);
    wire[0:0] s1107, in1107_1, in1107_2;
    wire c1107;
    assign in1107_1 = {c731};
    assign in1107_2 = {s735[3]};
    Half_Adder KS_1107(s1107, c1107, in1107_1, in1107_2);
    wire[3:0] s1108, in1108_1, in1108_2;
    wire c1108;
    assign in1108_1 = {c739,s761[0],c760,c755};
    assign in1108_2 = {c1079,s762[0],s761[1],s757[2]};
    CLA_4 KS_1108(s1108, c1108, in1108_1, in1108_2);
    wire[0:0] s1109, in1109_1, in1109_2;
    wire c1109;
    assign in1109_1 = {c1080};
    assign in1109_2 = {c1081};
    Half_Adder KS_1109(s1109, c1109, in1109_1, in1109_2);
    wire[1:0] s1110, in1110_1, in1110_2;
    wire c1110;
    assign in1110_1 = {c1082,s763[0]};
    assign in1110_2 = {c1083,s1097[1]};
    CLA_2 KS_1110(s1110, c1110, in1110_1, in1110_2);
    wire[0:0] s1111, in1111_1, in1111_2;
    wire c1111;
    assign in1111_1 = {c1084};
    assign in1111_2 = {c1085};
    Half_Adder KS_1111(s1111, c1111, in1111_1, in1111_2);
    wire[2:0] s1112, in1112_1, in1112_2;
    wire c1112;
    assign in1112_1 = {c1086,s1098[1],c762};
    assign in1112_2 = {c1087,s1099[1],s763[1]};
    CLA_3 KS_1112(s1112, c1112, in1112_1, in1112_2);
    wire[0:0] s1113, in1113_1, in1113_2;
    wire c1113;
    assign in1113_1 = {c1088};
    assign in1113_2 = {c1096};
    Half_Adder KS_1113(s1113, c1113, in1113_1, in1113_2);
    wire[1:0] s1114, in1114_1, in1114_2;
    wire c1114;
    assign in1114_1 = {s1097[0],s1100[1]};
    assign in1114_2 = {s1098[0],s1101[1]};
    CLA_2 KS_1114(s1114, c1114, in1114_1, in1114_2);
    wire[0:0] s1115, in1115_1, in1115_2;
    wire c1115;
    assign in1115_1 = {s1100[0]};
    assign in1115_2 = {s1101[0]};
    Full_Adder KS_1115(s1115, c1115, in1115_1, in1115_2, s1099[0]);
    wire[3:0] s1116, in1116_1, in1116_2;
    wire c1116;
    assign in1116_1 = {pp53[45],pp63[36],pp55[45],pp50[51]};
    assign in1116_2 = {pp54[44],c743,pp56[44],pp51[50]};
    CLA_4 KS_1116(s1116, c1116, in1116_1, in1116_2);
    wire[3:0] s1117, in1117_1, in1117_2;
    wire c1117;
    assign in1117_1 = {pp55[43],c744,pp57[43],pp52[49]};
    assign in1117_2 = {pp56[42],c745,pp58[42],pp53[48]};
    CLA_4 KS_1117(s1117, c1117, in1117_1, in1117_2);
    wire[3:0] s1118, in1118_1, in1118_2;
    wire c1118;
    assign in1118_1 = {pp57[41],c746,pp59[41],pp54[47]};
    assign in1118_2 = {pp58[40],c747,pp60[40],pp55[46]};
    CLA_4 KS_1118(s1118, c1118, in1118_1, in1118_2);
    wire[3:0] s1119, in1119_1, in1119_2;
    wire c1119;
    assign in1119_1 = {pp59[39],c748,pp61[39],pp56[45]};
    assign in1119_2 = {pp60[38],c749,pp62[38],pp57[44]};
    CLA_4 KS_1119(s1119, c1119, in1119_1, in1119_2);
    wire[3:0] s1120, in1120_1, in1120_2;
    wire c1120;
    assign in1120_1 = {pp61[37],c753,pp63[37],pp58[43]};
    assign in1120_2 = {pp62[36],c761,s764[1],pp59[42]};
    CLA_4 KS_1120(s1120, c1120, in1120_1, in1120_2);
    wire[3:0] s1121, in1121_1, in1121_2;
    wire c1121;
    assign in1121_1 = {pp63[35],s764[0],s765[1],pp60[41]};
    assign in1121_2 = {s743[3],s765[0],s766[1],pp61[40]};
    CLA_4 KS_1121(s1121, c1121, in1121_1, in1121_2);
    wire[3:0] s1122, in1122_1, in1122_2;
    wire c1122;
    assign in1122_1 = {s744[3],s766[0],s767[1],pp62[39]};
    assign in1122_2 = {s745[3],s767[0],s768[1],pp63[38]};
    CLA_4 KS_1122(s1122, c1122, in1122_1, in1122_2);
    wire[3:0] s1123, in1123_1, in1123_2;
    wire c1123;
    assign in1123_1 = {s746[3],s768[0],c769,s764[2]};
    assign in1123_2 = {s747[3],s769[0],s770[1],s765[2]};
    CLA_4 KS_1123(s1123, c1123, in1123_1, in1123_2);
    wire[3:0] s1124, in1124_1, in1124_2;
    wire c1124;
    assign in1124_1 = {s748[3],s770[0],c771,s766[2]};
    assign in1124_2 = {s749[3],s771[0],s772[1],s767[2]};
    CLA_4 KS_1124(s1124, c1124, in1124_1, in1124_2);
    wire[1:0] s1125, in1125_1, in1125_2;
    wire c1125;
    assign in1125_1 = {c750,s772[0]};
    assign in1125_2 = {s753[3],s773[0]};
    CLA_2 KS_1125(s1125, c1125, in1125_1, in1125_2);
    wire[0:0] s1126, in1126_1, in1126_2;
    wire c1126;
    assign in1126_1 = {c757};
    assign in1126_2 = {s761[3]};
    Half_Adder KS_1126(s1126, c1126, in1126_1, in1126_2);
    wire[3:0] s1127, in1127_1, in1127_2;
    wire c1127;
    assign in1127_1 = {c1097,s774[0],c773,c768};
    assign in1127_2 = {c1098,s775[0],s774[1],s770[2]};
    CLA_4 KS_1127(s1127, c1127, in1127_1, in1127_2);
    wire[0:0] s1128, in1128_1, in1128_2;
    wire c1128;
    assign in1128_1 = {c1099};
    assign in1128_2 = {c1100};
    Half_Adder KS_1128(s1128, c1128, in1128_1, in1128_2);
    wire[1:0] s1129, in1129_1, in1129_2;
    wire c1129;
    assign in1129_1 = {c1101,s776[0]};
    assign in1129_2 = {c1102,s1116[1]};
    CLA_2 KS_1129(s1129, c1129, in1129_1, in1129_2);
    wire[0:0] s1130, in1130_1, in1130_2;
    wire c1130;
    assign in1130_1 = {c1103};
    assign in1130_2 = {c1104};
    Half_Adder KS_1130(s1130, c1130, in1130_1, in1130_2);
    wire[2:0] s1131, in1131_1, in1131_2;
    wire c1131;
    assign in1131_1 = {c1105,s1117[1],c775};
    assign in1131_2 = {c1108,s1118[1],s776[1]};
    CLA_3 KS_1131(s1131, c1131, in1131_1, in1131_2);
    wire[0:0] s1132, in1132_1, in1132_2;
    wire c1132;
    assign in1132_1 = {s1117[0]};
    assign in1132_2 = {s1118[0]};
    Full_Adder KS_1132(s1132, c1132, in1132_1, in1132_2, s1116[0]);
    wire[3:0] s1133, in1133_1, in1133_2;
    wire c1133;
    assign in1133_1 = {pp47[55],pp49[54],pp45[59],pp44[61]};
    assign in1133_2 = {pp48[54],pp50[53],pp46[58],pp45[60]};
    CLA_4 KS_1133(s1133, c1133, in1133_1, in1133_2);
    wire[3:0] s1134, in1134_1, in1134_2;
    wire c1134;
    assign in1134_1 = {pp49[53],pp51[52],pp47[57],pp46[59]};
    assign in1134_2 = {pp50[52],pp52[51],pp48[56],pp47[58]};
    CLA_4 KS_1134(s1134, c1134, in1134_1, in1134_2);
    wire[3:0] s1135, in1135_1, in1135_2;
    wire c1135;
    assign in1135_1 = {pp51[51],pp53[50],pp49[55],pp48[57]};
    assign in1135_2 = {pp52[50],pp54[49],pp50[54],pp49[56]};
    CLA_4 KS_1135(s1135, c1135, in1135_1, in1135_2);
    wire[3:0] s1136, in1136_1, in1136_2;
    wire c1136;
    assign in1136_1 = {pp53[49],pp55[48],pp51[53],pp50[55]};
    assign in1136_2 = {pp54[48],pp56[47],pp52[52],pp51[54]};
    CLA_4 KS_1136(s1136, c1136, in1136_1, in1136_2);
    wire[3:0] s1137, in1137_1, in1137_2;
    wire c1137;
    assign in1137_1 = {pp55[47],pp57[46],pp53[51],pp52[53]};
    assign in1137_2 = {pp56[46],pp58[45],pp54[50],pp53[52]};
    CLA_4 KS_1137(s1137, c1137, in1137_1, in1137_2);
    wire[3:0] s1138, in1138_1, in1138_2;
    wire c1138;
    assign in1138_1 = {pp57[45],pp59[44],pp55[49],pp54[51]};
    assign in1138_2 = {pp58[44],pp60[43],pp56[48],pp55[50]};
    CLA_4 KS_1138(s1138, c1138, in1138_1, in1138_2);
    wire[3:0] s1139, in1139_1, in1139_2;
    wire c1139;
    assign in1139_1 = {pp59[43],pp61[42],pp57[47],pp56[49]};
    assign in1139_2 = {pp60[42],pp62[41],pp58[46],pp57[48]};
    CLA_4 KS_1139(s1139, c1139, in1139_1, in1139_2);
    wire[3:0] s1140, in1140_1, in1140_2;
    wire c1140;
    assign in1140_1 = {pp61[41],pp63[40],pp59[45],pp58[47]};
    assign in1140_2 = {pp62[40],c764,pp60[44],pp59[46]};
    CLA_4 KS_1140(s1140, c1140, in1140_1, in1140_2);
    wire[3:0] s1141, in1141_1, in1141_2;
    wire c1141;
    assign in1141_1 = {pp63[39],c765,pp61[43],pp60[45]};
    assign in1141_2 = {s764[3],c766,pp62[42],pp61[44]};
    CLA_4 KS_1141(s1141, c1141, in1141_1, in1141_2);
    wire[2:0] s1142, in1142_1, in1142_2;
    wire c1142;
    assign in1142_1 = {s765[3],c770,pp63[41]};
    assign in1142_2 = {s766[3],s777[0],s777[1]};
    CLA_3 KS_1142(s1142, c1142, in1142_1, in1142_2);
    wire[0:0] s1143, in1143_1, in1143_2;
    wire c1143;
    assign in1143_1 = {c767};
    assign in1143_2 = {s770[3]};
    Half_Adder KS_1143(s1143, c1143, in1143_1, in1143_2);
    wire[1:0] s1144, in1144_1, in1144_2;
    wire c1144;
    assign in1144_1 = {c774,s778[0]};
    assign in1144_2 = {c1116,s779[0]};
    CLA_2 KS_1144(s1144, c1144, in1144_1, in1144_2);
    wire[0:0] s1145, in1145_1, in1145_2;
    wire c1145;
    assign in1145_1 = {c1117};
    assign in1145_2 = {c1118};
    Half_Adder KS_1145(s1145, c1145, in1145_1, in1145_2);
    wire[3:0] s1146, in1146_1, in1146_2;
    wire c1146;
    assign in1146_1 = {c1119,s780[0],c778,pp62[43]};
    assign in1146_2 = {c1120,s1133[1],s779[1],pp63[42]};
    CLA_4 KS_1146(s1146, c1146, in1146_1, in1146_2);
    wire[0:0] s1147, in1147_1, in1147_2;
    wire c1147;
    assign in1147_1 = {c1121};
    assign in1147_2 = {c1122};
    Half_Adder KS_1147(s1147, c1147, in1147_1, in1147_2);
    wire[1:0] s1148, in1148_1, in1148_2;
    wire c1148;
    assign in1148_1 = {c1123,s1134[1]};
    assign in1148_2 = {c1124,s1135[1]};
    CLA_2 KS_1148(s1148, c1148, in1148_1, in1148_2);
    wire[0:0] s1149, in1149_1, in1149_2;
    wire c1149;
    assign in1149_1 = {c1127};
    assign in1149_2 = {s1133[0]};
    Half_Adder KS_1149(s1149, c1149, in1149_1, in1149_2);
    wire[2:0] s1150, in1150_1, in1150_2;
    wire c1150;
    assign in1150_1 = {s1135[0],s1136[1],c780};
    assign in1150_2 = {s1136[0],s1137[1],s1133[2]};
    CLA_3_c KS_1150(s1150, c1150, in1150_1, in1150_2, s1134[0]);
    wire[3:0] s1151, in1151_1, in1151_2;
    wire c1151;
    assign in1151_1 = {pp43[63],pp44[63],pp45[63],pp46[63]};
    assign in1151_2 = {pp44[62],pp45[62],pp46[62],pp47[62]};
    CLA_4 KS_1151(s1151, c1151, in1151_1, in1151_2);
    wire[3:0] s1152, in1152_1, in1152_2;
    wire c1152;
    assign in1152_1 = {pp45[61],pp46[61],pp47[61],pp48[61]};
    assign in1152_2 = {pp46[60],pp47[60],pp48[60],pp49[60]};
    CLA_4 KS_1152(s1152, c1152, in1152_1, in1152_2);
    wire[3:0] s1153, in1153_1, in1153_2;
    wire c1153;
    assign in1153_1 = {pp47[59],pp48[59],pp49[59],pp50[59]};
    assign in1153_2 = {pp48[58],pp49[58],pp50[58],pp51[58]};
    CLA_4 KS_1153(s1153, c1153, in1153_1, in1153_2);
    wire[3:0] s1154, in1154_1, in1154_2;
    wire c1154;
    assign in1154_1 = {pp49[57],pp50[57],pp51[57],pp52[57]};
    assign in1154_2 = {pp50[56],pp51[56],pp52[56],pp53[56]};
    CLA_4 KS_1154(s1154, c1154, in1154_1, in1154_2);
    wire[3:0] s1155, in1155_1, in1155_2;
    wire c1155;
    assign in1155_1 = {pp51[55],pp52[55],pp53[55],pp54[55]};
    assign in1155_2 = {pp52[54],pp53[54],pp54[54],pp55[54]};
    CLA_4 KS_1155(s1155, c1155, in1155_1, in1155_2);
    wire[2:0] s1156, in1156_1, in1156_2;
    wire c1156;
    assign in1156_1 = {pp53[53],pp54[53],pp55[53]};
    assign in1156_2 = {pp54[52],pp55[52],pp56[52]};
    CLA_3 KS_1156(s1156, c1156, in1156_1, in1156_2);
    wire[1:0] s1157, in1157_1, in1157_2;
    wire c1157;
    assign in1157_1 = {pp55[51],pp56[51]};
    assign in1157_2 = {pp56[50],pp57[50]};
    CLA_2 KS_1157(s1157, c1157, in1157_1, in1157_2);
    wire[0:0] s1158, in1158_1, in1158_2;
    wire c1158;
    assign in1158_1 = {pp57[49]};
    assign in1158_2 = {pp58[48]};
    Half_Adder KS_1158(s1158, c1158, in1158_1, in1158_2);
    wire[3:0] s1159, in1159_1, in1159_2;
    wire c1159;
    assign in1159_1 = {pp59[47],pp58[49],pp57[51],pp56[53]};
    assign in1159_2 = {pp60[46],pp59[48],pp58[50],pp57[52]};
    CLA_4 KS_1159(s1159, c1159, in1159_1, in1159_2);
    wire[0:0] s1160, in1160_1, in1160_2;
    wire c1160;
    assign in1160_1 = {pp61[45]};
    assign in1160_2 = {pp62[44]};
    Half_Adder KS_1160(s1160, c1160, in1160_1, in1160_2);
    wire[1:0] s1161, in1161_1, in1161_2;
    wire c1161;
    assign in1161_1 = {pp63[43],pp60[47]};
    assign in1161_2 = {c779,pp61[46]};
    CLA_2 KS_1161(s1161, c1161, in1161_1, in1161_2);
    wire[0:0] s1162, in1162_1, in1162_2;
    wire c1162;
    assign in1162_1 = {c1133};
    assign in1162_2 = {c1134};
    Half_Adder KS_1162(s1162, c1162, in1162_1, in1162_2);
    wire[2:0] s1163, in1163_1, in1163_2;
    wire c1163;
    assign in1163_1 = {c1135,pp62[45],pp59[49]};
    assign in1163_2 = {c1136,pp63[44],pp60[48]};
    CLA_3 KS_1163(s1163, c1163, in1163_1, in1163_2);
    wire[0:0] s1164, in1164_1, in1164_2;
    wire c1164;
    assign in1164_1 = {c1137};
    assign in1164_2 = {c1138};
    Half_Adder KS_1164(s1164, c1164, in1164_1, in1164_2);
    wire[1:0] s1165, in1165_1, in1165_2;
    wire c1165;
    assign in1165_1 = {c1139,s1151[1]};
    assign in1165_2 = {c1140,s1152[1]};
    CLA_2 KS_1165(s1165, c1165, in1165_1, in1165_2);
    wire[0:0] s1166, in1166_1, in1166_2;
    wire c1166;
    assign in1166_1 = {c1141};
    assign in1166_2 = {c1146};
    Half_Adder KS_1166(s1166, c1166, in1166_1, in1166_2);
    wire[3:0] s1167, in1167_1, in1167_2;
    wire c1167;
    assign in1167_1 = {s1152[0],s1153[1],pp61[47],pp58[51]};
    assign in1167_2 = {s1153[0],s1154[1],pp62[46],pp59[50]};
    CLA_4_c KS_1167(s1167, c1167, in1167_1, in1167_2, s1151[0]);
    wire[3:0] s1168, in1168_1, in1168_2;
    wire c1168;
    assign in1168_1 = {pp47[63],pp48[63],pp49[63],pp50[63]};
    assign in1168_2 = {pp48[62],pp49[62],pp50[62],pp51[62]};
    CLA_4 KS_1168(s1168, c1168, in1168_1, in1168_2);
    wire[2:0] s1169, in1169_1, in1169_2;
    wire c1169;
    assign in1169_1 = {pp49[61],pp50[61],pp51[61]};
    assign in1169_2 = {pp50[60],pp51[60],pp52[60]};
    CLA_3 KS_1169(s1169, c1169, in1169_1, in1169_2);
    wire[1:0] s1170, in1170_1, in1170_2;
    wire c1170;
    assign in1170_1 = {pp51[59],pp52[59]};
    assign in1170_2 = {pp52[58],pp53[58]};
    CLA_2 KS_1170(s1170, c1170, in1170_1, in1170_2);
    wire[0:0] s1171, in1171_1, in1171_2;
    wire c1171;
    assign in1171_1 = {pp53[57]};
    assign in1171_2 = {pp54[56]};
    Half_Adder KS_1171(s1171, c1171, in1171_1, in1171_2);
    wire[3:0] s1172, in1172_1, in1172_2;
    wire c1172;
    assign in1172_1 = {pp55[55],pp54[57],pp53[59],pp52[61]};
    assign in1172_2 = {pp56[54],pp55[56],pp54[58],pp53[60]};
    CLA_4 KS_1172(s1172, c1172, in1172_1, in1172_2);
    wire[0:0] s1173, in1173_1, in1173_2;
    wire c1173;
    assign in1173_1 = {pp57[53]};
    assign in1173_2 = {pp58[52]};
    Half_Adder KS_1173(s1173, c1173, in1173_1, in1173_2);
    wire[1:0] s1174, in1174_1, in1174_2;
    wire c1174;
    assign in1174_1 = {pp59[51],pp56[55]};
    assign in1174_2 = {pp60[50],pp57[54]};
    CLA_2 KS_1174(s1174, c1174, in1174_1, in1174_2);
    wire[0:0] s1175, in1175_1, in1175_2;
    wire c1175;
    assign in1175_1 = {pp61[49]};
    assign in1175_2 = {pp62[48]};
    Half_Adder KS_1175(s1175, c1175, in1175_1, in1175_2);
    wire[2:0] s1176, in1176_1, in1176_2;
    wire c1176;
    assign in1176_1 = {c1151,pp58[53],pp55[57]};
    assign in1176_2 = {c1152,pp59[52],pp56[56]};
    CLA_3_c KS_1176(s1176, c1176, in1176_1, in1176_2, pp63[47]);
    wire[0:0] s1177, in1177_1, in1177_2;
    wire c1177;
    assign in1177_1 = {pp51[63]};
    assign in1177_2 = {pp52[62]};
    Half_Adder KS_1177(s1177, c1177, in1177_1, in1177_2);

    /*Stage 4*/
    wire[3:0] s1178, in1178_1, in1178_2;
    wire c1178;
    assign in1178_1 = {pp0[9],pp0[10],pp0[11],pp0[12]};
    assign in1178_2 = {pp1[8],pp1[9],pp1[10],pp1[11]};
    CLA_4 KS_1178(s1178, c1178, in1178_1, in1178_2);
    wire[3:0] s1179, in1179_1, in1179_2;
    wire c1179;
    assign in1179_1 = {pp2[8],pp2[9],pp2[10],pp0[13]};
    assign in1179_2 = {pp3[7],pp3[8],pp3[9],pp1[12]};
    CLA_4 KS_1179(s1179, c1179, in1179_1, in1179_2);
    wire[3:0] s1180, in1180_1, in1180_2;
    wire c1180;
    assign in1180_1 = {pp4[7],pp4[8],pp2[11],pp2[12]};
    assign in1180_2 = {pp5[6],pp5[7],pp3[10],pp3[11]};
    CLA_4 KS_1180(s1180, c1180, in1180_1, in1180_2);
    wire[3:0] s1181, in1181_1, in1181_2;
    wire c1181;
    assign in1181_1 = {pp6[6],pp4[9],pp4[10],pp4[11]};
    assign in1181_2 = {pp7[5],pp5[8],pp5[9],pp5[10]};
    CLA_4 KS_1181(s1181, c1181, in1181_1, in1181_2);
    wire[3:0] s1182, in1182_1, in1182_2;
    wire c1182;
    assign in1182_1 = {pp6[7],pp6[8],pp6[9],pp6[10]};
    assign in1182_2 = {pp7[6],pp7[7],pp7[8],pp7[9]};
    CLA_4 KS_1182(s1182, c1182, in1182_1, in1182_2);
    wire[3:0] s1183, in1183_1, in1183_2;
    wire c1183;
    assign in1183_1 = {pp9[4],pp8[6],pp8[7],pp8[8]};
    assign in1183_2 = {pp10[3],pp9[5],pp9[6],pp9[7]};
    CLA_4_c KS_1183(s1183, c1183, in1183_1, in1183_2, pp8[5]);
    wire[3:0] s1184, in1184_1, in1184_2;
    wire c1184;
    assign in1184_1 = {pp11[3],pp10[5],pp10[6],pp8[9]};
    assign in1184_2 = {pp12[2],pp11[4],pp11[5],pp9[8]};
    CLA_4_c KS_1184(s1184, c1184, in1184_1, in1184_2, pp10[4]);
    wire[3:0] s1185, in1185_1, in1185_2;
    wire c1185;
    assign in1185_1 = {pp13[2],pp12[4],pp10[7],pp11[7]};
    assign in1185_2 = {pp14[1],pp13[3],pp11[6],pp12[6]};
    CLA_4_c KS_1185(s1185, c1185, in1185_1, in1185_2, pp12[3]);
    wire[3:0] s1186, in1186_1, in1186_2;
    wire c1186;
    assign in1186_1 = {pp15[1],pp12[5],pp13[5],pp13[6]};
    assign in1186_2 = {pp16[0],pp13[4],pp14[4],pp14[5]};
    CLA_4_c KS_1186(s1186, c1186, in1186_1, in1186_2, pp14[2]);
    wire[3:0] s1187, in1187_1, in1187_2;
    wire c1187;
    assign in1187_1 = {pp14[3],pp15[3],pp15[4],pp15[5]};
    assign in1187_2 = {pp15[2],pp16[2],pp16[3],pp16[4]};
    CLA_4 KS_1187(s1187, c1187, in1187_1, in1187_2);
    wire[3:0] s1188, in1188_1, in1188_2;
    wire c1188;
    assign in1188_1 = {pp16[1],pp17[1],pp17[2],pp17[3]};
    assign in1188_2 = {pp17[0],pp18[0],pp18[1],pp18[2]};
    CLA_4 KS_1188(s1188, c1188, in1188_1, in1188_2);
    wire[3:0] s1189, in1189_1, in1189_2;
    wire c1189;
    assign in1189_1 = {s782[2],c781,pp19[0],pp19[1]};
    assign in1189_2 = {s783[1],s782[3],c782,pp20[0]};
    CLA_4_c KS_1189(s1189, c1189, in1189_1, in1189_2, s781[3]);
    wire[3:0] s1190, in1190_1, in1190_2;
    wire c1190;
    assign in1190_1 = {s783[2],s783[3],c783,pp17[4]};
    assign in1190_2 = {s784[1],s784[2],s784[3],pp18[3]};
    CLA_4 KS_1190(s1190, c1190, in1190_1, in1190_2);
    wire[3:0] s1191, in1191_1, in1191_2;
    wire c1191;
    assign in1191_1 = {s785[1],s785[2],pp19[2],pp21[1]};
    assign in1191_2 = {s786[1],s786[2],pp20[1],pp22[0]};
    CLA_4 KS_1191(s1191, c1191, in1191_1, in1191_2);
    wire[3:0] s1192, in1192_1, in1192_2;
    wire c1192;
    assign in1192_1 = {s787[1],pp21[0],c785,pp23[0]};
    assign in1192_2 = {s788[1],c784,c786,s302[0]};
    CLA_4 KS_1192(s1192, c1192, in1192_1, in1192_2);
    wire[3:0] s1193, in1193_1, in1193_2;
    wire c1193;
    assign in1193_1 = {s785[3],s787[3],c787,s302[1]};
    assign in1193_2 = {s786[3],s788[3],c788,s303[0]};
    CLA_4 KS_1193(s1193, c1193, in1193_1, in1193_2);
    wire[3:0] s1194, in1194_1, in1194_2;
    wire c1194;
    assign in1194_1 = {s787[2],s789[2],s789[3],c789};
    assign in1194_2 = {s788[2],s790[2],s790[3],c790};
    CLA_4 KS_1194(s1194, c1194, in1194_1, in1194_2);
    wire[3:0] s1195, in1195_1, in1195_2;
    wire c1195;
    assign in1195_1 = {s789[1],s791[1],s791[2],s791[3]};
    assign in1195_2 = {s790[1],s792[1],s792[2],s792[3]};
    CLA_4 KS_1195(s1195, c1195, in1195_1, in1195_2);
    wire[3:0] s1196, in1196_1, in1196_2;
    wire c1196;
    assign in1196_1 = {s792[0],s793[0],s793[1],s793[2]};
    assign in1196_2 = {c1187,s794[0],s794[1],s794[2]};
    CLA_4_c KS_1196(s1196, c1196, in1196_1, in1196_2, s791[0]);
    wire[3:0] s1197, in1197_1, in1197_2;
    wire c1197;
    assign in1197_1 = {s795[1],s795[2],s303[1],c795};
    assign in1197_2 = {s796[1],s796[2],s304[0],c796};
    CLA_4 KS_1197(s1197, c1197, in1197_1, in1197_2);
    wire[3:0] s1198, in1198_1, in1198_2;
    wire c1198;
    assign in1198_1 = {s797[1],c791,s797[3],s307[0]};
    assign in1198_2 = {s798[1],c792,s798[3],c797};
    CLA_4 KS_1198(s1198, c1198, in1198_1, in1198_2);
    wire[3:0] s1199, in1199_1, in1199_2;
    wire c1199;
    assign in1199_1 = {s793[3],s799[2],c798,s308[0]};
    assign in1199_2 = {s794[3],s800[2],s799[3],s309[0]};
    CLA_4 KS_1199(s1199, c1199, in1199_1, in1199_2);
    wire[3:0] s1200, in1200_1, in1200_2;
    wire c1200;
    assign in1200_1 = {s795[3],s801[1],s800[3],c799};
    assign in1200_2 = {s796[3],s802[1],s801[2],c800};
    CLA_4 KS_1200(s1200, c1200, in1200_1, in1200_2);
    wire[3:0] s1201, in1201_1, in1201_2;
    wire c1201;
    assign in1201_1 = {s797[2],s803[0],s802[2],s801[3]};
    assign in1201_2 = {s798[2],s804[0],s803[1],s802[3]};
    CLA_4 KS_1201(s1201, c1201, in1201_1, in1201_2);
    wire[3:0] s1202, in1202_1, in1202_2;
    wire c1202;
    assign in1202_1 = {s799[1],s805[0],s804[1],s803[2]};
    assign in1202_2 = {s800[1],s806[0],s805[1],s804[2]};
    CLA_4 KS_1202(s1202, c1202, in1202_1, in1202_2);
    wire[0:0] s1203, in1203_1, in1203_2;
    wire c1203;
    assign in1203_1 = {s801[0]};
    assign in1203_2 = {s802[0]};
    Half_Adder KS_1203(s1203, c1203, in1203_1, in1203_2);
    wire[3:0] s1204, in1204_1, in1204_2;
    wire c1204;
    assign in1204_1 = {c1194,s807[0],s806[1],s805[2]};
    assign in1204_2 = {c1195,s808[0],s807[1],s806[2]};
    CLA_4_c KS_1204(s1204, c1204, in1204_1, in1204_2, c1193);
    wire[3:0] s1205, in1205_1, in1205_2;
    wire c1205;
    assign in1205_1 = {s807[2],s310[0],s809[3],s810[3]};
    assign in1205_2 = {s808[2],s311[0],s810[2],s811[2]};
    CLA_4 KS_1205(s1205, c1205, in1205_1, in1205_2);
    wire[3:0] s1206, in1206_1, in1206_2;
    wire c1206;
    assign in1206_1 = {c801,s811[1],s812[2],s320[0]};
    assign in1206_2 = {c802,s812[1],s813[1],c810};
    CLA_4 KS_1206(s1206, c1206, in1206_1, in1206_2);
    wire[3:0] s1207, in1207_1, in1207_2;
    wire c1207;
    assign in1207_1 = {s803[3],s813[0],s814[1],s811[3]};
    assign in1207_2 = {s804[3],s814[0],s815[1],s812[3]};
    CLA_4 KS_1207(s1207, c1207, in1207_1, in1207_2);
    wire[3:0] s1208, in1208_1, in1208_2;
    wire c1208;
    assign in1208_1 = {s805[3],s815[0],s816[1],s813[2]};
    assign in1208_2 = {s806[3],s816[0],s817[1],s814[2]};
    CLA_4 KS_1208(s1208, c1208, in1208_1, in1208_2);
    wire[3:0] s1209, in1209_1, in1209_2;
    wire c1209;
    assign in1209_1 = {s807[3],s817[0],s818[1],s815[2]};
    assign in1209_2 = {s808[3],s818[0],s819[1],s816[2]};
    CLA_4 KS_1209(s1209, c1209, in1209_1, in1209_2);
    wire[1:0] s1210, in1210_1, in1210_2;
    wire c1210;
    assign in1210_1 = {s809[2],s819[0]};
    assign in1210_2 = {s810[1],s820[0]};
    CLA_2 KS_1210(s1210, c1210, in1210_1, in1210_2);
    wire[0:0] s1211, in1211_1, in1211_2;
    wire c1211;
    assign in1211_1 = {s811[0]};
    assign in1211_2 = {s812[0]};
    Half_Adder KS_1211(s1211, c1211, in1211_1, in1211_2);
    wire[3:0] s1212, in1212_1, in1212_2;
    wire c1212;
    assign in1212_1 = {c1199,s821[0],s820[1],s817[2]};
    assign in1212_2 = {c1200,s822[0],c821,s818[2]};
    CLA_4 KS_1212(s1212, c1212, in1212_1, in1212_2);
    wire[0:0] s1213, in1213_1, in1213_2;
    wire c1213;
    assign in1213_1 = {c1202};
    assign in1213_2 = {c1204};
    Full_Adder KS_1213(s1213, c1213, in1213_1, in1213_2, c1201);
    wire[3:0] s1214, in1214_1, in1214_2;
    wire c1214;
    assign in1214_1 = {s322[0],s826[0],s826[1],s336[0]};
    assign in1214_2 = {s323[0],s827[0],s827[1],s823[3]};
    CLA_4 KS_1214(s1214, c1214, in1214_1, in1214_2);
    wire[3:0] s1215, in1215_1, in1215_2;
    wire c1215;
    assign in1215_1 = {c811,s828[0],s828[1],s824[2]};
    assign in1215_2 = {c812,s829[0],s829[1],s825[2]};
    CLA_4 KS_1215(s1215, c1215, in1215_1, in1215_2);
    wire[3:0] s1216, in1216_1, in1216_2;
    wire c1216;
    assign in1216_1 = {s813[3],s830[0],s830[1],s826[2]};
    assign in1216_2 = {s814[3],s831[0],s831[1],s827[2]};
    CLA_4 KS_1216(s1216, c1216, in1216_1, in1216_2);
    wire[3:0] s1217, in1217_1, in1217_2;
    wire c1217;
    assign in1217_1 = {s815[3],s832[0],s832[1],s828[2]};
    assign in1217_2 = {s816[3],s833[0],c833,s829[2]};
    CLA_4 KS_1217(s1217, c1217, in1217_1, in1217_2);
    wire[3:0] s1218, in1218_1, in1218_2;
    wire c1218;
    assign in1218_1 = {s817[3],s834[0],s834[1],s830[2]};
    assign in1218_2 = {s818[3],s835[0],c835,s831[2]};
    CLA_4 KS_1218(s1218, c1218, in1218_1, in1218_2);
    wire[3:0] s1219, in1219_1, in1219_2;
    wire c1219;
    assign in1219_1 = {s819[3],s836[0],s836[1],s832[2]};
    assign in1219_2 = {s820[3],s837[0],c837,c834};
    CLA_4 KS_1219(s1219, c1219, in1219_1, in1219_2);
    wire[0:0] s1220, in1220_1, in1220_2;
    wire c1220;
    assign in1220_1 = {s822[3]};
    assign in1220_2 = {s823[0]};
    Half_Adder KS_1220(s1220, c1220, in1220_1, in1220_2);
    wire[1:0] s1221, in1221_1, in1221_2;
    wire c1221;
    assign in1221_1 = {c1206,s838[0]};
    assign in1221_2 = {c1207,s839[0]};
    CLA_2 KS_1221(s1221, c1221, in1221_1, in1221_2);
    wire[0:0] s1222, in1222_1, in1222_2;
    wire c1222;
    assign in1222_1 = {c1209};
    assign in1222_2 = {c1212};
    Full_Adder KS_1222(s1222, c1222, in1222_1, in1222_2, c1208);
    wire[3:0] s1223, in1223_1, in1223_2;
    wire c1223;
    assign in1223_1 = {s338[0],s844[0],s845[1],s841[2]};
    assign in1223_2 = {s339[0],s845[0],s846[1],s842[2]};
    CLA_4 KS_1223(s1223, c1223, in1223_1, in1223_2);
    wire[3:0] s1224, in1224_1, in1224_2;
    wire c1224;
    assign in1224_1 = {s340[0],s846[0],s847[1],s843[2]};
    assign in1224_2 = {c823,s847[0],s848[1],s844[2]};
    CLA_4 KS_1224(s1224, c1224, in1224_1, in1224_2);
    wire[3:0] s1225, in1225_1, in1225_2;
    wire c1225;
    assign in1225_1 = {s824[3],s848[0],s849[1],s845[2]};
    assign in1225_2 = {s825[3],s849[0],c850,s846[2]};
    CLA_4 KS_1225(s1225, c1225, in1225_1, in1225_2);
    wire[3:0] s1226, in1226_1, in1226_2;
    wire c1226;
    assign in1226_1 = {s826[3],s850[0],s851[1],s847[2]};
    assign in1226_2 = {s827[3],s851[0],c852,s848[2]};
    CLA_4 KS_1226(s1226, c1226, in1226_1, in1226_2);
    wire[3:0] s1227, in1227_1, in1227_2;
    wire c1227;
    assign in1227_1 = {s828[3],s852[0],s853[1],s849[2]};
    assign in1227_2 = {s829[3],s853[0],c854,c851};
    CLA_4 KS_1227(s1227, c1227, in1227_1, in1227_2);
    wire[1:0] s1228, in1228_1, in1228_2;
    wire c1228;
    assign in1228_1 = {s830[3],s854[0]};
    assign in1228_2 = {s831[3],s855[0]};
    CLA_2 KS_1228(s1228, c1228, in1228_1, in1228_2);
    wire[0:0] s1229, in1229_1, in1229_2;
    wire c1229;
    assign in1229_1 = {s832[3]};
    assign in1229_2 = {s836[3]};
    Half_Adder KS_1229(s1229, c1229, in1229_1, in1229_2);
    wire[2:0] s1230, in1230_1, in1230_2;
    wire c1230;
    assign in1230_1 = {c1214,s856[0],s855[1]};
    assign in1230_2 = {c1215,s857[0],c856};
    CLA_3 KS_1230(s1230, c1230, in1230_1, in1230_2);
    wire[0:0] s1231, in1231_1, in1231_2;
    wire c1231;
    assign in1231_1 = {c1216};
    assign in1231_2 = {c1217};
    Half_Adder KS_1231(s1231, c1231, in1231_1, in1231_2);
    wire[1:0] s1232, in1232_1, in1232_2;
    wire c1232;
    assign in1232_1 = {c1219,s1223[1]};
    assign in1232_2 = {s1223[0],s1224[1]};
    CLA_2_c KS_1232(s1232, c1232, in1232_1, in1232_2, c1218);
    wire[3:0] s1233, in1233_1, in1233_2;
    wire c1233;
    assign in1233_1 = {s358[0],s863[0],s863[1],s859[2]};
    assign in1233_2 = {s840[3],s864[0],s864[1],s860[2]};
    CLA_4 KS_1233(s1233, c1233, in1233_1, in1233_2);
    wire[3:0] s1234, in1234_1, in1234_2;
    wire c1234;
    assign in1234_1 = {s841[3],s865[0],s865[1],s861[2]};
    assign in1234_2 = {s842[3],s866[0],s866[1],s862[2]};
    CLA_4 KS_1234(s1234, c1234, in1234_1, in1234_2);
    wire[3:0] s1235, in1235_1, in1235_2;
    wire c1235;
    assign in1235_1 = {s843[3],s867[0],s867[1],s863[2]};
    assign in1235_2 = {s844[3],s868[0],c868,s864[2]};
    CLA_4 KS_1235(s1235, c1235, in1235_1, in1235_2);
    wire[3:0] s1236, in1236_1, in1236_2;
    wire c1236;
    assign in1236_1 = {s845[3],s869[0],s869[1],s865[2]};
    assign in1236_2 = {s846[3],s870[0],c870,s866[2]};
    CLA_4 KS_1236(s1236, c1236, in1236_1, in1236_2);
    wire[3:0] s1237, in1237_1, in1237_2;
    wire c1237;
    assign in1237_1 = {s847[3],s871[0],s871[1],s867[2]};
    assign in1237_2 = {s848[3],s872[0],c872,c869};
    CLA_4 KS_1237(s1237, c1237, in1237_1, in1237_2);
    wire[2:0] s1238, in1238_1, in1238_2;
    wire c1238;
    assign in1238_1 = {s849[3],s873[0],s873[1]};
    assign in1238_2 = {c853,s874[0],c874};
    CLA_3 KS_1238(s1238, c1238, in1238_1, in1238_2);
    wire[0:0] s1239, in1239_1, in1239_2;
    wire c1239;
    assign in1239_1 = {s857[3]};
    assign in1239_2 = {c1223};
    Half_Adder KS_1239(s1239, c1239, in1239_1, in1239_2);
    wire[1:0] s1240, in1240_1, in1240_2;
    wire c1240;
    assign in1240_1 = {c1225,s875[0]};
    assign in1240_2 = {c1226,s876[0]};
    CLA_2_c KS_1240(s1240, c1240, in1240_1, in1240_2, c1224);
    wire[3:0] s1241, in1241_1, in1241_2;
    wire c1241;
    assign in1241_1 = {s381[0],s882[0],s882[1],s877[2]};
    assign in1241_2 = {s858[3],s883[0],s883[1],s878[2]};
    CLA_4 KS_1241(s1241, c1241, in1241_1, in1241_2);
    wire[3:0] s1242, in1242_1, in1242_2;
    wire c1242;
    assign in1242_1 = {s859[3],s884[0],s884[1],s879[2]};
    assign in1242_2 = {s860[3],s885[0],s885[1],s880[2]};
    CLA_4 KS_1242(s1242, c1242, in1242_1, in1242_2);
    wire[3:0] s1243, in1243_1, in1243_2;
    wire c1243;
    assign in1243_1 = {s861[3],s886[0],s886[1],s881[2]};
    assign in1243_2 = {s862[3],s887[0],c887,s882[2]};
    CLA_4 KS_1243(s1243, c1243, in1243_1, in1243_2);
    wire[3:0] s1244, in1244_1, in1244_2;
    wire c1244;
    assign in1244_1 = {s863[3],s888[0],s888[1],s883[2]};
    assign in1244_2 = {s864[3],s889[0],c889,s884[2]};
    CLA_4 KS_1244(s1244, c1244, in1244_1, in1244_2);
    wire[3:0] s1245, in1245_1, in1245_2;
    wire c1245;
    assign in1245_1 = {s865[3],s890[0],s890[1],s885[2]};
    assign in1245_2 = {s866[3],s891[0],c891,c886};
    CLA_4 KS_1245(s1245, c1245, in1245_1, in1245_2);
    wire[3:0] s1246, in1246_1, in1246_2;
    wire c1246;
    assign in1246_1 = {s867[3],s892[0],s892[1],s888[2]};
    assign in1246_2 = {c871,s893[0],c893,c890};
    CLA_4 KS_1246(s1246, c1246, in1246_1, in1246_2);
    wire[0:0] s1247, in1247_1, in1247_2;
    wire c1247;
    assign in1247_1 = {s875[3]};
    assign in1247_2 = {c1233};
    Half_Adder KS_1247(s1247, c1247, in1247_1, in1247_2);
    wire[1:0] s1248, in1248_1, in1248_2;
    wire c1248;
    assign in1248_1 = {c1235,s894[0]};
    assign in1248_2 = {c1236,s895[0]};
    CLA_2_c KS_1248(s1248, c1248, in1248_1, in1248_2, c1234);
    wire[3:0] s1249, in1249_1, in1249_2;
    wire c1249;
    assign in1249_1 = {c405,s900[0],s901[1],s897[2]};
    assign in1249_2 = {s407[2],s901[0],s902[1],s898[2]};
    CLA_4 KS_1249(s1249, c1249, in1249_1, in1249_2);
    wire[3:0] s1250, in1250_1, in1250_2;
    wire c1250;
    assign in1250_1 = {s877[3],s902[0],s903[1],s899[2]};
    assign in1250_2 = {s878[3],s903[0],s904[1],s900[2]};
    CLA_4 KS_1250(s1250, c1250, in1250_1, in1250_2);
    wire[3:0] s1251, in1251_1, in1251_2;
    wire c1251;
    assign in1251_1 = {s879[3],s904[0],s905[1],s901[2]};
    assign in1251_2 = {s880[3],s905[0],c906,s902[2]};
    CLA_4 KS_1251(s1251, c1251, in1251_1, in1251_2);
    wire[3:0] s1252, in1252_1, in1252_2;
    wire c1252;
    assign in1252_1 = {s881[3],s906[0],s907[1],s903[2]};
    assign in1252_2 = {s882[3],s907[0],c908,s904[2]};
    CLA_4 KS_1252(s1252, c1252, in1252_1, in1252_2);
    wire[3:0] s1253, in1253_1, in1253_2;
    wire c1253;
    assign in1253_1 = {s883[3],s908[0],s909[1],s905[2]};
    assign in1253_2 = {s884[3],s909[0],c910,c907};
    CLA_4 KS_1253(s1253, c1253, in1253_1, in1253_2);
    wire[1:0] s1254, in1254_1, in1254_2;
    wire c1254;
    assign in1254_1 = {s885[3],s910[0]};
    assign in1254_2 = {c888,s911[0]};
    CLA_2 KS_1254(s1254, c1254, in1254_1, in1254_2);
    wire[0:0] s1255, in1255_1, in1255_2;
    wire c1255;
    assign in1255_1 = {s892[3]};
    assign in1255_2 = {c1241};
    Half_Adder KS_1255(s1255, c1255, in1255_1, in1255_2);
    wire[2:0] s1256, in1256_1, in1256_2;
    wire c1256;
    assign in1256_1 = {c1242,s912[0],s911[1]};
    assign in1256_2 = {c1243,s913[0],c912};
    CLA_3 KS_1256(s1256, c1256, in1256_1, in1256_2);
    wire[0:0] s1257, in1257_1, in1257_2;
    wire c1257;
    assign in1257_1 = {c1245};
    assign in1257_2 = {c1246};
    Full_Adder KS_1257(s1257, c1257, in1257_1, in1257_2, c1244);
    wire[3:0] s1258, in1258_1, in1258_2;
    wire c1258;
    assign in1258_1 = {c437,s919[0],s919[1],s915[2]};
    assign in1258_2 = {s896[3],s920[0],s920[1],s916[2]};
    CLA_4 KS_1258(s1258, c1258, in1258_1, in1258_2);
    wire[3:0] s1259, in1259_1, in1259_2;
    wire c1259;
    assign in1259_1 = {s897[3],s921[0],s921[1],s917[2]};
    assign in1259_2 = {s898[3],s922[0],s922[1],s918[2]};
    CLA_4 KS_1259(s1259, c1259, in1259_1, in1259_2);
    wire[3:0] s1260, in1260_1, in1260_2;
    wire c1260;
    assign in1260_1 = {s899[3],s923[0],s923[1],s919[2]};
    assign in1260_2 = {s900[3],s924[0],c924,s920[2]};
    CLA_4 KS_1260(s1260, c1260, in1260_1, in1260_2);
    wire[3:0] s1261, in1261_1, in1261_2;
    wire c1261;
    assign in1261_1 = {s901[3],s925[0],s925[1],s921[2]};
    assign in1261_2 = {s902[3],s926[0],c926,s922[2]};
    CLA_4 KS_1261(s1261, c1261, in1261_1, in1261_2);
    wire[3:0] s1262, in1262_1, in1262_2;
    wire c1262;
    assign in1262_1 = {s903[3],s927[0],s927[1],s923[2]};
    assign in1262_2 = {s904[3],s928[0],c928,c925};
    CLA_4 KS_1262(s1262, c1262, in1262_1, in1262_2);
    wire[2:0] s1263, in1263_1, in1263_2;
    wire c1263;
    assign in1263_1 = {s905[3],s929[0],s929[1]};
    assign in1263_2 = {c909,s930[0],c930};
    CLA_3 KS_1263(s1263, c1263, in1263_1, in1263_2);
    wire[0:0] s1264, in1264_1, in1264_2;
    wire c1264;
    assign in1264_1 = {s913[3]};
    assign in1264_2 = {c1249};
    Half_Adder KS_1264(s1264, c1264, in1264_1, in1264_2);
    wire[1:0] s1265, in1265_1, in1265_2;
    wire c1265;
    assign in1265_1 = {c1251,s931[0]};
    assign in1265_2 = {c1252,s932[0]};
    CLA_2_c KS_1265(s1265, c1265, in1265_1, in1265_2, c1250);
    wire[3:0] s1266, in1266_1, in1266_2;
    wire c1266;
    assign in1266_1 = {c468,s938[0],s938[1],s934[2]};
    assign in1266_2 = {s914[3],s939[0],s939[1],s935[2]};
    CLA_4 KS_1266(s1266, c1266, in1266_1, in1266_2);
    wire[3:0] s1267, in1267_1, in1267_2;
    wire c1267;
    assign in1267_1 = {s915[3],s940[0],s940[1],s936[2]};
    assign in1267_2 = {s916[3],s941[0],s941[1],s937[2]};
    CLA_4 KS_1267(s1267, c1267, in1267_1, in1267_2);
    wire[3:0] s1268, in1268_1, in1268_2;
    wire c1268;
    assign in1268_1 = {s917[3],s942[0],s942[1],s938[2]};
    assign in1268_2 = {s918[3],s943[0],c943,s939[2]};
    CLA_4 KS_1268(s1268, c1268, in1268_1, in1268_2);
    wire[3:0] s1269, in1269_1, in1269_2;
    wire c1269;
    assign in1269_1 = {s919[3],s944[0],s944[1],s940[2]};
    assign in1269_2 = {s920[3],s945[0],c945,s941[2]};
    CLA_4 KS_1269(s1269, c1269, in1269_1, in1269_2);
    wire[3:0] s1270, in1270_1, in1270_2;
    wire c1270;
    assign in1270_1 = {s921[3],s946[0],s946[1],s942[2]};
    assign in1270_2 = {s922[3],s947[0],c947,c944};
    CLA_4 KS_1270(s1270, c1270, in1270_1, in1270_2);
    wire[2:0] s1271, in1271_1, in1271_2;
    wire c1271;
    assign in1271_1 = {s923[3],s948[0],s948[1]};
    assign in1271_2 = {c927,s949[0],c949};
    CLA_3 KS_1271(s1271, c1271, in1271_1, in1271_2);
    wire[0:0] s1272, in1272_1, in1272_2;
    wire c1272;
    assign in1272_1 = {s931[3]};
    assign in1272_2 = {c1258};
    Half_Adder KS_1272(s1272, c1272, in1272_1, in1272_2);
    wire[1:0] s1273, in1273_1, in1273_2;
    wire c1273;
    assign in1273_1 = {c1260,s950[0]};
    assign in1273_2 = {c1261,s951[0]};
    CLA_2_c KS_1273(s1273, c1273, in1273_1, in1273_2, c1259);
    wire[3:0] s1274, in1274_1, in1274_2;
    wire c1274;
    assign in1274_1 = {c499,s957[0],s957[1],s952[2]};
    assign in1274_2 = {s933[3],s958[0],s958[1],s953[2]};
    CLA_4 KS_1274(s1274, c1274, in1274_1, in1274_2);
    wire[3:0] s1275, in1275_1, in1275_2;
    wire c1275;
    assign in1275_1 = {s934[3],s959[0],s959[1],s954[2]};
    assign in1275_2 = {s935[3],s960[0],s960[1],s955[2]};
    CLA_4 KS_1275(s1275, c1275, in1275_1, in1275_2);
    wire[3:0] s1276, in1276_1, in1276_2;
    wire c1276;
    assign in1276_1 = {s936[3],s961[0],s961[1],s956[2]};
    assign in1276_2 = {s937[3],s962[0],c962,s957[2]};
    CLA_4 KS_1276(s1276, c1276, in1276_1, in1276_2);
    wire[3:0] s1277, in1277_1, in1277_2;
    wire c1277;
    assign in1277_1 = {s938[3],s963[0],s963[1],s958[2]};
    assign in1277_2 = {s939[3],s964[0],c964,s959[2]};
    CLA_4 KS_1277(s1277, c1277, in1277_1, in1277_2);
    wire[3:0] s1278, in1278_1, in1278_2;
    wire c1278;
    assign in1278_1 = {s940[3],s965[0],s965[1],s960[2]};
    assign in1278_2 = {s941[3],s966[0],c966,c961};
    CLA_4 KS_1278(s1278, c1278, in1278_1, in1278_2);
    wire[3:0] s1279, in1279_1, in1279_2;
    wire c1279;
    assign in1279_1 = {s942[3],s967[0],s967[1],s963[2]};
    assign in1279_2 = {c946,s968[0],c968,c965};
    CLA_4 KS_1279(s1279, c1279, in1279_1, in1279_2);
    wire[0:0] s1280, in1280_1, in1280_2;
    wire c1280;
    assign in1280_1 = {s950[3]};
    assign in1280_2 = {c1266};
    Half_Adder KS_1280(s1280, c1280, in1280_1, in1280_2);
    wire[1:0] s1281, in1281_1, in1281_2;
    wire c1281;
    assign in1281_1 = {c1268,s969[0]};
    assign in1281_2 = {c1269,s970[0]};
    CLA_2_c KS_1281(s1281, c1281, in1281_1, in1281_2, c1267);
    wire[3:0] s1282, in1282_1, in1282_2;
    wire c1282;
    assign in1282_1 = {c526,s975[0],s976[1],s972[2]};
    assign in1282_2 = {s528[2],s976[0],s977[1],s973[2]};
    CLA_4 KS_1282(s1282, c1282, in1282_1, in1282_2);
    wire[3:0] s1283, in1283_1, in1283_2;
    wire c1283;
    assign in1283_1 = {c530,s977[0],s978[1],s974[2]};
    assign in1283_2 = {s952[3],s978[0],s979[1],s975[2]};
    CLA_4 KS_1283(s1283, c1283, in1283_1, in1283_2);
    wire[3:0] s1284, in1284_1, in1284_2;
    wire c1284;
    assign in1284_1 = {s953[3],s979[0],s980[1],s976[2]};
    assign in1284_2 = {s954[3],s980[0],c981,s977[2]};
    CLA_4 KS_1284(s1284, c1284, in1284_1, in1284_2);
    wire[3:0] s1285, in1285_1, in1285_2;
    wire c1285;
    assign in1285_1 = {s955[3],s981[0],s982[1],s978[2]};
    assign in1285_2 = {s956[3],s982[0],c983,s979[2]};
    CLA_4 KS_1285(s1285, c1285, in1285_1, in1285_2);
    wire[3:0] s1286, in1286_1, in1286_2;
    wire c1286;
    assign in1286_1 = {s957[3],s983[0],s984[1],s980[2]};
    assign in1286_2 = {s958[3],s984[0],c985,c982};
    CLA_4 KS_1286(s1286, c1286, in1286_1, in1286_2);
    wire[1:0] s1287, in1287_1, in1287_2;
    wire c1287;
    assign in1287_1 = {s959[3],s985[0]};
    assign in1287_2 = {s960[3],s986[0]};
    CLA_2 KS_1287(s1287, c1287, in1287_1, in1287_2);
    wire[0:0] s1288, in1288_1, in1288_2;
    wire c1288;
    assign in1288_1 = {s963[3]};
    assign in1288_2 = {c967};
    Half_Adder KS_1288(s1288, c1288, in1288_1, in1288_2);
    wire[2:0] s1289, in1289_1, in1289_2;
    wire c1289;
    assign in1289_1 = {c1274,s987[0],s986[1]};
    assign in1289_2 = {c1275,s988[0],c987};
    CLA_3 KS_1289(s1289, c1289, in1289_1, in1289_2);
    wire[0:0] s1290, in1290_1, in1290_2;
    wire c1290;
    assign in1290_1 = {c1276};
    assign in1290_2 = {c1277};
    Half_Adder KS_1290(s1290, c1290, in1290_1, in1290_2);
    wire[1:0] s1291, in1291_1, in1291_2;
    wire c1291;
    assign in1291_1 = {c1279,s1282[1]};
    assign in1291_2 = {s1282[0],s1283[1]};
    CLA_2_c KS_1291(s1291, c1291, in1291_1, in1291_2, c1278);
    wire[3:0] s1292, in1292_1, in1292_2;
    wire c1292;
    assign in1292_1 = {c557,s993[0],s994[1],s990[2]};
    assign in1292_2 = {s559[2],s994[0],s995[1],s991[2]};
    CLA_4 KS_1292(s1292, c1292, in1292_1, in1292_2);
    wire[3:0] s1293, in1293_1, in1293_2;
    wire c1293;
    assign in1293_1 = {s971[3],s995[0],s996[1],s992[2]};
    assign in1293_2 = {s972[3],s996[0],s997[1],s993[2]};
    CLA_4 KS_1293(s1293, c1293, in1293_1, in1293_2);
    wire[3:0] s1294, in1294_1, in1294_2;
    wire c1294;
    assign in1294_1 = {s973[3],s997[0],s998[1],s994[2]};
    assign in1294_2 = {s974[3],s998[0],c999,s995[2]};
    CLA_4 KS_1294(s1294, c1294, in1294_1, in1294_2);
    wire[3:0] s1295, in1295_1, in1295_2;
    wire c1295;
    assign in1295_1 = {s975[3],s999[0],s1000[1],s996[2]};
    assign in1295_2 = {s976[3],s1000[0],c1001,s997[2]};
    CLA_4 KS_1295(s1295, c1295, in1295_1, in1295_2);
    wire[3:0] s1296, in1296_1, in1296_2;
    wire c1296;
    assign in1296_1 = {s977[3],s1001[0],s1002[1],s998[2]};
    assign in1296_2 = {s978[3],s1002[0],c1003,c1000};
    CLA_4 KS_1296(s1296, c1296, in1296_1, in1296_2);
    wire[1:0] s1297, in1297_1, in1297_2;
    wire c1297;
    assign in1297_1 = {s979[3],s1003[0]};
    assign in1297_2 = {c980,s1004[0]};
    CLA_2 KS_1297(s1297, c1297, in1297_1, in1297_2);
    wire[0:0] s1298, in1298_1, in1298_2;
    wire c1298;
    assign in1298_1 = {s984[3]};
    assign in1298_2 = {c988};
    Half_Adder KS_1298(s1298, c1298, in1298_1, in1298_2);
    wire[2:0] s1299, in1299_1, in1299_2;
    wire c1299;
    assign in1299_1 = {c1282,s1005[0],s1004[1]};
    assign in1299_2 = {c1283,s1006[0],c1005};
    CLA_3 KS_1299(s1299, c1299, in1299_1, in1299_2);
    wire[0:0] s1300, in1300_1, in1300_2;
    wire c1300;
    assign in1300_1 = {c1285};
    assign in1300_2 = {c1286};
    Full_Adder KS_1300(s1300, c1300, in1300_1, in1300_2, c1284);
    wire[3:0] s1301, in1301_1, in1301_2;
    wire c1301;
    assign in1301_1 = {c587,s1011[0],s1012[1],s1007[2]};
    assign in1301_2 = {s589[2],s1012[0],s1013[1],s1008[2]};
    CLA_4 KS_1301(s1301, c1301, in1301_1, in1301_2);
    wire[3:0] s1302, in1302_1, in1302_2;
    wire c1302;
    assign in1302_1 = {s989[3],s1013[0],s1014[1],s1009[2]};
    assign in1302_2 = {s990[3],s1014[0],s1015[1],s1010[2]};
    CLA_4 KS_1302(s1302, c1302, in1302_1, in1302_2);
    wire[3:0] s1303, in1303_1, in1303_2;
    wire c1303;
    assign in1303_1 = {s991[3],s1015[0],s1016[1],s1011[2]};
    assign in1303_2 = {s992[3],s1016[0],c1017,s1012[2]};
    CLA_4 KS_1303(s1303, c1303, in1303_1, in1303_2);
    wire[3:0] s1304, in1304_1, in1304_2;
    wire c1304;
    assign in1304_1 = {s993[3],s1017[0],s1018[1],s1013[2]};
    assign in1304_2 = {s994[3],s1018[0],c1019,s1014[2]};
    CLA_4 KS_1304(s1304, c1304, in1304_1, in1304_2);
    wire[3:0] s1305, in1305_1, in1305_2;
    wire c1305;
    assign in1305_1 = {s995[3],s1019[0],s1020[1],s1015[2]};
    assign in1305_2 = {s996[3],s1020[0],c1021,c1016};
    CLA_4 KS_1305(s1305, c1305, in1305_1, in1305_2);
    wire[1:0] s1306, in1306_1, in1306_2;
    wire c1306;
    assign in1306_1 = {s997[3],s1021[0]};
    assign in1306_2 = {c998,s1022[0]};
    CLA_2 KS_1306(s1306, c1306, in1306_1, in1306_2);
    wire[0:0] s1307, in1307_1, in1307_2;
    wire c1307;
    assign in1307_1 = {s1002[3]};
    assign in1307_2 = {c1006};
    Half_Adder KS_1307(s1307, c1307, in1307_1, in1307_2);
    wire[3:0] s1308, in1308_1, in1308_2;
    wire c1308;
    assign in1308_1 = {c1292,s1023[0],s1022[1],s1018[2]};
    assign in1308_2 = {c1293,s1024[0],c1023,c1020};
    CLA_4 KS_1308(s1308, c1308, in1308_1, in1308_2);
    wire[0:0] s1309, in1309_1, in1309_2;
    wire c1309;
    assign in1309_1 = {c1295};
    assign in1309_2 = {c1296};
    Full_Adder KS_1309(s1309, c1309, in1309_1, in1309_2, c1294);
    wire[3:0] s1310, in1310_1, in1310_2;
    wire c1310;
    assign in1310_1 = {c619,s1029[0],s1030[1],s1025[2]};
    assign in1310_2 = {s621[2],s1030[0],s1031[1],s1026[2]};
    CLA_4 KS_1310(s1310, c1310, in1310_1, in1310_2);
    wire[3:0] s1311, in1311_1, in1311_2;
    wire c1311;
    assign in1311_1 = {s1007[3],s1031[0],s1032[1],s1027[2]};
    assign in1311_2 = {s1008[3],s1032[0],s1033[1],s1028[2]};
    CLA_4 KS_1311(s1311, c1311, in1311_1, in1311_2);
    wire[3:0] s1312, in1312_1, in1312_2;
    wire c1312;
    assign in1312_1 = {s1009[3],s1033[0],s1034[1],s1029[2]};
    assign in1312_2 = {s1010[3],s1034[0],c1035,s1030[2]};
    CLA_4 KS_1312(s1312, c1312, in1312_1, in1312_2);
    wire[3:0] s1313, in1313_1, in1313_2;
    wire c1313;
    assign in1313_1 = {s1011[3],s1035[0],s1036[1],s1031[2]};
    assign in1313_2 = {s1012[3],s1036[0],c1037,s1032[2]};
    CLA_4 KS_1313(s1313, c1313, in1313_1, in1313_2);
    wire[3:0] s1314, in1314_1, in1314_2;
    wire c1314;
    assign in1314_1 = {s1013[3],s1037[0],s1038[1],s1033[2]};
    assign in1314_2 = {s1014[3],s1038[0],c1039,c1034};
    CLA_4 KS_1314(s1314, c1314, in1314_1, in1314_2);
    wire[1:0] s1315, in1315_1, in1315_2;
    wire c1315;
    assign in1315_1 = {s1015[3],s1039[0]};
    assign in1315_2 = {c1018,s1040[0]};
    CLA_2 KS_1315(s1315, c1315, in1315_1, in1315_2);
    wire[0:0] s1316, in1316_1, in1316_2;
    wire c1316;
    assign in1316_1 = {s1022[3]};
    assign in1316_2 = {c1301};
    Half_Adder KS_1316(s1316, c1316, in1316_1, in1316_2);
    wire[3:0] s1317, in1317_1, in1317_2;
    wire c1317;
    assign in1317_1 = {c1302,s1041[0],s1040[1],s1036[2]};
    assign in1317_2 = {c1303,s1042[0],c1041,c1038};
    CLA_4 KS_1317(s1317, c1317, in1317_1, in1317_2);
    wire[0:0] s1318, in1318_1, in1318_2;
    wire c1318;
    assign in1318_1 = {c1305};
    assign in1318_2 = {c1308};
    Full_Adder KS_1318(s1318, c1318, in1318_1, in1318_2, c1304);
    wire[3:0] s1319, in1319_1, in1319_2;
    wire c1319;
    assign in1319_1 = {c648,s1047[0],s1048[1],s1044[2]};
    assign in1319_2 = {s650[2],s1048[0],s1049[1],s1045[2]};
    CLA_4 KS_1319(s1319, c1319, in1319_1, in1319_2);
    wire[3:0] s1320, in1320_1, in1320_2;
    wire c1320;
    assign in1320_1 = {c652,s1049[0],s1050[1],s1046[2]};
    assign in1320_2 = {s1025[3],s1050[0],s1051[1],s1047[2]};
    CLA_4 KS_1320(s1320, c1320, in1320_1, in1320_2);
    wire[3:0] s1321, in1321_1, in1321_2;
    wire c1321;
    assign in1321_1 = {s1026[3],s1051[0],s1052[1],s1048[2]};
    assign in1321_2 = {s1027[3],s1052[0],c1053,s1049[2]};
    CLA_4 KS_1321(s1321, c1321, in1321_1, in1321_2);
    wire[3:0] s1322, in1322_1, in1322_2;
    wire c1322;
    assign in1322_1 = {s1028[3],s1053[0],s1054[1],s1050[2]};
    assign in1322_2 = {s1029[3],s1054[0],c1055,s1051[2]};
    CLA_4 KS_1322(s1322, c1322, in1322_1, in1322_2);
    wire[3:0] s1323, in1323_1, in1323_2;
    wire c1323;
    assign in1323_1 = {s1030[3],s1055[0],s1056[1],s1052[2]};
    assign in1323_2 = {s1031[3],s1056[0],c1057,c1054};
    CLA_4 KS_1323(s1323, c1323, in1323_1, in1323_2);
    wire[1:0] s1324, in1324_1, in1324_2;
    wire c1324;
    assign in1324_1 = {s1032[3],s1057[0]};
    assign in1324_2 = {s1033[3],s1058[0]};
    CLA_2 KS_1324(s1324, c1324, in1324_1, in1324_2);
    wire[0:0] s1325, in1325_1, in1325_2;
    wire c1325;
    assign in1325_1 = {s1036[3]};
    assign in1325_2 = {c1040};
    Half_Adder KS_1325(s1325, c1325, in1325_1, in1325_2);
    wire[2:0] s1326, in1326_1, in1326_2;
    wire c1326;
    assign in1326_1 = {c1310,s1059[0],s1058[1]};
    assign in1326_2 = {c1311,s1060[0],c1059};
    CLA_3 KS_1326(s1326, c1326, in1326_1, in1326_2);
    wire[0:0] s1327, in1327_1, in1327_2;
    wire c1327;
    assign in1327_1 = {c1312};
    assign in1327_2 = {c1313};
    Half_Adder KS_1327(s1327, c1327, in1327_1, in1327_2);
    wire[1:0] s1328, in1328_1, in1328_2;
    wire c1328;
    assign in1328_1 = {c1317,s1319[1]};
    assign in1328_2 = {s1319[0],s1320[1]};
    CLA_2_c KS_1328(s1328, c1328, in1328_1, in1328_2, c1314);
    wire[3:0] s1329, in1329_1, in1329_2;
    wire c1329;
    assign in1329_1 = {c681,s1065[0],s1066[1],s1062[2]};
    assign in1329_2 = {s1043[3],s1066[0],s1067[1],s1063[2]};
    CLA_4 KS_1329(s1329, c1329, in1329_1, in1329_2);
    wire[3:0] s1330, in1330_1, in1330_2;
    wire c1330;
    assign in1330_1 = {s1044[3],s1067[0],s1068[1],s1064[2]};
    assign in1330_2 = {s1045[3],s1068[0],s1069[1],s1065[2]};
    CLA_4 KS_1330(s1330, c1330, in1330_1, in1330_2);
    wire[3:0] s1331, in1331_1, in1331_2;
    wire c1331;
    assign in1331_1 = {s1046[3],s1069[0],s1070[1],s1066[2]};
    assign in1331_2 = {s1047[3],s1070[0],c1071,s1067[2]};
    CLA_4 KS_1331(s1331, c1331, in1331_1, in1331_2);
    wire[3:0] s1332, in1332_1, in1332_2;
    wire c1332;
    assign in1332_1 = {s1048[3],s1071[0],s1072[1],s1068[2]};
    assign in1332_2 = {s1049[3],s1072[0],c1073,s1069[2]};
    CLA_4 KS_1332(s1332, c1332, in1332_1, in1332_2);
    wire[3:0] s1333, in1333_1, in1333_2;
    wire c1333;
    assign in1333_1 = {s1050[3],s1073[0],s1074[1],s1070[2]};
    assign in1333_2 = {s1051[3],s1074[0],c1075,c1072};
    CLA_4 KS_1333(s1333, c1333, in1333_1, in1333_2);
    wire[1:0] s1334, in1334_1, in1334_2;
    wire c1334;
    assign in1334_1 = {s1052[3],s1075[0]};
    assign in1334_2 = {c1056,s1076[0]};
    CLA_2 KS_1334(s1334, c1334, in1334_1, in1334_2);
    wire[0:0] s1335, in1335_1, in1335_2;
    wire c1335;
    assign in1335_1 = {s1060[3]};
    assign in1335_2 = {c1319};
    Half_Adder KS_1335(s1335, c1335, in1335_1, in1335_2);
    wire[2:0] s1336, in1336_1, in1336_2;
    wire c1336;
    assign in1336_1 = {c1321,s1077[0],s1076[1]};
    assign in1336_2 = {c1322,s1078[0],c1077};
    CLA_3_c KS_1336(s1336, c1336, in1336_1, in1336_2, c1320);
    wire[3:0] s1337, in1337_1, in1337_2;
    wire c1337;
    assign in1337_1 = {c709,s1083[0],s1084[1],s1080[2]};
    assign in1337_2 = {s711[2],s1084[0],s1085[1],s1081[2]};
    CLA_4 KS_1337(s1337, c1337, in1337_1, in1337_2);
    wire[3:0] s1338, in1338_1, in1338_2;
    wire c1338;
    assign in1338_1 = {s1061[3],s1085[0],s1086[1],s1082[2]};
    assign in1338_2 = {s1062[3],s1086[0],s1087[1],s1083[2]};
    CLA_4 KS_1338(s1338, c1338, in1338_1, in1338_2);
    wire[3:0] s1339, in1339_1, in1339_2;
    wire c1339;
    assign in1339_1 = {s1063[3],s1087[0],s1088[1],s1084[2]};
    assign in1339_2 = {s1064[3],s1088[0],c1089,s1085[2]};
    CLA_4 KS_1339(s1339, c1339, in1339_1, in1339_2);
    wire[3:0] s1340, in1340_1, in1340_2;
    wire c1340;
    assign in1340_1 = {s1065[3],s1089[0],s1090[1],s1086[2]};
    assign in1340_2 = {s1066[3],s1090[0],c1091,s1087[2]};
    CLA_4 KS_1340(s1340, c1340, in1340_1, in1340_2);
    wire[3:0] s1341, in1341_1, in1341_2;
    wire c1341;
    assign in1341_1 = {s1067[3],s1091[0],s1092[1],s1088[2]};
    assign in1341_2 = {s1068[3],s1092[0],c1093,c1090};
    CLA_4 KS_1341(s1341, c1341, in1341_1, in1341_2);
    wire[1:0] s1342, in1342_1, in1342_2;
    wire c1342;
    assign in1342_1 = {s1069[3],s1093[0]};
    assign in1342_2 = {c1070,s1094[0]};
    CLA_2 KS_1342(s1342, c1342, in1342_1, in1342_2);
    wire[0:0] s1343, in1343_1, in1343_2;
    wire c1343;
    assign in1343_1 = {s1074[3]};
    assign in1343_2 = {c1078};
    Half_Adder KS_1343(s1343, c1343, in1343_1, in1343_2);
    wire[2:0] s1344, in1344_1, in1344_2;
    wire c1344;
    assign in1344_1 = {c1329,s1095[0],s1094[1]};
    assign in1344_2 = {c1330,s1096[0],c1095};
    CLA_3 KS_1344(s1344, c1344, in1344_1, in1344_2);
    wire[0:0] s1345, in1345_1, in1345_2;
    wire c1345;
    assign in1345_1 = {c1332};
    assign in1345_2 = {c1333};
    Full_Adder KS_1345(s1345, c1345, in1345_1, in1345_2, c1331);
    wire[3:0] s1346, in1346_1, in1346_2;
    wire c1346;
    assign in1346_1 = {c741,s1102[0],s1102[1],s1097[2]};
    assign in1346_2 = {s1079[3],s1103[0],s1103[1],s1098[2]};
    CLA_4 KS_1346(s1346, c1346, in1346_1, in1346_2);
    wire[3:0] s1347, in1347_1, in1347_2;
    wire c1347;
    assign in1347_1 = {s1080[3],s1104[0],s1104[1],s1099[2]};
    assign in1347_2 = {s1081[3],s1105[0],s1105[1],s1100[2]};
    CLA_4 KS_1347(s1347, c1347, in1347_1, in1347_2);
    wire[3:0] s1348, in1348_1, in1348_2;
    wire c1348;
    assign in1348_1 = {s1082[3],s1106[0],s1106[1],s1101[2]};
    assign in1348_2 = {s1083[3],s1107[0],c1107,s1102[2]};
    CLA_4 KS_1348(s1348, c1348, in1348_1, in1348_2);
    wire[3:0] s1349, in1349_1, in1349_2;
    wire c1349;
    assign in1349_1 = {s1084[3],s1108[0],s1108[1],s1103[2]};
    assign in1349_2 = {s1085[3],s1109[0],c1109,s1104[2]};
    CLA_4 KS_1349(s1349, c1349, in1349_1, in1349_2);
    wire[3:0] s1350, in1350_1, in1350_2;
    wire c1350;
    assign in1350_1 = {s1086[3],s1110[0],s1110[1],s1105[2]};
    assign in1350_2 = {s1087[3],s1111[0],c1111,c1106};
    CLA_4 KS_1350(s1350, c1350, in1350_1, in1350_2);
    wire[3:0] s1351, in1351_1, in1351_2;
    wire c1351;
    assign in1351_1 = {s1088[3],s1112[0],s1112[1],s1108[2]};
    assign in1351_2 = {c1092,s1113[0],c1113,c1110};
    CLA_4 KS_1351(s1351, c1351, in1351_1, in1351_2);
    wire[0:0] s1352, in1352_1, in1352_2;
    wire c1352;
    assign in1352_1 = {s1096[3]};
    assign in1352_2 = {c1337};
    Half_Adder KS_1352(s1352, c1352, in1352_1, in1352_2);
    wire[1:0] s1353, in1353_1, in1353_2;
    wire c1353;
    assign in1353_1 = {c1339,s1114[0]};
    assign in1353_2 = {c1340,s1115[0]};
    CLA_2_c KS_1353(s1353, c1353, in1353_1, in1353_2, c1338);
    wire[3:0] s1354, in1354_1, in1354_2;
    wire c1354;
    assign in1354_1 = {c759,s1119[0],s1119[1],s1116[2]};
    assign in1354_2 = {s761[2],s1120[0],s1120[1],s1117[2]};
    CLA_4 KS_1354(s1354, c1354, in1354_1, in1354_2);
    wire[3:0] s1355, in1355_1, in1355_2;
    wire c1355;
    assign in1355_1 = {c763,s1121[0],s1121[1],s1118[2]};
    assign in1355_2 = {s1097[3],s1122[0],s1122[1],s1119[2]};
    CLA_4 KS_1355(s1355, c1355, in1355_1, in1355_2);
    wire[3:0] s1356, in1356_1, in1356_2;
    wire c1356;
    assign in1356_1 = {s1098[3],s1123[0],s1123[1],s1120[2]};
    assign in1356_2 = {s1099[3],s1124[0],s1124[1],s1121[2]};
    CLA_4 KS_1356(s1356, c1356, in1356_1, in1356_2);
    wire[3:0] s1357, in1357_1, in1357_2;
    wire c1357;
    assign in1357_1 = {s1100[3],s1125[0],s1125[1],s1122[2]};
    assign in1357_2 = {s1101[3],s1126[0],c1126,s1123[2]};
    CLA_4 KS_1357(s1357, c1357, in1357_1, in1357_2);
    wire[3:0] s1358, in1358_1, in1358_2;
    wire c1358;
    assign in1358_1 = {s1102[3],s1127[0],s1127[1],s1124[2]};
    assign in1358_2 = {s1103[3],s1128[0],c1128,c1125};
    CLA_4 KS_1358(s1358, c1358, in1358_1, in1358_2);
    wire[2:0] s1359, in1359_1, in1359_2;
    wire c1359;
    assign in1359_1 = {s1104[3],s1129[0],s1129[1]};
    assign in1359_2 = {s1105[3],s1130[0],c1130};
    CLA_3 KS_1359(s1359, c1359, in1359_1, in1359_2);
    wire[0:0] s1360, in1360_1, in1360_2;
    wire c1360;
    assign in1360_1 = {s1108[3]};
    assign in1360_2 = {c1112};
    Half_Adder KS_1360(s1360, c1360, in1360_1, in1360_2);
    wire[1:0] s1361, in1361_1, in1361_2;
    wire c1361;
    assign in1361_1 = {c1346,s1131[0]};
    assign in1361_2 = {c1347,s1132[0]};
    CLA_2 KS_1361(s1361, c1361, in1361_1, in1361_2);
    wire[0:0] s1362, in1362_1, in1362_2;
    wire c1362;
    assign in1362_1 = {c1348};
    assign in1362_2 = {c1349};
    Half_Adder KS_1362(s1362, c1362, in1362_1, in1362_2);
    wire[3:0] s1363, in1363_1, in1363_2;
    wire c1363;
    assign in1363_1 = {c1351,s1354[1],s1131[1],s1127[2]};
    assign in1363_2 = {s1354[0],s1355[1],c1132,c1129};
    CLA_4_c KS_1363(s1363, c1363, in1363_1, in1363_2, c1350);
    wire[3:0] s1364, in1364_1, in1364_2;
    wire c1364;
    assign in1364_1 = {c772,s1137[0],s1138[1],s1134[2]};
    assign in1364_2 = {s774[2],s1138[0],s1139[1],s1135[2]};
    CLA_4 KS_1364(s1364, c1364, in1364_1, in1364_2);
    wire[3:0] s1365, in1365_1, in1365_2;
    wire c1365;
    assign in1365_1 = {c776,s1139[0],s1140[1],s1136[2]};
    assign in1365_2 = {s1116[3],s1140[0],s1141[1],s1137[2]};
    CLA_4 KS_1365(s1365, c1365, in1365_1, in1365_2);
    wire[3:0] s1366, in1366_1, in1366_2;
    wire c1366;
    assign in1366_1 = {s1117[3],s1141[0],s1142[1],s1138[2]};
    assign in1366_2 = {s1118[3],s1142[0],c1143,s1139[2]};
    CLA_4 KS_1366(s1366, c1366, in1366_1, in1366_2);
    wire[3:0] s1367, in1367_1, in1367_2;
    wire c1367;
    assign in1367_1 = {s1119[3],s1143[0],s1144[1],s1140[2]};
    assign in1367_2 = {s1120[3],s1144[0],c1145,s1141[2]};
    CLA_4 KS_1367(s1367, c1367, in1367_1, in1367_2);
    wire[3:0] s1368, in1368_1, in1368_2;
    wire c1368;
    assign in1368_1 = {s1121[3],s1145[0],s1146[1],s1142[2]};
    assign in1368_2 = {s1122[3],s1146[0],c1147,c1144};
    CLA_4 KS_1368(s1368, c1368, in1368_1, in1368_2);
    wire[1:0] s1369, in1369_1, in1369_2;
    wire c1369;
    assign in1369_1 = {s1123[3],s1147[0]};
    assign in1369_2 = {s1124[3],s1148[0]};
    CLA_2 KS_1369(s1369, c1369, in1369_1, in1369_2);
    wire[0:0] s1370, in1370_1, in1370_2;
    wire c1370;
    assign in1370_1 = {s1127[3]};
    assign in1370_2 = {c1131};
    Half_Adder KS_1370(s1370, c1370, in1370_1, in1370_2);
    wire[2:0] s1371, in1371_1, in1371_2;
    wire c1371;
    assign in1371_1 = {c1354,s1149[0],s1148[1]};
    assign in1371_2 = {c1355,s1150[0],c1149};
    CLA_3 KS_1371(s1371, c1371, in1371_1, in1371_2);
    wire[0:0] s1372, in1372_1, in1372_2;
    wire c1372;
    assign in1372_1 = {c1356};
    assign in1372_2 = {c1357};
    Half_Adder KS_1372(s1372, c1372, in1372_1, in1372_2);
    wire[1:0] s1373, in1373_1, in1373_2;
    wire c1373;
    assign in1373_1 = {c1363,s1364[1]};
    assign in1373_2 = {s1364[0],s1365[1]};
    CLA_2_c KS_1373(s1373, c1373, in1373_1, in1373_2, c1358);
    wire[3:0] s1374, in1374_1, in1374_2;
    wire c1374;
    assign in1374_1 = {c777,s1154[0],s1155[1],pp63[45]};
    assign in1374_2 = {s779[2],s1155[0],s1156[1],s1151[2]};
    CLA_4 KS_1374(s1374, c1374, in1374_1, in1374_2);
    wire[3:0] s1375, in1375_1, in1375_2;
    wire c1375;
    assign in1375_1 = {s1133[3],s1156[0],s1157[1],s1152[2]};
    assign in1375_2 = {s1134[3],s1157[0],c1158,s1153[2]};
    CLA_4 KS_1375(s1375, c1375, in1375_1, in1375_2);
    wire[3:0] s1376, in1376_1, in1376_2;
    wire c1376;
    assign in1376_1 = {s1135[3],s1158[0],s1159[1],s1154[2]};
    assign in1376_2 = {s1136[3],s1159[0],c1160,s1155[2]};
    CLA_4 KS_1376(s1376, c1376, in1376_1, in1376_2);
    wire[3:0] s1377, in1377_1, in1377_2;
    wire c1377;
    assign in1377_1 = {s1137[3],s1160[0],s1161[1],s1156[2]};
    assign in1377_2 = {s1138[3],s1161[0],c1162,c1157};
    CLA_4 KS_1377(s1377, c1377, in1377_1, in1377_2);
    wire[3:0] s1378, in1378_1, in1378_2;
    wire c1378;
    assign in1378_1 = {s1139[3],s1162[0],s1163[1],s1159[2]};
    assign in1378_2 = {s1140[3],s1163[0],c1164,c1161};
    CLA_4 KS_1378(s1378, c1378, in1378_1, in1378_2);
    wire[1:0] s1379, in1379_1, in1379_2;
    wire c1379;
    assign in1379_1 = {s1141[3],s1164[0]};
    assign in1379_2 = {c1142,s1165[0]};
    CLA_2 KS_1379(s1379, c1379, in1379_1, in1379_2);
    wire[0:0] s1380, in1380_1, in1380_2;
    wire c1380;
    assign in1380_1 = {s1146[3]};
    assign in1380_2 = {c1150};
    Half_Adder KS_1380(s1380, c1380, in1380_1, in1380_2);
    wire[2:0] s1381, in1381_1, in1381_2;
    wire c1381;
    assign in1381_1 = {c1364,s1166[0],s1165[1]};
    assign in1381_2 = {c1365,s1167[0],c1166};
    CLA_3 KS_1381(s1381, c1381, in1381_1, in1381_2);
    wire[0:0] s1382, in1382_1, in1382_2;
    wire c1382;
    assign in1382_1 = {c1367};
    assign in1382_2 = {c1368};
    Full_Adder KS_1382(s1382, c1382, in1382_1, in1382_2, c1366);
    wire[3:0] s1383, in1383_1, in1383_2;
    wire c1383;
    assign in1383_1 = {pp60[49],c1153,pp60[51],pp57[55]};
    assign in1383_2 = {pp61[48],c1154,pp61[50],pp58[54]};
    CLA_4 KS_1383(s1383, c1383, in1383_1, in1383_2);
    wire[3:0] s1384, in1384_1, in1384_2;
    wire c1384;
    assign in1384_1 = {pp62[47],c1155,pp62[49],pp59[53]};
    assign in1384_2 = {pp63[46],c1159,pp63[48],pp60[52]};
    CLA_4 KS_1384(s1384, c1384, in1384_1, in1384_2);
    wire[3:0] s1385, in1385_1, in1385_2;
    wire c1385;
    assign in1385_1 = {s1151[3],c1167,s1168[1],pp61[51]};
    assign in1385_2 = {s1152[3],s1168[0],s1169[1],pp62[50]};
    CLA_4 KS_1385(s1385, c1385, in1385_1, in1385_2);
    wire[3:0] s1386, in1386_1, in1386_2;
    wire c1386;
    assign in1386_1 = {s1153[3],s1169[0],s1170[1],pp63[49]};
    assign in1386_2 = {s1154[3],s1170[0],c1171,s1168[2]};
    CLA_4 KS_1386(s1386, c1386, in1386_1, in1386_2);
    wire[3:0] s1387, in1387_1, in1387_2;
    wire c1387;
    assign in1387_1 = {s1155[3],s1171[0],s1172[1],s1169[2]};
    assign in1387_2 = {c1156,s1172[0],c1173,c1170};
    CLA_4 KS_1387(s1387, c1387, in1387_1, in1387_2);
    wire[1:0] s1388, in1388_1, in1388_2;
    wire c1388;
    assign in1388_1 = {s1159[3],s1173[0]};
    assign in1388_2 = {c1163,s1174[0]};
    CLA_2 KS_1388(s1388, c1388, in1388_1, in1388_2);
    wire[0:0] s1389, in1389_1, in1389_2;
    wire c1389;
    assign in1389_1 = {s1167[3]};
    assign in1389_2 = {c1374};
    Half_Adder KS_1389(s1389, c1389, in1389_1, in1389_2);
    wire[2:0] s1390, in1390_1, in1390_2;
    wire c1390;
    assign in1390_1 = {c1376,s1175[0],s1174[1]};
    assign in1390_2 = {c1377,s1176[0],c1175};
    CLA_3_c KS_1390(s1390, c1390, in1390_1, in1390_2, c1375);
    wire[3:0] s1391, in1391_1, in1391_2;
    wire c1391;
    assign in1391_1 = {pp54[59],pp53[61],pp52[63],pp53[63]};
    assign in1391_2 = {pp55[58],pp54[60],pp53[62],pp54[62]};
    CLA_4 KS_1391(s1391, c1391, in1391_1, in1391_2);
    wire[3:0] s1392, in1392_1, in1392_2;
    wire c1392;
    assign in1392_1 = {pp56[57],pp55[59],pp54[61],pp55[61]};
    assign in1392_2 = {pp57[56],pp56[58],pp55[60],pp56[60]};
    CLA_4 KS_1392(s1392, c1392, in1392_1, in1392_2);
    wire[3:0] s1393, in1393_1, in1393_2;
    wire c1393;
    assign in1393_1 = {pp58[55],pp57[57],pp56[59],pp57[59]};
    assign in1393_2 = {pp59[54],pp58[56],pp57[58],pp58[58]};
    CLA_4 KS_1393(s1393, c1393, in1393_1, in1393_2);
    wire[2:0] s1394, in1394_1, in1394_2;
    wire c1394;
    assign in1394_1 = {pp60[53],pp59[55],pp58[57]};
    assign in1394_2 = {pp61[52],pp60[54],pp59[56]};
    CLA_3 KS_1394(s1394, c1394, in1394_1, in1394_2);
    wire[3:0] s1395, in1395_1, in1395_2;
    wire c1395;
    assign in1395_1 = {pp62[51],pp61[53],pp60[55],pp59[57]};
    assign in1395_2 = {pp63[50],pp62[52],pp61[54],pp60[56]};
    CLA_4 KS_1395(s1395, c1395, in1395_1, in1395_2);
    wire[1:0] s1396, in1396_1, in1396_2;
    wire c1396;
    assign in1396_1 = {s1168[3],pp63[51]};
    assign in1396_2 = {c1169,c1168};
    CLA_2 KS_1396(s1396, c1396, in1396_1, in1396_2);
    wire[0:0] s1397, in1397_1, in1397_2;
    wire c1397;
    assign in1397_1 = {s1172[3]};
    assign in1397_2 = {c1176};
    Half_Adder KS_1397(s1397, c1397, in1397_1, in1397_2);
    wire[2:0] s1398, in1398_1, in1398_2;
    wire c1398;
    assign in1398_1 = {c1383,c1172,pp62[53]};
    assign in1398_2 = {c1384,s1177[0],pp63[52]};
    CLA_3 KS_1398(s1398, c1398, in1398_1, in1398_2);
    wire[0:0] s1399, in1399_1, in1399_2;
    wire c1399;
    assign in1399_1 = {c1386};
    assign in1399_2 = {c1387};
    Full_Adder KS_1399(s1399, c1399, in1399_1, in1399_2, c1385);
    wire[1:0] s1400, in1400_1, in1400_2;
    wire c1400;
    assign in1400_1 = {pp54[63],pp55[63]};
    assign in1400_2 = {pp55[62],pp56[62]};
    CLA_2 KS_1400(s1400, c1400, in1400_1, in1400_2);
    wire[0:0] s1401, in1401_1, in1401_2;
    wire c1401;
    assign in1401_1 = {pp56[61]};
    assign in1401_2 = {pp57[60]};
    Half_Adder KS_1401(s1401, c1401, in1401_1, in1401_2);
    wire[2:0] s1402, in1402_1, in1402_2;
    wire c1402;
    assign in1402_1 = {pp58[59],pp57[61],pp56[63]};
    assign in1402_2 = {pp59[58],pp58[60],pp57[62]};
    CLA_3 KS_1402(s1402, c1402, in1402_1, in1402_2);
    wire[0:0] s1403, in1403_1, in1403_2;
    wire c1403;
    assign in1403_1 = {pp61[56]};
    assign in1403_2 = {pp62[55]};
    Full_Adder KS_1403(s1403, c1403, in1403_1, in1403_2, pp60[57]);

    /*Stage 5*/
    wire[3:0] s1404, in1404_1, in1404_2;
    wire c1404;
    assign in1404_1 = {pp0[6],pp0[7],pp0[8],pp2[7]};
    assign in1404_2 = {pp1[5],pp1[6],pp1[7],pp3[6]};
    CLA_4 KS_1404(s1404, c1404, in1404_1, in1404_2);
    wire[3:0] s1405, in1405_1, in1405_2;
    wire c1405;
    assign in1405_1 = {pp2[5],pp2[6],pp4[5],pp4[6]};
    assign in1405_2 = {pp3[4],pp3[5],pp5[4],pp5[5]};
    CLA_4 KS_1405(s1405, c1405, in1405_1, in1405_2);
    wire[3:0] s1406, in1406_1, in1406_2;
    wire c1406;
    assign in1406_1 = {pp4[4],pp6[3],pp6[4],pp6[5]};
    assign in1406_2 = {pp5[3],pp7[2],pp7[3],pp7[4]};
    CLA_4 KS_1406(s1406, c1406, in1406_1, in1406_2);
    wire[3:0] s1407, in1407_1, in1407_2;
    wire c1407;
    assign in1407_1 = {pp9[1],pp8[3],pp8[4],pp11[2]};
    assign in1407_2 = {pp10[0],pp9[2],pp9[3],pp12[1]};
    CLA_4_c KS_1407(s1407, c1407, in1407_1, in1407_2, pp8[2]);
    wire[3:0] s1408, in1408_1, in1408_2;
    wire c1408;
    assign in1408_1 = {pp11[0],pp10[2],pp13[0],pp13[1]};
    assign in1408_2 = {s1178[2],pp11[1],c1178,pp14[0]};
    CLA_4_c KS_1408(s1408, c1408, in1408_1, in1408_2, pp10[1]);
    wire[3:0] s1409, in1409_1, in1409_2;
    wire c1409;
    assign in1409_1 = {s1178[3],s1179[3],s781[0],pp15[0]};
    assign in1409_2 = {s1179[2],s1180[2],c1179,s781[1]};
    CLA_4_c KS_1409(s1409, c1409, in1409_1, in1409_2, pp12[0]);
    wire[3:0] s1410, in1410_1, in1410_2;
    wire c1410;
    assign in1410_1 = {s1181[2],s782[0],s781[2],s784[0]};
    assign in1410_2 = {s1182[1],c1180,s782[1],c1182};
    CLA_4_c KS_1410(s1410, c1410, in1410_1, in1410_2, s1180[3]);
    wire[3:0] s1411, in1411_1, in1411_2;
    wire c1411;
    assign in1411_1 = {s1182[2],s783[0],c1183,s785[0]};
    assign in1411_2 = {s1183[2],c1181,s1184[3],s786[0]};
    CLA_4_c KS_1411(s1411, c1411, in1411_1, in1411_2, s1181[3]);
    wire[3:0] s1412, in1412_1, in1412_2;
    wire c1412;
    assign in1412_1 = {s1183[3],s1185[2],c1184,s787[0]};
    assign in1412_2 = {s1184[2],s1186[1],s1185[3],s788[0]};
    CLA_4_c KS_1412(s1412, c1412, in1412_1, in1412_2, s1182[3]);
    wire[3:0] s1413, in1413_1, in1413_2;
    wire c1413;
    assign in1413_1 = {s1187[1],c1185,s789[0],c1188};
    assign in1413_2 = {s1188[1],s1186[3],s790[0],c1189};
    CLA_4_c KS_1413(s1413, c1413, in1413_1, in1413_2, s1186[2]);
    wire[3:0] s1414, in1414_1, in1414_2;
    wire c1414;
    assign in1414_1 = {s1188[2],c1186,s1190[3],s795[0]};
    assign in1414_2 = {s1189[2],s1187[3],s1191[2],s796[0]};
    CLA_4_c KS_1414(s1414, c1414, in1414_1, in1414_2, s1187[2]);
    wire[3:0] s1415, in1415_1, in1415_2;
    wire c1415;
    assign in1415_1 = {s1189[3],s1192[1],c1190,s797[0]};
    assign in1415_2 = {s1190[2],s1193[0],s1191[3],s798[0]};
    CLA_4_c KS_1415(s1415, c1415, in1415_1, in1415_2, s1188[3]);
    wire[3:0] s1416, in1416_1, in1416_2;
    wire c1416;
    assign in1416_1 = {s1193[1],c1191,s799[0],c1196};
    assign in1416_2 = {s1194[1],s1192[3],s800[0],s1197[2]};
    CLA_4_c KS_1416(s1416, c1416, in1416_1, in1416_2, s1192[2]);
    wire[3:0] s1417, in1417_1, in1417_2;
    wire c1417;
    assign in1417_1 = {s1194[2],c1192,s1198[1],s1197[3]};
    assign in1417_2 = {s1195[2],s1193[3],s1199[0],s1198[2]};
    CLA_4_c KS_1417(s1417, c1417, in1417_1, in1417_2, s1193[2]);
    wire[3:0] s1418, in1418_1, in1418_2;
    wire c1418;
    assign in1418_1 = {s1195[3],s1200[0],s1199[1],s808[1]};
    assign in1418_2 = {s1196[3],s1201[0],s1200[1],s809[0]};
    CLA_4_c KS_1418(s1418, c1418, in1418_1, in1418_2, s1194[3]);
    wire[3:0] s1419, in1419_1, in1419_2;
    wire c1419;
    assign in1419_1 = {s1201[1],c1197,s809[1],s1205[1]};
    assign in1419_2 = {s1202[1],s1198[3],s810[0],s1206[0]};
    CLA_4 KS_1419(s1419, c1419, in1419_1, in1419_2);
    wire[3:0] s1420, in1420_1, in1420_2;
    wire c1420;
    assign in1420_1 = {s1200[2],c1198,s1207[0],s1205[2]};
    assign in1420_2 = {s1201[2],s1199[3],s1208[0],s1206[1]};
    CLA_4_c KS_1420(s1420, c1420, in1420_1, in1420_2, s1199[2]);
    wire[3:0] s1421, in1421_1, in1421_2;
    wire c1421;
    assign in1421_1 = {s1201[3],s1209[0],s1207[1],s822[1]};
    assign in1421_2 = {s1202[3],s1210[0],s1208[1],s1205[3]};
    CLA_4_c KS_1421(s1421, c1421, in1421_1, in1421_2, s1200[3]);
    wire[3:0] s1422, in1422_1, in1422_2;
    wire c1422;
    assign in1422_1 = {s1210[1],s1206[2],s819[2],s1214[0]};
    assign in1422_2 = {c1211,s1207[2],s820[2],s1215[0]};
    CLA_4_c KS_1422(s1422, c1422, in1422_1, in1422_2, s1209[1]);
    wire[3:0] s1423, in1423_1, in1423_2;
    wire c1423;
    assign in1423_1 = {s1208[2],s822[2],s1216[0],s1214[1]};
    assign in1423_2 = {s1209[2],c1205,s1217[0],s1215[1]};
    CLA_4 KS_1423(s1423, c1423, in1423_1, in1423_2);
    wire[3:0] s1424, in1424_1, in1424_2;
    wire c1424;
    assign in1424_1 = {s1207[3],s1218[0],s1216[1],s838[1]};
    assign in1424_2 = {s1208[3],s1219[0],s1217[1],c839};
    CLA_4_c KS_1424(s1424, c1424, in1424_1, in1424_2, s1206[3]);
    wire[3:0] s1425, in1425_1, in1425_2;
    wire c1425;
    assign in1425_1 = {s1219[1],s1214[2],s836[2],s1224[0]};
    assign in1425_2 = {c1220,s1215[2],c838,s1225[0]};
    CLA_4_c KS_1425(s1425, c1425, in1425_1, in1425_2, s1218[1]);
    wire[3:0] s1426, in1426_1, in1426_2;
    wire c1426;
    assign in1426_1 = {s1217[2],s1214[3],s1226[0],s1225[1]};
    assign in1426_2 = {s1218[2],s1215[3],s1227[0],s1226[1]};
    CLA_4_c KS_1426(s1426, c1426, in1426_1, in1426_2, s1216[2]);
    wire[3:0] s1427, in1427_1, in1427_2;
    wire c1427;
    assign in1427_1 = {s1216[3],s1228[0],s1227[1],s857[1]};
    assign in1427_2 = {s1217[3],s1229[0],s1228[1],s1223[2]};
    CLA_4 KS_1427(s1427, c1427, in1427_1, in1427_2);
    wire[3:0] s1428, in1428_1, in1428_2;
    wire c1428;
    assign in1428_1 = {c1229,s1224[2],s853[2],c1227};
    assign in1428_2 = {s1230[1],s1225[2],c855,s1233[0]};
    CLA_4 KS_1428(s1428, c1428, in1428_1, in1428_2);
    wire[3:0] s1429, in1429_1, in1429_2;
    wire c1429;
    assign in1429_1 = {s1227[2],s857[2],s1234[0],s1233[1]};
    assign in1429_2 = {c1228,s1223[3],s1235[0],s1234[1]};
    CLA_4_c KS_1429(s1429, c1429, in1429_1, in1429_2, s1226[2]);
    wire[3:0] s1430, in1430_1, in1430_2;
    wire c1430;
    assign in1430_1 = {s1225[3],s1236[0],s1235[1],s875[1]};
    assign in1430_2 = {s1226[3],s1237[0],s1236[1],c876};
    CLA_4_c KS_1430(s1430, c1430, in1430_1, in1430_2, s1224[3]);
    wire[3:0] s1431, in1431_1, in1431_2;
    wire c1431;
    assign in1431_1 = {s1237[1],s1233[2],s871[2],c1237};
    assign in1431_2 = {s1238[1],s1234[2],c873,s1241[0]};
    CLA_4 KS_1431(s1431, c1431, in1431_1, in1431_2);
    wire[3:0] s1432, in1432_1, in1432_2;
    wire c1432;
    assign in1432_1 = {s1236[2],s875[2],s1242[0],s1241[1]};
    assign in1432_2 = {s1237[2],s1233[3],s1243[0],s1242[1]};
    CLA_4_c KS_1432(s1432, c1432, in1432_1, in1432_2, s1235[2]);
    wire[3:0] s1433, in1433_1, in1433_2;
    wire c1433;
    assign in1433_1 = {s1235[3],s1244[0],s1243[1],s894[1]};
    assign in1433_2 = {s1236[3],s1245[0],s1244[1],c895};
    CLA_4_c KS_1433(s1433, c1433, in1433_1, in1433_2, s1234[3]);
    wire[3:0] s1434, in1434_1, in1434_2;
    wire c1434;
    assign in1434_1 = {s1245[1],s1241[2],s892[2],s1249[0]};
    assign in1434_2 = {s1246[1],s1242[2],c894,s1250[0]};
    CLA_4 KS_1434(s1434, c1434, in1434_1, in1434_2);
    wire[3:0] s1435, in1435_1, in1435_2;
    wire c1435;
    assign in1435_1 = {s1244[2],s1241[3],s1251[0],s1249[1]};
    assign in1435_2 = {s1245[2],s1242[3],s1252[0],s1250[1]};
    CLA_4_c KS_1435(s1435, c1435, in1435_1, in1435_2, s1243[2]);
    wire[3:0] s1436, in1436_1, in1436_2;
    wire c1436;
    assign in1436_1 = {s1243[3],s1253[0],s1251[1],s913[1]};
    assign in1436_2 = {s1244[3],s1254[0],s1252[1],s1249[2]};
    CLA_4 KS_1436(s1436, c1436, in1436_1, in1436_2);
    wire[3:0] s1437, in1437_1, in1437_2;
    wire c1437;
    assign in1437_1 = {s1254[1],s1250[2],s909[2],c1253};
    assign in1437_2 = {c1255,s1251[2],c911,s1258[0]};
    CLA_4_c KS_1437(s1437, c1437, in1437_1, in1437_2, s1253[1]);
    wire[3:0] s1438, in1438_1, in1438_2;
    wire c1438;
    assign in1438_1 = {s1252[2],s913[2],s1259[0],s1258[1]};
    assign in1438_2 = {s1253[2],s1249[3],s1260[0],s1259[1]};
    CLA_4 KS_1438(s1438, c1438, in1438_1, in1438_2);
    wire[3:0] s1439, in1439_1, in1439_2;
    wire c1439;
    assign in1439_1 = {s1251[3],s1261[0],s1260[1],s931[1]};
    assign in1439_2 = {s1252[3],s1262[0],s1261[1],c932};
    CLA_4_c KS_1439(s1439, c1439, in1439_1, in1439_2, s1250[3]);
    wire[3:0] s1440, in1440_1, in1440_2;
    wire c1440;
    assign in1440_1 = {s1262[1],s1258[2],s927[2],c1262};
    assign in1440_2 = {s1263[1],s1259[2],c929,s1266[0]};
    CLA_4 KS_1440(s1440, c1440, in1440_1, in1440_2);
    wire[3:0] s1441, in1441_1, in1441_2;
    wire c1441;
    assign in1441_1 = {s1261[2],s931[2],s1267[0],s1266[1]};
    assign in1441_2 = {s1262[2],s1258[3],s1268[0],s1267[1]};
    CLA_4_c KS_1441(s1441, c1441, in1441_1, in1441_2, s1260[2]);
    wire[3:0] s1442, in1442_1, in1442_2;
    wire c1442;
    assign in1442_1 = {s1260[3],s1269[0],s1268[1],s950[1]};
    assign in1442_2 = {s1261[3],s1270[0],s1269[1],c951};
    CLA_4_c KS_1442(s1442, c1442, in1442_1, in1442_2, s1259[3]);
    wire[3:0] s1443, in1443_1, in1443_2;
    wire c1443;
    assign in1443_1 = {s1270[1],s1266[2],s946[2],c1270};
    assign in1443_2 = {s1271[1],s1267[2],c948,s1274[0]};
    CLA_4 KS_1443(s1443, c1443, in1443_1, in1443_2);
    wire[3:0] s1444, in1444_1, in1444_2;
    wire c1444;
    assign in1444_1 = {s1269[2],s950[2],s1275[0],s1274[1]};
    assign in1444_2 = {s1270[2],s1266[3],s1276[0],s1275[1]};
    CLA_4_c KS_1444(s1444, c1444, in1444_1, in1444_2, s1268[2]);
    wire[3:0] s1445, in1445_1, in1445_2;
    wire c1445;
    assign in1445_1 = {s1268[3],s1277[0],s1276[1],s969[1]};
    assign in1445_2 = {s1269[3],s1278[0],s1277[1],c970};
    CLA_4_c KS_1445(s1445, c1445, in1445_1, in1445_2, s1267[3]);
    wire[3:0] s1446, in1446_1, in1446_2;
    wire c1446;
    assign in1446_1 = {s1278[1],s1274[2],s967[2],s1283[0]};
    assign in1446_2 = {s1279[1],s1275[2],c969,s1284[0]};
    CLA_4 KS_1446(s1446, c1446, in1446_1, in1446_2);
    wire[3:0] s1447, in1447_1, in1447_2;
    wire c1447;
    assign in1447_1 = {s1277[2],s1274[3],s1285[0],s1284[1]};
    assign in1447_2 = {s1278[2],s1275[3],s1286[0],s1285[1]};
    CLA_4_c KS_1447(s1447, c1447, in1447_1, in1447_2, s1276[2]);
    wire[3:0] s1448, in1448_1, in1448_2;
    wire c1448;
    assign in1448_1 = {s1276[3],s1287[0],s1286[1],s988[1]};
    assign in1448_2 = {s1277[3],s1288[0],s1287[1],s1282[2]};
    CLA_4 KS_1448(s1448, c1448, in1448_1, in1448_2);
    wire[3:0] s1449, in1449_1, in1449_2;
    wire c1449;
    assign in1449_1 = {c1288,s1283[2],s984[2],s1292[0]};
    assign in1449_2 = {s1289[1],s1284[2],c986,s1293[0]};
    CLA_4 KS_1449(s1449, c1449, in1449_1, in1449_2);
    wire[3:0] s1450, in1450_1, in1450_2;
    wire c1450;
    assign in1450_1 = {s1286[2],s988[2],s1294[0],s1292[1]};
    assign in1450_2 = {c1287,s1282[3],s1295[0],s1293[1]};
    CLA_4_c KS_1450(s1450, c1450, in1450_1, in1450_2, s1285[2]);
    wire[3:0] s1451, in1451_1, in1451_2;
    wire c1451;
    assign in1451_1 = {s1284[3],s1296[0],s1294[1],s1006[1]};
    assign in1451_2 = {s1285[3],s1297[0],s1295[1],s1292[2]};
    CLA_4_c KS_1451(s1451, c1451, in1451_1, in1451_2, s1283[3]);
    wire[3:0] s1452, in1452_1, in1452_2;
    wire c1452;
    assign in1452_1 = {s1297[1],s1293[2],s1002[2],s1301[0]};
    assign in1452_2 = {c1298,s1294[2],c1004,s1302[0]};
    CLA_4_c KS_1452(s1452, c1452, in1452_1, in1452_2, s1296[1]);
    wire[3:0] s1453, in1453_1, in1453_2;
    wire c1453;
    assign in1453_1 = {s1295[2],s1006[2],s1303[0],s1301[1]};
    assign in1453_2 = {s1296[2],s1292[3],s1304[0],s1302[1]};
    CLA_4 KS_1453(s1453, c1453, in1453_1, in1453_2);
    wire[3:0] s1454, in1454_1, in1454_2;
    wire c1454;
    assign in1454_1 = {s1294[3],s1305[0],s1303[1],s1024[1]};
    assign in1454_2 = {s1295[3],s1306[0],s1304[1],s1301[2]};
    CLA_4_c KS_1454(s1454, c1454, in1454_1, in1454_2, s1293[3]);
    wire[3:0] s1455, in1455_1, in1455_2;
    wire c1455;
    assign in1455_1 = {s1306[1],s1302[2],s1022[2],s1310[0]};
    assign in1455_2 = {c1307,s1303[2],c1024,s1311[0]};
    CLA_4_c KS_1455(s1455, c1455, in1455_1, in1455_2, s1305[1]);
    wire[3:0] s1456, in1456_1, in1456_2;
    wire c1456;
    assign in1456_1 = {s1304[2],s1301[3],s1312[0],s1310[1]};
    assign in1456_2 = {s1305[2],s1302[3],s1313[0],s1311[1]};
    CLA_4 KS_1456(s1456, c1456, in1456_1, in1456_2);
    wire[3:0] s1457, in1457_1, in1457_2;
    wire c1457;
    assign in1457_1 = {s1303[3],s1314[0],s1312[1],s1042[1]};
    assign in1457_2 = {s1304[3],s1315[0],s1313[1],s1310[2]};
    CLA_4 KS_1457(s1457, c1457, in1457_1, in1457_2);
    wire[3:0] s1458, in1458_1, in1458_2;
    wire c1458;
    assign in1458_1 = {s1315[1],s1311[2],s1040[2],s1320[0]};
    assign in1458_2 = {c1316,s1312[2],c1042,s1321[0]};
    CLA_4_c KS_1458(s1458, c1458, in1458_1, in1458_2, s1314[1]);
    wire[3:0] s1459, in1459_1, in1459_2;
    wire c1459;
    assign in1459_1 = {s1313[2],s1310[3],s1322[0],s1321[1]};
    assign in1459_2 = {s1314[2],s1311[3],s1323[0],s1322[1]};
    CLA_4 KS_1459(s1459, c1459, in1459_1, in1459_2);
    wire[3:0] s1460, in1460_1, in1460_2;
    wire c1460;
    assign in1460_1 = {s1312[3],s1324[0],s1323[1],s1060[1]};
    assign in1460_2 = {s1313[3],s1325[0],s1324[1],s1319[2]};
    CLA_4 KS_1460(s1460, c1460, in1460_1, in1460_2);
    wire[3:0] s1461, in1461_1, in1461_2;
    wire c1461;
    assign in1461_1 = {c1325,s1320[2],s1056[2],c1323};
    assign in1461_2 = {s1326[1],s1321[2],c1058,s1329[0]};
    CLA_4 KS_1461(s1461, c1461, in1461_1, in1461_2);
    wire[3:0] s1462, in1462_1, in1462_2;
    wire c1462;
    assign in1462_1 = {s1323[2],s1060[2],s1330[0],s1329[1]};
    assign in1462_2 = {c1324,s1319[3],s1331[0],s1330[1]};
    CLA_4_c KS_1462(s1462, c1462, in1462_1, in1462_2, s1322[2]);
    wire[3:0] s1463, in1463_1, in1463_2;
    wire c1463;
    assign in1463_1 = {s1321[3],s1332[0],s1331[1],s1078[1]};
    assign in1463_2 = {s1322[3],s1333[0],s1332[1],s1329[2]};
    CLA_4_c KS_1463(s1463, c1463, in1463_1, in1463_2, s1320[3]);
    wire[3:0] s1464, in1464_1, in1464_2;
    wire c1464;
    assign in1464_1 = {s1333[1],s1330[2],s1074[2],s1337[0]};
    assign in1464_2 = {s1334[1],s1331[2],c1076,s1338[0]};
    CLA_4 KS_1464(s1464, c1464, in1464_1, in1464_2);
    wire[3:0] s1465, in1465_1, in1465_2;
    wire c1465;
    assign in1465_1 = {s1332[2],s1078[2],s1339[0],s1337[1]};
    assign in1465_2 = {s1333[2],s1329[3],s1340[0],s1338[1]};
    CLA_4 KS_1465(s1465, c1465, in1465_1, in1465_2);
    wire[3:0] s1466, in1466_1, in1466_2;
    wire c1466;
    assign in1466_1 = {s1331[3],s1341[0],s1339[1],s1096[1]};
    assign in1466_2 = {s1332[3],s1342[0],s1340[1],s1337[2]};
    CLA_4_c KS_1466(s1466, c1466, in1466_1, in1466_2, s1330[3]);
    wire[3:0] s1467, in1467_1, in1467_2;
    wire c1467;
    assign in1467_1 = {s1342[1],s1338[2],s1092[2],c1341};
    assign in1467_2 = {c1343,s1339[2],c1094,s1346[0]};
    CLA_4_c KS_1467(s1467, c1467, in1467_1, in1467_2, s1341[1]);
    wire[3:0] s1468, in1468_1, in1468_2;
    wire c1468;
    assign in1468_1 = {s1340[2],s1096[2],s1347[0],s1346[1]};
    assign in1468_2 = {s1341[2],s1337[3],s1348[0],s1347[1]};
    CLA_4 KS_1468(s1468, c1468, in1468_1, in1468_2);
    wire[3:0] s1469, in1469_1, in1469_2;
    wire c1469;
    assign in1469_1 = {s1339[3],s1349[0],s1348[1],s1114[1]};
    assign in1469_2 = {s1340[3],s1350[0],s1349[1],c1115};
    CLA_4_c KS_1469(s1469, c1469, in1469_1, in1469_2, s1338[3]);
    wire[3:0] s1470, in1470_1, in1470_2;
    wire c1470;
    assign in1470_1 = {s1350[1],s1346[2],s1112[2],s1355[0]};
    assign in1470_2 = {s1351[1],s1347[2],c1114,s1356[0]};
    CLA_4 KS_1470(s1470, c1470, in1470_1, in1470_2);
    wire[3:0] s1471, in1471_1, in1471_2;
    wire c1471;
    assign in1471_1 = {s1349[2],s1346[3],s1357[0],s1356[1]};
    assign in1471_2 = {s1350[2],s1347[3],s1358[0],s1357[1]};
    CLA_4_c KS_1471(s1471, c1471, in1471_1, in1471_2, s1348[2]);
    wire[3:0] s1472, in1472_1, in1472_2;
    wire c1472;
    assign in1472_1 = {s1348[3],s1359[0],s1358[1],s1354[2]};
    assign in1472_2 = {s1349[3],s1360[0],s1359[1],s1355[2]};
    CLA_4 KS_1472(s1472, c1472, in1472_1, in1472_2);
    wire[3:0] s1473, in1473_1, in1473_2;
    wire c1473;
    assign in1473_1 = {c1360,s1356[2],s1131[2],s1365[0]};
    assign in1473_2 = {s1361[1],s1357[2],s1354[3],s1366[0]};
    CLA_4 KS_1473(s1473, c1473, in1473_1, in1473_2);
    wire[3:0] s1474, in1474_1, in1474_2;
    wire c1474;
    assign in1474_1 = {s1358[2],s1355[3],s1367[0],s1366[1]};
    assign in1474_2 = {s1359[2],s1356[3],s1368[0],s1367[1]};
    CLA_4 KS_1474(s1474, c1474, in1474_1, in1474_2);
    wire[3:0] s1475, in1475_1, in1475_2;
    wire c1475;
    assign in1475_1 = {s1357[3],s1369[0],s1368[1],s1150[1]};
    assign in1475_2 = {s1358[3],s1370[0],s1369[1],s1364[2]};
    CLA_4 KS_1475(s1475, c1475, in1475_1, in1475_2);
    wire[3:0] s1476, in1476_1, in1476_2;
    wire c1476;
    assign in1476_1 = {c1370,s1365[2],s1146[2],s1374[0]};
    assign in1476_2 = {s1371[1],s1366[2],c1148,s1375[0]};
    CLA_4 KS_1476(s1476, c1476, in1476_1, in1476_2);
    wire[3:0] s1477, in1477_1, in1477_2;
    wire c1477;
    assign in1477_1 = {s1368[2],s1150[2],s1376[0],s1374[1]};
    assign in1477_2 = {c1369,s1364[3],s1377[0],s1375[1]};
    CLA_4_c KS_1477(s1477, c1477, in1477_1, in1477_2, s1367[2]);
    wire[3:0] s1478, in1478_1, in1478_2;
    wire c1478;
    assign in1478_1 = {s1366[3],s1378[0],s1376[1],s1167[1]};
    assign in1478_2 = {s1367[3],s1379[0],s1377[1],s1374[2]};
    CLA_4_c KS_1478(s1478, c1478, in1478_1, in1478_2, s1365[3]);
    wire[3:0] s1479, in1479_1, in1479_2;
    wire c1479;
    assign in1479_1 = {s1379[1],s1375[2],s1163[2],c1378};
    assign in1479_2 = {c1380,s1376[2],c1165,s1383[0]};
    CLA_4_c KS_1479(s1479, c1479, in1479_1, in1479_2, s1378[1]);
    wire[3:0] s1480, in1480_1, in1480_2;
    wire c1480;
    assign in1480_1 = {s1377[2],s1167[2],s1384[0],s1383[1]};
    assign in1480_2 = {s1378[2],s1374[3],s1385[0],s1384[1]};
    CLA_4 KS_1480(s1480, c1480, in1480_1, in1480_2);
    wire[3:0] s1481, in1481_1, in1481_2;
    wire c1481;
    assign in1481_1 = {s1376[3],s1386[0],s1385[1],s1176[1]};
    assign in1481_2 = {s1377[3],s1387[0],s1386[1],s1383[2]};
    CLA_4_c KS_1481(s1481, c1481, in1481_1, in1481_2, s1375[3]);
    wire[3:0] s1482, in1482_1, in1482_2;
    wire c1482;
    assign in1482_1 = {s1387[1],s1384[2],s1172[2],s1391[0]};
    assign in1482_2 = {s1388[1],s1385[2],c1174,s1392[0]};
    CLA_4 KS_1482(s1482, c1482, in1482_1, in1482_2);
    wire[3:0] s1483, in1483_1, in1483_2;
    wire c1483;
    assign in1483_1 = {s1386[2],s1176[2],s1393[0],s1391[1]};
    assign in1483_2 = {s1387[2],s1383[3],s1394[0],s1392[1]};
    CLA_4 KS_1483(s1483, c1483, in1483_1, in1483_2);
    wire[3:0] s1484, in1484_1, in1484_2;
    wire c1484;
    assign in1484_1 = {s1385[3],s1395[0],s1393[1],c1177};
    assign in1484_2 = {s1386[3],s1396[0],s1394[1],s1391[2]};
    CLA_4_c KS_1484(s1484, c1484, in1484_1, in1484_2, s1384[3]);
    wire[3:0] s1485, in1485_1, in1485_2;
    wire c1485;
    assign in1485_1 = {s1396[1],s1392[2],pp61[55],pp63[54]};
    assign in1485_2 = {c1397,s1393[2],pp62[54],c1391};
    CLA_4_c KS_1485(s1485, c1485, in1485_1, in1485_2, s1395[1]);
    wire[3:0] s1486, in1486_1, in1486_2;
    wire c1486;
    assign in1486_1 = {s1394[2],pp63[53],c1392,pp59[59]};
    assign in1486_2 = {s1395[2],s1391[3],c1393,pp60[58]};
    CLA_4 KS_1486(s1486, c1486, in1486_1, in1486_2);
    wire[3:0] s1487, in1487_1, in1487_2;
    wire c1487;
    assign in1487_1 = {s1393[3],c1395,pp61[57],pp58[61]};
    assign in1487_2 = {c1394,s1400[0],pp62[56],pp59[60]};
    CLA_4_c KS_1487(s1487, c1487, in1487_1, in1487_2, s1392[3]);
    wire[3:0] s1488, in1488_1, in1488_2;
    wire c1488;
    assign in1488_1 = {s1400[1],pp60[59],pp57[63],pp58[63]};
    assign in1488_2 = {c1401,pp61[58],pp58[62],pp59[62]};
    CLA_4_c KS_1488(s1488, c1488, in1488_1, in1488_2, pp63[55]);
    wire[1:0] s1489, in1489_1, in1489_2;
    wire c1489;
    assign in1489_1 = {pp62[57],pp59[61]};
    assign in1489_2 = {pp63[56],pp60[60]};
    CLA_2 KS_1489(s1489, c1489, in1489_1, in1489_2);
    wire[2:0] s1490, in1490_1, in1490_2;
    wire c1490;
    assign in1490_1 = {pp61[59],pp60[61],pp59[63]};
    assign in1490_2 = {pp62[58],pp61[60],pp60[62]};
    CLA_3 KS_1490(s1490, c1490, in1490_1, in1490_2);

    /*Stage 6*/
    wire[3:0] s1491, in1491_1, in1491_2;
    wire c1491;
    assign in1491_1 = {pp0[4],pp0[5],pp2[4],pp4[3]};
    assign in1491_2 = {pp1[3],pp1[4],pp3[3],pp5[2]};
    CLA_4 KS_1491(s1491, c1491, in1491_1, in1491_2);
    wire[3:0] s1492, in1492_1, in1492_2;
    wire c1492;
    assign in1492_1 = {pp2[3],pp4[2],pp6[1],pp6[2]};
    assign in1492_2 = {pp3[2],pp5[1],pp7[0],pp7[1]};
    CLA_4 KS_1492(s1492, c1492, in1492_1, in1492_2);
    wire[3:0] s1493, in1493_1, in1493_2;
    wire c1493;
    assign in1493_1 = {s1404[2],pp8[1],s1178[1],s1179[1]};
    assign in1493_2 = {s1405[1],pp9[0],s1179[0],s1180[0]};
    CLA_4_c KS_1493(s1493, c1493, in1493_1, in1493_2, pp8[0]);
    wire[3:0] s1494, in1494_1, in1494_2;
    wire c1494;
    assign in1494_1 = {s1404[3],c1404,c1405,s1180[1]};
    assign in1494_2 = {s1405[2],s1405[3],s1406[3],s1181[0]};
    CLA_4_c KS_1494(s1494, c1494, in1494_1, in1494_2, s1178[0]);
    wire[3:0] s1495, in1495_1, in1495_2;
    wire c1495;
    assign in1495_1 = {s1407[2],s1181[1],s1183[1],s1184[1]};
    assign in1495_2 = {s1408[1],s1182[0],s1184[0],s1185[0]};
    CLA_4_c KS_1495(s1495, c1495, in1495_1, in1495_2, c1406);
    wire[3:0] s1496, in1496_1, in1496_2;
    wire c1496;
    assign in1496_1 = {s1407[3],c1407,c1408,s1185[1]};
    assign in1496_2 = {s1408[2],s1408[3],s1409[3],s1186[0]};
    CLA_4_c KS_1496(s1496, c1496, in1496_1, in1496_2, s1183[0]);
    wire[3:0] s1497, in1497_1, in1497_2;
    wire c1497;
    assign in1497_1 = {s1410[2],s1187[0],s1189[1],s1190[1]};
    assign in1497_2 = {s1411[1],s1188[0],s1190[0],s1191[0]};
    CLA_4_c KS_1497(s1497, c1497, in1497_1, in1497_2, c1409);
    wire[3:0] s1498, in1498_1, in1498_2;
    wire c1498;
    assign in1498_1 = {s1410[3],c1410,c1411,s1191[1]};
    assign in1498_2 = {s1411[2],s1411[3],s1412[3],s1192[0]};
    CLA_4_c KS_1498(s1498, c1498, in1498_1, in1498_2, s1189[0]);
    wire[3:0] s1499, in1499_1, in1499_2;
    wire c1499;
    assign in1499_1 = {s1413[2],s1194[0],s1195[1],s1196[2]};
    assign in1499_2 = {s1414[1],s1195[0],s1196[1],s1197[0]};
    CLA_4_c KS_1499(s1499, c1499, in1499_1, in1499_2, c1412);
    wire[3:0] s1500, in1500_1, in1500_2;
    wire c1500;
    assign in1500_1 = {s1413[3],c1413,c1414,s1197[1]};
    assign in1500_2 = {s1414[2],s1414[3],s1415[3],s1198[0]};
    CLA_4_c KS_1500(s1500, c1500, in1500_1, in1500_2, s1196[0]);
    wire[3:0] s1501, in1501_1, in1501_2;
    wire c1501;
    assign in1501_1 = {s1416[2],s1202[0],c1203,s1202[2]};
    assign in1501_2 = {s1417[1],s1203[0],s1204[1],s1204[2]};
    CLA_4_c KS_1501(s1501, c1501, in1501_1, in1501_2, c1415);
    wire[3:0] s1502, in1502_1, in1502_2;
    wire c1502;
    assign in1502_1 = {s1416[3],c1416,c1417,s1204[3]};
    assign in1502_2 = {s1417[2],s1417[3],s1418[3],s1205[0]};
    CLA_4_c KS_1502(s1502, c1502, in1502_1, in1502_2, s1204[0]);
    wire[3:0] s1503, in1503_1, in1503_2;
    wire c1503;
    assign in1503_1 = {s1419[2],s1211[0],s1212[1],c1210};
    assign in1503_2 = {s1420[1],s1212[0],c1213,s1212[2]};
    CLA_4_c KS_1503(s1503, c1503, in1503_1, in1503_2, c1418);
    wire[3:0] s1504, in1504_1, in1504_2;
    wire c1504;
    assign in1504_1 = {s1419[3],c1419,c1420,s1209[3]};
    assign in1504_2 = {s1420[2],s1420[3],s1421[3],s1212[3]};
    CLA_4_c KS_1504(s1504, c1504, in1504_1, in1504_2, s1213[0]);
    wire[3:0] s1505, in1505_1, in1505_2;
    wire c1505;
    assign in1505_1 = {s1422[2],s1220[0],s1221[1],s1219[2]};
    assign in1505_2 = {s1423[1],s1221[0],c1222,c1221};
    CLA_4_c KS_1505(s1505, c1505, in1505_1, in1505_2, c1421);
    wire[3:0] s1506, in1506_1, in1506_2;
    wire c1506;
    assign in1506_1 = {s1422[3],c1422,c1423,s1218[3]};
    assign in1506_2 = {s1423[2],s1423[3],s1424[3],s1219[3]};
    CLA_4_c KS_1506(s1506, c1506, in1506_1, in1506_2, s1222[0]);
    wire[3:0] s1507, in1507_1, in1507_2;
    wire c1507;
    assign in1507_1 = {s1425[2],s1230[0],c1231,s1230[2]};
    assign in1507_2 = {s1426[1],s1231[0],s1232[1],c1232};
    CLA_4_c KS_1507(s1507, c1507, in1507_1, in1507_2, c1424);
    wire[3:0] s1508, in1508_1, in1508_2;
    wire c1508;
    assign in1508_1 = {s1425[3],c1425,c1426,s1227[3]};
    assign in1508_2 = {s1426[2],s1426[3],s1427[3],c1230};
    CLA_4_c KS_1508(s1508, c1508, in1508_1, in1508_2, s1232[0]);
    wire[3:0] s1509, in1509_1, in1509_2;
    wire c1509;
    assign in1509_1 = {s1428[2],s1238[0],c1239,s1238[2]};
    assign in1509_2 = {s1429[1],s1239[0],s1240[1],c1240};
    CLA_4_c KS_1509(s1509, c1509, in1509_1, in1509_2, c1427);
    wire[3:0] s1510, in1510_1, in1510_2;
    wire c1510;
    assign in1510_1 = {s1428[3],c1428,c1429,s1237[3]};
    assign in1510_2 = {s1429[2],s1429[3],s1430[3],c1238};
    CLA_4_c KS_1510(s1510, c1510, in1510_1, in1510_2, s1240[0]);
    wire[3:0] s1511, in1511_1, in1511_2;
    wire c1511;
    assign in1511_1 = {s1431[2],s1246[0],c1247,s1246[2]};
    assign in1511_2 = {s1432[1],s1247[0],s1248[1],c1248};
    CLA_4_c KS_1511(s1511, c1511, in1511_1, in1511_2, c1430);
    wire[3:0] s1512, in1512_1, in1512_2;
    wire c1512;
    assign in1512_1 = {s1431[3],c1431,c1432,s1245[3]};
    assign in1512_2 = {s1432[2],s1432[3],s1433[3],s1246[3]};
    CLA_4_c KS_1512(s1512, c1512, in1512_1, in1512_2, s1248[0]);
    wire[3:0] s1513, in1513_1, in1513_2;
    wire c1513;
    assign in1513_1 = {s1434[2],s1255[0],s1256[1],c1254};
    assign in1513_2 = {s1435[1],s1256[0],c1257,s1256[2]};
    CLA_4_c KS_1513(s1513, c1513, in1513_1, in1513_2, c1433);
    wire[3:0] s1514, in1514_1, in1514_2;
    wire c1514;
    assign in1514_1 = {s1434[3],c1434,c1435,s1253[3]};
    assign in1514_2 = {s1435[2],s1435[3],s1436[3],c1256};
    CLA_4_c KS_1514(s1514, c1514, in1514_1, in1514_2, s1257[0]);
    wire[3:0] s1515, in1515_1, in1515_2;
    wire c1515;
    assign in1515_1 = {s1437[2],s1263[0],c1264,s1263[2]};
    assign in1515_2 = {s1438[1],s1264[0],s1265[1],c1265};
    CLA_4_c KS_1515(s1515, c1515, in1515_1, in1515_2, c1436);
    wire[3:0] s1516, in1516_1, in1516_2;
    wire c1516;
    assign in1516_1 = {s1437[3],c1437,c1438,s1262[3]};
    assign in1516_2 = {s1438[2],s1438[3],s1439[3],c1263};
    CLA_4_c KS_1516(s1516, c1516, in1516_1, in1516_2, s1265[0]);
    wire[3:0] s1517, in1517_1, in1517_2;
    wire c1517;
    assign in1517_1 = {s1440[2],s1271[0],c1272,s1271[2]};
    assign in1517_2 = {s1441[1],s1272[0],s1273[1],c1273};
    CLA_4_c KS_1517(s1517, c1517, in1517_1, in1517_2, c1439);
    wire[3:0] s1518, in1518_1, in1518_2;
    wire c1518;
    assign in1518_1 = {s1440[3],c1440,c1441,s1270[3]};
    assign in1518_2 = {s1441[2],s1441[3],s1442[3],c1271};
    CLA_4_c KS_1518(s1518, c1518, in1518_1, in1518_2, s1273[0]);
    wire[3:0] s1519, in1519_1, in1519_2;
    wire c1519;
    assign in1519_1 = {s1443[2],s1279[0],c1280,s1279[2]};
    assign in1519_2 = {s1444[1],s1280[0],s1281[1],c1281};
    CLA_4_c KS_1519(s1519, c1519, in1519_1, in1519_2, c1442);
    wire[3:0] s1520, in1520_1, in1520_2;
    wire c1520;
    assign in1520_1 = {s1443[3],c1443,c1444,s1278[3]};
    assign in1520_2 = {s1444[2],s1444[3],s1445[3],s1279[3]};
    CLA_4_c KS_1520(s1520, c1520, in1520_1, in1520_2, s1281[0]);
    wire[3:0] s1521, in1521_1, in1521_2;
    wire c1521;
    assign in1521_1 = {s1446[2],s1289[0],c1290,s1289[2]};
    assign in1521_2 = {s1447[1],s1290[0],s1291[1],c1291};
    CLA_4_c KS_1521(s1521, c1521, in1521_1, in1521_2, c1445);
    wire[3:0] s1522, in1522_1, in1522_2;
    wire c1522;
    assign in1522_1 = {s1446[3],c1446,c1447,s1286[3]};
    assign in1522_2 = {s1447[2],s1447[3],s1448[3],c1289};
    CLA_4_c KS_1522(s1522, c1522, in1522_1, in1522_2, s1291[0]);
    wire[3:0] s1523, in1523_1, in1523_2;
    wire c1523;
    assign in1523_1 = {s1449[2],s1298[0],s1299[1],c1297};
    assign in1523_2 = {s1450[1],s1299[0],c1300,s1299[2]};
    CLA_4_c KS_1523(s1523, c1523, in1523_1, in1523_2, c1448);
    wire[3:0] s1524, in1524_1, in1524_2;
    wire c1524;
    assign in1524_1 = {s1449[3],c1449,c1450,s1296[3]};
    assign in1524_2 = {s1450[2],s1450[3],s1451[3],c1299};
    CLA_4_c KS_1524(s1524, c1524, in1524_1, in1524_2, s1300[0]);
    wire[3:0] s1525, in1525_1, in1525_2;
    wire c1525;
    assign in1525_1 = {s1452[2],s1307[0],s1308[1],c1306};
    assign in1525_2 = {s1453[1],s1308[0],c1309,s1308[2]};
    CLA_4_c KS_1525(s1525, c1525, in1525_1, in1525_2, c1451);
    wire[3:0] s1526, in1526_1, in1526_2;
    wire c1526;
    assign in1526_1 = {s1452[3],c1452,c1453,s1305[3]};
    assign in1526_2 = {s1453[2],s1453[3],s1454[3],s1308[3]};
    CLA_4_c KS_1526(s1526, c1526, in1526_1, in1526_2, s1309[0]);
    wire[3:0] s1527, in1527_1, in1527_2;
    wire c1527;
    assign in1527_1 = {s1455[2],s1316[0],s1317[1],c1315};
    assign in1527_2 = {s1456[1],s1317[0],c1318,s1317[2]};
    CLA_4_c KS_1527(s1527, c1527, in1527_1, in1527_2, c1454);
    wire[3:0] s1528, in1528_1, in1528_2;
    wire c1528;
    assign in1528_1 = {s1455[3],c1455,c1456,s1314[3]};
    assign in1528_2 = {s1456[2],s1456[3],s1457[3],s1317[3]};
    CLA_4_c KS_1528(s1528, c1528, in1528_1, in1528_2, s1318[0]);
    wire[3:0] s1529, in1529_1, in1529_2;
    wire c1529;
    assign in1529_1 = {s1458[2],s1326[0],c1327,s1326[2]};
    assign in1529_2 = {s1459[1],s1327[0],s1328[1],c1328};
    CLA_4_c KS_1529(s1529, c1529, in1529_1, in1529_2, c1457);
    wire[3:0] s1530, in1530_1, in1530_2;
    wire c1530;
    assign in1530_1 = {s1458[3],c1458,c1459,s1323[3]};
    assign in1530_2 = {s1459[2],s1459[3],s1460[3],c1326};
    CLA_4_c KS_1530(s1530, c1530, in1530_1, in1530_2, s1328[0]);
    wire[3:0] s1531, in1531_1, in1531_2;
    wire c1531;
    assign in1531_1 = {s1461[2],s1334[0],c1335,c1334};
    assign in1531_2 = {s1462[1],s1335[0],s1336[1],s1336[2]};
    CLA_4_c KS_1531(s1531, c1531, in1531_1, in1531_2, c1460);
    wire[3:0] s1532, in1532_1, in1532_2;
    wire c1532;
    assign in1532_1 = {s1461[3],c1461,c1462,s1333[3]};
    assign in1532_2 = {s1462[2],s1462[3],s1463[3],c1336};
    CLA_4_c KS_1532(s1532, c1532, in1532_1, in1532_2, s1336[0]);
    wire[3:0] s1533, in1533_1, in1533_2;
    wire c1533;
    assign in1533_1 = {s1464[2],s1343[0],s1344[1],c1342};
    assign in1533_2 = {s1465[1],s1344[0],c1345,s1344[2]};
    CLA_4_c KS_1533(s1533, c1533, in1533_1, in1533_2, c1463);
    wire[3:0] s1534, in1534_1, in1534_2;
    wire c1534;
    assign in1534_1 = {s1464[3],c1464,c1465,s1341[3]};
    assign in1534_2 = {s1465[2],s1465[3],s1466[3],c1344};
    CLA_4_c KS_1534(s1534, c1534, in1534_1, in1534_2, s1345[0]);
    wire[3:0] s1535, in1535_1, in1535_2;
    wire c1535;
    assign in1535_1 = {s1467[2],s1351[0],c1352,s1351[2]};
    assign in1535_2 = {s1468[1],s1352[0],s1353[1],c1353};
    CLA_4_c KS_1535(s1535, c1535, in1535_1, in1535_2, c1466);
    wire[3:0] s1536, in1536_1, in1536_2;
    wire c1536;
    assign in1536_1 = {s1467[3],c1467,c1468,s1350[3]};
    assign in1536_2 = {s1468[2],s1468[3],s1469[3],s1351[3]};
    CLA_4_c KS_1536(s1536, c1536, in1536_1, in1536_2, s1353[0]);
    wire[3:0] s1537, in1537_1, in1537_2;
    wire c1537;
    assign in1537_1 = {s1470[2],s1361[0],c1362,c1361};
    assign in1537_2 = {s1471[1],s1362[0],s1363[1],s1363[2]};
    CLA_4_c KS_1537(s1537, c1537, in1537_1, in1537_2, c1469);
    wire[3:0] s1538, in1538_1, in1538_2;
    wire c1538;
    assign in1538_1 = {s1470[3],c1470,c1471,c1359};
    assign in1538_2 = {s1471[2],s1471[3],s1472[3],s1363[3]};
    CLA_4_c KS_1538(s1538, c1538, in1538_1, in1538_2, s1363[0]);
    wire[3:0] s1539, in1539_1, in1539_2;
    wire c1539;
    assign in1539_1 = {s1473[2],s1371[0],c1372,s1371[2]};
    assign in1539_2 = {s1474[1],s1372[0],s1373[1],c1373};
    CLA_4_c KS_1539(s1539, c1539, in1539_1, in1539_2, c1472);
    wire[3:0] s1540, in1540_1, in1540_2;
    wire c1540;
    assign in1540_1 = {s1473[3],c1473,c1474,s1368[3]};
    assign in1540_2 = {s1474[2],s1474[3],s1475[3],c1371};
    CLA_4_c KS_1540(s1540, c1540, in1540_1, in1540_2, s1373[0]);
    wire[3:0] s1541, in1541_1, in1541_2;
    wire c1541;
    assign in1541_1 = {s1476[2],s1380[0],s1381[1],c1379};
    assign in1541_2 = {s1477[1],s1381[0],c1382,s1381[2]};
    CLA_4_c KS_1541(s1541, c1541, in1541_1, in1541_2, c1475);
    wire[3:0] s1542, in1542_1, in1542_2;
    wire c1542;
    assign in1542_1 = {s1476[3],c1476,c1477,s1378[3]};
    assign in1542_2 = {s1477[2],s1477[3],s1478[3],c1381};
    CLA_4_c KS_1542(s1542, c1542, in1542_1, in1542_2, s1382[0]);
    wire[3:0] s1543, in1543_1, in1543_2;
    wire c1543;
    assign in1543_1 = {s1479[2],s1388[0],c1389,c1388};
    assign in1543_2 = {s1480[1],s1389[0],s1390[1],s1390[2]};
    CLA_4_c KS_1543(s1543, c1543, in1543_1, in1543_2, c1478);
    wire[3:0] s1544, in1544_1, in1544_2;
    wire c1544;
    assign in1544_1 = {s1479[3],c1479,c1480,s1387[3]};
    assign in1544_2 = {s1480[2],s1480[3],s1481[3],c1390};
    CLA_4_c KS_1544(s1544, c1544, in1544_1, in1544_2, s1390[0]);
    wire[3:0] s1545, in1545_1, in1545_2;
    wire c1545;
    assign in1545_1 = {s1482[2],s1397[0],s1398[1],c1396};
    assign in1545_2 = {s1483[1],s1398[0],c1399,s1398[2]};
    CLA_4_c KS_1545(s1545, c1545, in1545_1, in1545_2, c1481);
    wire[3:0] s1546, in1546_1, in1546_2;
    wire c1546;
    assign in1546_1 = {s1482[3],c1482,c1483,s1395[3]};
    assign in1546_2 = {s1483[2],s1483[3],s1484[3],c1398};
    CLA_4_c KS_1546(s1546, c1546, in1546_1, in1546_2, s1399[0]);
    wire[3:0] s1547, in1547_1, in1547_2;
    wire c1547;
    assign in1547_1 = {s1485[2],s1401[0],s1402[1],c1400};
    assign in1547_2 = {s1486[1],s1402[0],c1403,s1402[2]};
    CLA_4_c KS_1547(s1547, c1547, in1547_1, in1547_2, c1484);
    wire[3:0] s1548, in1548_1, in1548_2;
    wire c1548;
    assign in1548_1 = {s1485[3],c1485,c1486,pp63[57]};
    assign in1548_2 = {s1486[2],s1486[3],s1487[3],c1402};
    CLA_4_c KS_1548(s1548, c1548, in1548_1, in1548_2, s1403[0]);
    wire[3:0] s1549, in1549_1, in1549_2;
    wire c1549;
    assign in1549_1 = {s1488[2],pp62[59],pp61[61],pp60[63]};
    assign in1549_2 = {s1489[1],pp63[58],pp62[60],pp61[62]};
    CLA_4_c KS_1549(s1549, c1549, in1549_1, in1549_2, c1487);
    wire[3:0] s1550, in1550_1, in1550_2;
    wire c1550;
    assign in1550_1 = {s1488[3],pp63[59],pp62[61],pp61[63]};
    assign in1550_2 = {c1489,c1488,pp63[60],pp62[62]};
    CLA_4 KS_1550(s1550, c1550, in1550_1, in1550_2);

    /*Stage 7*/
    wire[3:0] s1551, in1551_1, in1551_2;
    wire c1551;
    assign in1551_1 = {pp0[3],pp2[2],pp4[1],pp6[0]};
    assign in1551_2 = {pp1[2],pp3[1],pp5[0],s1404[0]};
    CLA_4 KS_1551(s1551, c1551, in1551_1, in1551_2);
    wire[3:0] s1552, in1552_1, in1552_2;
    wire c1552;
    assign in1552_1 = {s1405[0],s1406[0],s1406[1],s1406[2]};
    assign in1552_2 = {s1491[3],c1491,c1492,s1407[0]};
    CLA_4_c KS_1552(s1552, c1552, in1552_1, in1552_2, s1404[1]);
    wire[3:0] s1553, in1553_1, in1553_2;
    wire c1553;
    assign in1553_1 = {s1408[0],s1409[0],s1409[1],s1409[2]};
    assign in1553_2 = {s1493[3],c1493,c1494,s1410[0]};
    CLA_4_c KS_1553(s1553, c1553, in1553_1, in1553_2, s1407[1]);
    wire[3:0] s1554, in1554_1, in1554_2;
    wire c1554;
    assign in1554_1 = {s1411[0],s1412[0],s1412[1],s1412[2]};
    assign in1554_2 = {s1495[3],c1495,c1496,s1413[0]};
    CLA_4_c KS_1554(s1554, c1554, in1554_1, in1554_2, s1410[1]);
    wire[3:0] s1555, in1555_1, in1555_2;
    wire c1555;
    assign in1555_1 = {s1414[0],s1415[0],s1415[1],s1415[2]};
    assign in1555_2 = {s1497[3],c1497,c1498,s1416[0]};
    CLA_4_c KS_1555(s1555, c1555, in1555_1, in1555_2, s1413[1]);
    wire[3:0] s1556, in1556_1, in1556_2;
    wire c1556;
    assign in1556_1 = {s1417[0],s1418[0],s1418[1],s1418[2]};
    assign in1556_2 = {s1499[3],c1499,c1500,s1419[0]};
    CLA_4_c KS_1556(s1556, c1556, in1556_1, in1556_2, s1416[1]);
    wire[3:0] s1557, in1557_1, in1557_2;
    wire c1557;
    assign in1557_1 = {s1420[0],s1421[0],s1421[1],s1421[2]};
    assign in1557_2 = {s1501[3],c1501,c1502,s1422[0]};
    CLA_4_c KS_1557(s1557, c1557, in1557_1, in1557_2, s1419[1]);
    wire[3:0] s1558, in1558_1, in1558_2;
    wire c1558;
    assign in1558_1 = {s1423[0],s1424[0],s1424[1],s1424[2]};
    assign in1558_2 = {s1503[3],c1503,c1504,s1425[0]};
    CLA_4_c KS_1558(s1558, c1558, in1558_1, in1558_2, s1422[1]);
    wire[3:0] s1559, in1559_1, in1559_2;
    wire c1559;
    assign in1559_1 = {s1426[0],s1427[0],s1427[1],s1427[2]};
    assign in1559_2 = {s1505[3],c1505,c1506,s1428[0]};
    CLA_4_c KS_1559(s1559, c1559, in1559_1, in1559_2, s1425[1]);
    wire[3:0] s1560, in1560_1, in1560_2;
    wire c1560;
    assign in1560_1 = {s1429[0],s1430[0],s1430[1],s1430[2]};
    assign in1560_2 = {s1507[3],c1507,c1508,s1431[0]};
    CLA_4_c KS_1560(s1560, c1560, in1560_1, in1560_2, s1428[1]);
    wire[3:0] s1561, in1561_1, in1561_2;
    wire c1561;
    assign in1561_1 = {s1432[0],s1433[0],s1433[1],s1433[2]};
    assign in1561_2 = {s1509[3],c1509,c1510,s1434[0]};
    CLA_4_c KS_1561(s1561, c1561, in1561_1, in1561_2, s1431[1]);
    wire[3:0] s1562, in1562_1, in1562_2;
    wire c1562;
    assign in1562_1 = {s1435[0],s1436[0],s1436[1],s1436[2]};
    assign in1562_2 = {s1511[3],c1511,c1512,s1437[0]};
    CLA_4_c KS_1562(s1562, c1562, in1562_1, in1562_2, s1434[1]);
    wire[3:0] s1563, in1563_1, in1563_2;
    wire c1563;
    assign in1563_1 = {s1438[0],s1439[0],s1439[1],s1439[2]};
    assign in1563_2 = {s1513[3],c1513,c1514,s1440[0]};
    CLA_4_c KS_1563(s1563, c1563, in1563_1, in1563_2, s1437[1]);
    wire[3:0] s1564, in1564_1, in1564_2;
    wire c1564;
    assign in1564_1 = {s1441[0],s1442[0],s1442[1],s1442[2]};
    assign in1564_2 = {s1515[3],c1515,c1516,s1443[0]};
    CLA_4_c KS_1564(s1564, c1564, in1564_1, in1564_2, s1440[1]);
    wire[3:0] s1565, in1565_1, in1565_2;
    wire c1565;
    assign in1565_1 = {s1444[0],s1445[0],s1445[1],s1445[2]};
    assign in1565_2 = {s1517[3],c1517,c1518,s1446[0]};
    CLA_4_c KS_1565(s1565, c1565, in1565_1, in1565_2, s1443[1]);
    wire[3:0] s1566, in1566_1, in1566_2;
    wire c1566;
    assign in1566_1 = {s1447[0],s1448[0],s1448[1],s1448[2]};
    assign in1566_2 = {s1519[3],c1519,c1520,s1449[0]};
    CLA_4_c KS_1566(s1566, c1566, in1566_1, in1566_2, s1446[1]);
    wire[3:0] s1567, in1567_1, in1567_2;
    wire c1567;
    assign in1567_1 = {s1450[0],s1451[0],s1451[1],s1451[2]};
    assign in1567_2 = {s1521[3],c1521,c1522,s1452[0]};
    CLA_4_c KS_1567(s1567, c1567, in1567_1, in1567_2, s1449[1]);
    wire[3:0] s1568, in1568_1, in1568_2;
    wire c1568;
    assign in1568_1 = {s1453[0],s1454[0],s1454[1],s1454[2]};
    assign in1568_2 = {s1523[3],c1523,c1524,s1455[0]};
    CLA_4_c KS_1568(s1568, c1568, in1568_1, in1568_2, s1452[1]);
    wire[3:0] s1569, in1569_1, in1569_2;
    wire c1569;
    assign in1569_1 = {s1456[0],s1457[0],s1457[1],s1457[2]};
    assign in1569_2 = {s1525[3],c1525,c1526,s1458[0]};
    CLA_4_c KS_1569(s1569, c1569, in1569_1, in1569_2, s1455[1]);
    wire[3:0] s1570, in1570_1, in1570_2;
    wire c1570;
    assign in1570_1 = {s1459[0],s1460[0],s1460[1],s1460[2]};
    assign in1570_2 = {s1527[3],c1527,c1528,s1461[0]};
    CLA_4_c KS_1570(s1570, c1570, in1570_1, in1570_2, s1458[1]);
    wire[3:0] s1571, in1571_1, in1571_2;
    wire c1571;
    assign in1571_1 = {s1462[0],s1463[0],s1463[1],s1463[2]};
    assign in1571_2 = {s1529[3],c1529,c1530,s1464[0]};
    CLA_4_c KS_1571(s1571, c1571, in1571_1, in1571_2, s1461[1]);
    wire[3:0] s1572, in1572_1, in1572_2;
    wire c1572;
    assign in1572_1 = {s1465[0],s1466[0],s1466[1],s1466[2]};
    assign in1572_2 = {s1531[3],c1531,c1532,s1467[0]};
    CLA_4_c KS_1572(s1572, c1572, in1572_1, in1572_2, s1464[1]);
    wire[3:0] s1573, in1573_1, in1573_2;
    wire c1573;
    assign in1573_1 = {s1468[0],s1469[0],s1469[1],s1469[2]};
    assign in1573_2 = {s1533[3],c1533,c1534,s1470[0]};
    CLA_4_c KS_1573(s1573, c1573, in1573_1, in1573_2, s1467[1]);
    wire[3:0] s1574, in1574_1, in1574_2;
    wire c1574;
    assign in1574_1 = {s1471[0],s1472[0],s1472[1],s1472[2]};
    assign in1574_2 = {s1535[3],c1535,c1536,s1473[0]};
    CLA_4_c KS_1574(s1574, c1574, in1574_1, in1574_2, s1470[1]);
    wire[3:0] s1575, in1575_1, in1575_2;
    wire c1575;
    assign in1575_1 = {s1474[0],s1475[0],s1475[1],s1475[2]};
    assign in1575_2 = {s1537[3],c1537,c1538,s1476[0]};
    CLA_4_c KS_1575(s1575, c1575, in1575_1, in1575_2, s1473[1]);
    wire[3:0] s1576, in1576_1, in1576_2;
    wire c1576;
    assign in1576_1 = {s1477[0],s1478[0],s1478[1],s1478[2]};
    assign in1576_2 = {s1539[3],c1539,c1540,s1479[0]};
    CLA_4_c KS_1576(s1576, c1576, in1576_1, in1576_2, s1476[1]);
    wire[3:0] s1577, in1577_1, in1577_2;
    wire c1577;
    assign in1577_1 = {s1480[0],s1481[0],s1481[1],s1481[2]};
    assign in1577_2 = {s1541[3],c1541,c1542,s1482[0]};
    CLA_4_c KS_1577(s1577, c1577, in1577_1, in1577_2, s1479[1]);
    wire[3:0] s1578, in1578_1, in1578_2;
    wire c1578;
    assign in1578_1 = {s1483[0],s1484[0],s1484[1],s1484[2]};
    assign in1578_2 = {s1543[3],c1543,c1544,s1485[0]};
    CLA_4_c KS_1578(s1578, c1578, in1578_1, in1578_2, s1482[1]);
    wire[3:0] s1579, in1579_1, in1579_2;
    wire c1579;
    assign in1579_1 = {s1486[0],s1487[0],s1487[1],s1487[2]};
    assign in1579_2 = {s1545[3],c1545,c1546,s1488[0]};
    CLA_4_c KS_1579(s1579, c1579, in1579_1, in1579_2, s1485[1]);
    wire[3:0] s1580, in1580_1, in1580_2;
    wire c1580;
    assign in1580_1 = {s1489[0],s1490[0],s1490[1],s1490[2]};
    assign in1580_2 = {s1547[3],c1547,c1548,s1549[2]};
    CLA_4_c KS_1580(s1580, c1580, in1580_1, in1580_2, s1488[1]);
    wire[2:0] s1581, in1581_1, in1581_2;
    wire c1581;
    assign in1581_1 = {c1490,pp63[61],pp62[63]};
    assign in1581_2 = {s1549[3],c1549,pp63[62]};
    CLA_3 KS_1581(s1581, c1581, in1581_1, in1581_2);

    /*Stage 8*/
    wire[3:0] s1582, in1582_1, in1582_2;
    wire c1582;
    assign in1582_1 = {pp0[2],pp2[1],pp4[0],s1491[1]};
    assign in1582_2 = {pp1[1],pp3[0],s1491[0],s1492[0]};
    CLA_4 KS_1582(s1582, c1582, in1582_1, in1582_2);
    wire[3:0] s1583, in1583_1, in1583_2;
    wire c1583;
    assign in1583_1 = {s1492[1],s1492[2],s1492[3],s1493[1]};
    assign in1583_2 = {s1551[3],c1551,s1493[0],s1494[0]};
    CLA_4_c KS_1583(s1583, c1583, in1583_1, in1583_2, s1491[2]);
    wire[3:0] s1584, in1584_1, in1584_2;
    wire c1584;
    assign in1584_1 = {s1494[1],s1494[2],s1494[3],s1495[1]};
    assign in1584_2 = {s1552[3],c1552,s1495[0],s1496[0]};
    CLA_4_c KS_1584(s1584, c1584, in1584_1, in1584_2, s1493[2]);
    wire[3:0] s1585, in1585_1, in1585_2;
    wire c1585;
    assign in1585_1 = {s1496[1],s1496[2],s1496[3],s1497[1]};
    assign in1585_2 = {s1553[3],c1553,s1497[0],s1498[0]};
    CLA_4_c KS_1585(s1585, c1585, in1585_1, in1585_2, s1495[2]);
    wire[3:0] s1586, in1586_1, in1586_2;
    wire c1586;
    assign in1586_1 = {s1498[1],s1498[2],s1498[3],s1499[1]};
    assign in1586_2 = {s1554[3],c1554,s1499[0],s1500[0]};
    CLA_4_c KS_1586(s1586, c1586, in1586_1, in1586_2, s1497[2]);
    wire[3:0] s1587, in1587_1, in1587_2;
    wire c1587;
    assign in1587_1 = {s1500[1],s1500[2],s1500[3],s1501[1]};
    assign in1587_2 = {s1555[3],c1555,s1501[0],s1502[0]};
    CLA_4_c KS_1587(s1587, c1587, in1587_1, in1587_2, s1499[2]);
    wire[3:0] s1588, in1588_1, in1588_2;
    wire c1588;
    assign in1588_1 = {s1502[1],s1502[2],s1502[3],s1503[1]};
    assign in1588_2 = {s1556[3],c1556,s1503[0],s1504[0]};
    CLA_4_c KS_1588(s1588, c1588, in1588_1, in1588_2, s1501[2]);
    wire[3:0] s1589, in1589_1, in1589_2;
    wire c1589;
    assign in1589_1 = {s1504[1],s1504[2],s1504[3],s1505[1]};
    assign in1589_2 = {s1557[3],c1557,s1505[0],s1506[0]};
    CLA_4_c KS_1589(s1589, c1589, in1589_1, in1589_2, s1503[2]);
    wire[3:0] s1590, in1590_1, in1590_2;
    wire c1590;
    assign in1590_1 = {s1506[1],s1506[2],s1506[3],s1507[1]};
    assign in1590_2 = {s1558[3],c1558,s1507[0],s1508[0]};
    CLA_4_c KS_1590(s1590, c1590, in1590_1, in1590_2, s1505[2]);
    wire[3:0] s1591, in1591_1, in1591_2;
    wire c1591;
    assign in1591_1 = {s1508[1],s1508[2],s1508[3],s1509[1]};
    assign in1591_2 = {s1559[3],c1559,s1509[0],s1510[0]};
    CLA_4_c KS_1591(s1591, c1591, in1591_1, in1591_2, s1507[2]);
    wire[3:0] s1592, in1592_1, in1592_2;
    wire c1592;
    assign in1592_1 = {s1510[1],s1510[2],s1510[3],s1511[1]};
    assign in1592_2 = {s1560[3],c1560,s1511[0],s1512[0]};
    CLA_4_c KS_1592(s1592, c1592, in1592_1, in1592_2, s1509[2]);
    wire[3:0] s1593, in1593_1, in1593_2;
    wire c1593;
    assign in1593_1 = {s1512[1],s1512[2],s1512[3],s1513[1]};
    assign in1593_2 = {s1561[3],c1561,s1513[0],s1514[0]};
    CLA_4_c KS_1593(s1593, c1593, in1593_1, in1593_2, s1511[2]);
    wire[3:0] s1594, in1594_1, in1594_2;
    wire c1594;
    assign in1594_1 = {s1514[1],s1514[2],s1514[3],s1515[1]};
    assign in1594_2 = {s1562[3],c1562,s1515[0],s1516[0]};
    CLA_4_c KS_1594(s1594, c1594, in1594_1, in1594_2, s1513[2]);
    wire[3:0] s1595, in1595_1, in1595_2;
    wire c1595;
    assign in1595_1 = {s1516[1],s1516[2],s1516[3],s1517[1]};
    assign in1595_2 = {s1563[3],c1563,s1517[0],s1518[0]};
    CLA_4_c KS_1595(s1595, c1595, in1595_1, in1595_2, s1515[2]);
    wire[3:0] s1596, in1596_1, in1596_2;
    wire c1596;
    assign in1596_1 = {s1518[1],s1518[2],s1518[3],s1519[1]};
    assign in1596_2 = {s1564[3],c1564,s1519[0],s1520[0]};
    CLA_4_c KS_1596(s1596, c1596, in1596_1, in1596_2, s1517[2]);
    wire[3:0] s1597, in1597_1, in1597_2;
    wire c1597;
    assign in1597_1 = {s1520[1],s1520[2],s1520[3],s1521[1]};
    assign in1597_2 = {s1565[3],c1565,s1521[0],s1522[0]};
    CLA_4_c KS_1597(s1597, c1597, in1597_1, in1597_2, s1519[2]);
    wire[3:0] s1598, in1598_1, in1598_2;
    wire c1598;
    assign in1598_1 = {s1522[1],s1522[2],s1522[3],s1523[1]};
    assign in1598_2 = {s1566[3],c1566,s1523[0],s1524[0]};
    CLA_4_c KS_1598(s1598, c1598, in1598_1, in1598_2, s1521[2]);
    wire[3:0] s1599, in1599_1, in1599_2;
    wire c1599;
    assign in1599_1 = {s1524[1],s1524[2],s1524[3],s1525[1]};
    assign in1599_2 = {s1567[3],c1567,s1525[0],s1526[0]};
    CLA_4_c KS_1599(s1599, c1599, in1599_1, in1599_2, s1523[2]);
    wire[3:0] s1600, in1600_1, in1600_2;
    wire c1600;
    assign in1600_1 = {s1526[1],s1526[2],s1526[3],s1527[1]};
    assign in1600_2 = {s1568[3],c1568,s1527[0],s1528[0]};
    CLA_4_c KS_1600(s1600, c1600, in1600_1, in1600_2, s1525[2]);
    wire[3:0] s1601, in1601_1, in1601_2;
    wire c1601;
    assign in1601_1 = {s1528[1],s1528[2],s1528[3],s1529[1]};
    assign in1601_2 = {s1569[3],c1569,s1529[0],s1530[0]};
    CLA_4_c KS_1601(s1601, c1601, in1601_1, in1601_2, s1527[2]);
    wire[3:0] s1602, in1602_1, in1602_2;
    wire c1602;
    assign in1602_1 = {s1530[1],s1530[2],s1530[3],s1531[1]};
    assign in1602_2 = {s1570[3],c1570,s1531[0],s1532[0]};
    CLA_4_c KS_1602(s1602, c1602, in1602_1, in1602_2, s1529[2]);
    wire[3:0] s1603, in1603_1, in1603_2;
    wire c1603;
    assign in1603_1 = {s1532[1],s1532[2],s1532[3],s1533[1]};
    assign in1603_2 = {s1571[3],c1571,s1533[0],s1534[0]};
    CLA_4_c KS_1603(s1603, c1603, in1603_1, in1603_2, s1531[2]);
    wire[3:0] s1604, in1604_1, in1604_2;
    wire c1604;
    assign in1604_1 = {s1534[1],s1534[2],s1534[3],s1535[1]};
    assign in1604_2 = {s1572[3],c1572,s1535[0],s1536[0]};
    CLA_4_c KS_1604(s1604, c1604, in1604_1, in1604_2, s1533[2]);
    wire[3:0] s1605, in1605_1, in1605_2;
    wire c1605;
    assign in1605_1 = {s1536[1],s1536[2],s1536[3],s1537[1]};
    assign in1605_2 = {s1573[3],c1573,s1537[0],s1538[0]};
    CLA_4_c KS_1605(s1605, c1605, in1605_1, in1605_2, s1535[2]);
    wire[3:0] s1606, in1606_1, in1606_2;
    wire c1606;
    assign in1606_1 = {s1538[1],s1538[2],s1538[3],s1539[1]};
    assign in1606_2 = {s1574[3],c1574,s1539[0],s1540[0]};
    CLA_4_c KS_1606(s1606, c1606, in1606_1, in1606_2, s1537[2]);
    wire[3:0] s1607, in1607_1, in1607_2;
    wire c1607;
    assign in1607_1 = {s1540[1],s1540[2],s1540[3],s1541[1]};
    assign in1607_2 = {s1575[3],c1575,s1541[0],s1542[0]};
    CLA_4_c KS_1607(s1607, c1607, in1607_1, in1607_2, s1539[2]);
    wire[3:0] s1608, in1608_1, in1608_2;
    wire c1608;
    assign in1608_1 = {s1542[1],s1542[2],s1542[3],s1543[1]};
    assign in1608_2 = {s1576[3],c1576,s1543[0],s1544[0]};
    CLA_4_c KS_1608(s1608, c1608, in1608_1, in1608_2, s1541[2]);
    wire[3:0] s1609, in1609_1, in1609_2;
    wire c1609;
    assign in1609_1 = {s1544[1],s1544[2],s1544[3],s1545[1]};
    assign in1609_2 = {s1577[3],c1577,s1545[0],s1546[0]};
    CLA_4_c KS_1609(s1609, c1609, in1609_1, in1609_2, s1543[2]);
    wire[3:0] s1610, in1610_1, in1610_2;
    wire c1610;
    assign in1610_1 = {s1546[1],s1546[2],s1546[3],s1547[1]};
    assign in1610_2 = {s1578[3],c1578,s1547[0],s1548[0]};
    CLA_4_c KS_1610(s1610, c1610, in1610_1, in1610_2, s1545[2]);
    wire[3:0] s1611, in1611_1, in1611_2;
    wire c1611;
    assign in1611_1 = {s1548[1],s1548[2],s1548[3],s1549[1]};
    assign in1611_2 = {s1579[3],c1579,s1549[0],s1550[0]};
    CLA_4_c KS_1611(s1611, c1611, in1611_1, in1611_2, s1547[2]);
    wire[3:0] s1612, in1612_1, in1612_2;
    wire c1612;
    assign in1612_1 = {s1550[1],s1550[2],s1550[3],c1550};
    assign in1612_2 = {s1580[3],c1580,s1581[1],s1581[2]};
    CLA_4 KS_1612(s1612, c1612, in1612_1, in1612_2);


    /*Final Stage 8*/
    wire[125:0] s, in_1, in_2;
    wire c;
    assign in_1 = {pp0[1],pp2[0],s1551[0],s1551[1],s1551[2],c1582,s1552[0],s1552[1],s1552[2],c1583,s1553[0],s1553[1],s1553[2],c1584,s1554[0],s1554[1],s1554[2],c1585,s1555[0],s1555[1],s1555[2],c1586,s1556[0],s1556[1],s1556[2],c1587,s1557[0],s1557[1],s1557[2],c1588,s1558[0],s1558[1],s1558[2],c1589,s1559[0],s1559[1],s1559[2],c1590,s1560[0],s1560[1],s1560[2],c1591,s1561[0],s1561[1],s1561[2],c1592,s1562[0],s1562[1],s1562[2],c1593,s1563[0],s1563[1],s1563[2],c1594,s1564[0],s1564[1],s1564[2],c1595,s1565[0],s1565[1],s1565[2],c1596,s1566[0],s1566[1],s1566[2],c1597,s1567[0],s1567[1],s1567[2],c1598,s1568[0],s1568[1],s1568[2],c1599,s1569[0],s1569[1],s1569[2],c1600,s1570[0],s1570[1],s1570[2],c1601,s1571[0],s1571[1],s1571[2],c1602,s1572[0],s1572[1],s1572[2],c1603,s1573[0],s1573[1],s1573[2],c1604,s1574[0],s1574[1],s1574[2],c1605,s1575[0],s1575[1],s1575[2],c1606,s1576[0],s1576[1],s1576[2],c1607,s1577[0],s1577[1],s1577[2],c1608,s1578[0],s1578[1],s1578[2],c1609,s1579[0],s1579[1],s1579[2],c1610,s1580[0],s1580[1],s1580[2],c1611,s1581[0],s1612[2],s1612[3],c1612};
    assign in_2 = {pp1[0],s1582[0],s1582[1],s1582[2],s1582[3],s1583[0],s1583[1],s1583[2],s1583[3],s1584[0],s1584[1],s1584[2],s1584[3],s1585[0],s1585[1],s1585[2],s1585[3],s1586[0],s1586[1],s1586[2],s1586[3],s1587[0],s1587[1],s1587[2],s1587[3],s1588[0],s1588[1],s1588[2],s1588[3],s1589[0],s1589[1],s1589[2],s1589[3],s1590[0],s1590[1],s1590[2],s1590[3],s1591[0],s1591[1],s1591[2],s1591[3],s1592[0],s1592[1],s1592[2],s1592[3],s1593[0],s1593[1],s1593[2],s1593[3],s1594[0],s1594[1],s1594[2],s1594[3],s1595[0],s1595[1],s1595[2],s1595[3],s1596[0],s1596[1],s1596[2],s1596[3],s1597[0],s1597[1],s1597[2],s1597[3],s1598[0],s1598[1],s1598[2],s1598[3],s1599[0],s1599[1],s1599[2],s1599[3],s1600[0],s1600[1],s1600[2],s1600[3],s1601[0],s1601[1],s1601[2],s1601[3],s1602[0],s1602[1],s1602[2],s1602[3],s1603[0],s1603[1],s1603[2],s1603[3],s1604[0],s1604[1],s1604[2],s1604[3],s1605[0],s1605[1],s1605[2],s1605[3],s1606[0],s1606[1],s1606[2],s1606[3],s1607[0],s1607[1],s1607[2],s1607[3],s1608[0],s1608[1],s1608[2],s1608[3],s1609[0],s1609[1],s1609[2],s1609[3],s1610[0],s1610[1],s1610[2],s1610[3],s1611[0],s1611[1],s1611[2],s1611[3],s1612[0],s1612[1],1'b0,1'b0,1'b0};
    CLA_126(s, c, in_1, in_2);

    assign product[0] = pp0[0];
    assign product[1] = s[0];
    assign product[2] = s[1];
    assign product[3] = s[2];
    assign product[4] = s[3];
    assign product[5] = s[4];
    assign product[6] = s[5];
    assign product[7] = s[6];
    assign product[8] = s[7];
    assign product[9] = s[8];
    assign product[10] = s[9];
    assign product[11] = s[10];
    assign product[12] = s[11];
    assign product[13] = s[12];
    assign product[14] = s[13];
    assign product[15] = s[14];
    assign product[16] = s[15];
    assign product[17] = s[16];
    assign product[18] = s[17];
    assign product[19] = s[18];
    assign product[20] = s[19];
    assign product[21] = s[20];
    assign product[22] = s[21];
    assign product[23] = s[22];
    assign product[24] = s[23];
    assign product[25] = s[24];
    assign product[26] = s[25];
    assign product[27] = s[26];
    assign product[28] = s[27];
    assign product[29] = s[28];
    assign product[30] = s[29];
    assign product[31] = s[30];
    assign product[32] = s[31];
    assign product[33] = s[32];
    assign product[34] = s[33];
    assign product[35] = s[34];
    assign product[36] = s[35];
    assign product[37] = s[36];
    assign product[38] = s[37];
    assign product[39] = s[38];
    assign product[40] = s[39];
    assign product[41] = s[40];
    assign product[42] = s[41];
    assign product[43] = s[42];
    assign product[44] = s[43];
    assign product[45] = s[44];
    assign product[46] = s[45];
    assign product[47] = s[46];
    assign product[48] = s[47];
    assign product[49] = s[48];
    assign product[50] = s[49];
    assign product[51] = s[50];
    assign product[52] = s[51];
    assign product[53] = s[52];
    assign product[54] = s[53];
    assign product[55] = s[54];
    assign product[56] = s[55];
    assign product[57] = s[56];
    assign product[58] = s[57];
    assign product[59] = s[58];
    assign product[60] = s[59];
    assign product[61] = s[60];
    assign product[62] = s[61];
    assign product[63] = s[62];
    assign product[64] = s[63];
    assign product[65] = s[64];
    assign product[66] = s[65];
    assign product[67] = s[66];
    assign product[68] = s[67];
    assign product[69] = s[68];
    assign product[70] = s[69];
    assign product[71] = s[70];
    assign product[72] = s[71];
    assign product[73] = s[72];
    assign product[74] = s[73];
    assign product[75] = s[74];
    assign product[76] = s[75];
    assign product[77] = s[76];
    assign product[78] = s[77];
    assign product[79] = s[78];
    assign product[80] = s[79];
    assign product[81] = s[80];
    assign product[82] = s[81];
    assign product[83] = s[82];
    assign product[84] = s[83];
    assign product[85] = s[84];
    assign product[86] = s[85];
    assign product[87] = s[86];
    assign product[88] = s[87];
    assign product[89] = s[88];
    assign product[90] = s[89];
    assign product[91] = s[90];
    assign product[92] = s[91];
    assign product[93] = s[92];
    assign product[94] = s[93];
    assign product[95] = s[94];
    assign product[96] = s[95];
    assign product[97] = s[96];
    assign product[98] = s[97];
    assign product[99] = s[98];
    assign product[100] = s[99];
    assign product[101] = s[100];
    assign product[102] = s[101];
    assign product[103] = s[102];
    assign product[104] = s[103];
    assign product[105] = s[104];
    assign product[106] = s[105];
    assign product[107] = s[106];
    assign product[108] = s[107];
    assign product[109] = s[108];
    assign product[110] = s[109];
    assign product[111] = s[110];
    assign product[112] = s[111];
    assign product[113] = s[112];
    assign product[114] = s[113];
    assign product[115] = s[114];
    assign product[116] = s[115];
    assign product[117] = s[116];
    assign product[118] = s[117];
    assign product[119] = s[118];
    assign product[120] = s[119];
    assign product[121] = s[120];
    assign product[122] = s[121];
    assign product[123] = s[122];
    assign product[124] = s[123];
    assign product[125] = s[124];
    assign product[126] = s[125];
    assign product[127] = c;
endmodule


module CLA_2(output [1:0] sum, output cout, input [1:0] in1, input [1:0] in2);

    wire[1:0] G;
    wire[1:0] C;
    wire[1:0] P;

    assign G[0] = in1[1] & in2[1];
    assign P[0] = in1[1] ^ in2[1];
    assign G[1] = in1[0] & in2[0];
    assign P[1] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign cout = G[1] | (P[1] & C[1]);
    assign sum = P ^ C;
endmodule


module CLA_2_c(output [1:0] sum,
            output cout,
            input [1:0] in1, in2,
            input cin);

    wire [1:0] G; /* Generate */
    wire [1:0] P; /* Propagate */
    wire [1:0] C; /* Carry */

    assign G[0] = in1[1] & in2[1]; /*Generate    Gi = Ai * Bi */
    assign G[1] = in1[0] & in2[0];

    assign P[0] = in1[1] ^ in2[1];
    assign P[1] = in1[0] ^ in2[0];

    assign C[0] = cin;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign cout = G[1] | (P[1] & C[1]);
    assign sum = P ^ C;
endmodule


module CLA_3(output [2:0] sum, output cout, input [2:0] in1, input [2:0] in2);

    wire[2:0] G;
    wire[2:0] C;
    wire[2:0] P;

    assign G[0] = in1[2] & in2[2];
    assign P[0] = in1[2] ^ in2[2];
    assign G[1] = in1[1] & in2[1];
    assign P[1] = in1[1] ^ in2[1];
    assign G[2] = in1[0] & in2[0];
    assign P[2] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign cout = G[2] | (P[2] & C[2]);
    assign sum = P ^ C;
endmodule

module CLA_3_c(output [2:0] sum, output cout, input [2:0] in1, input [2:0] in2, input cin);

    wire[2:0] G;
    wire[2:0] C;
    wire[2:0] P;

    assign G[0] = in1[2] & in2[2];
    assign P[0] = in1[2] ^ in2[2];
    assign G[1] = in1[1] & in2[1];
    assign P[1] = in1[1] ^ in2[1];
    assign G[2] = in1[0] & in2[0];
    assign P[2] = in1[0] ^ in2[0];


    assign C[0] = cin;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign cout = G[2] | (P[2] & C[2]);
    assign sum = P ^ C;
endmodule

module CLA_4(output [3:0] sum,
            output cout,
            input [3:0] in1, in2);

    wire [3:0] G; /* Generate */
    wire [3:0] P; /* Propagate */
    wire [3:0] C; /* Carry */

    assign G[0] = in1[3] & in2[3]; /*Generate    Gi = Ai * Bi */
    assign G[1] = in1[2] & in2[2];
    assign G[2] = in1[1] & in2[1];
    assign G[3] = in1[0] & in2[0];
    assign P[0] = in1[3] ^ in2[3]; /*Propagate   Pi = Ai + Bi */
    assign P[1] = in1[2] ^ in2[2];
    assign P[2] = in1[1] ^ in2[1];
    assign P[3] = in1[0] ^ in2[0];

    assign C[0] = 0;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign cout = G[3] | (P[3] & C[3]);
    assign sum = P ^ C;
endmodule

module CLA_4_c(output [3:0] sum,
            output cout,
            input [3:0] in1, in2,
            input cin);

    wire [3:0] G; /* Generate */
    wire [3:0] P; /* Propagate */
    wire [3:0] C; /* Carry */

    assign G[0] = in1[3] & in2[3]; /*Generate    Gi = Ai * Bi */
    assign G[1] = in1[2] & in2[2];
    assign G[2] = in1[1] & in2[1];
    assign G[3] = in1[0] & in2[0];
    assign P[0] = in1[3] ^ in2[3]; /*Propagate   Pi = Ai + Bi */
    assign P[1] = in1[2] ^ in2[2];
    assign P[2] = in1[1] ^ in2[1];
    assign P[3] = in1[0] ^ in2[0];

    assign C[0] = cin;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign cout = G[3] | (P[3] & C[3]);
    assign sum = P ^ C;
endmodule

module Half_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2);
    xor(sum, in1, in2);
    and(cout, in1, in2);
endmodule

module Full_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2,
                  input wire cin);
    wire temp1;
    wire temp2;
    wire temp3;
    xor(sum, in1, in2, cin);
    and(temp1,in1,in2);
    and(temp2,in1,cin);
    and(temp3,in2,cin);
    or(cout,temp1,temp2,temp3);
endmodule


module CLA_126(output [125:0] sum, output cout, input [125:0] in1, input [125:0] in2);

    wire[125:0] G;
    wire[125:0] C;
    wire[125:0] P;

    assign G[0] = in1[125] & in2[125];
    assign P[0] = in1[125] ^ in2[125];
    assign G[1] = in1[124] & in2[124];
    assign P[1] = in1[124] ^ in2[124];
    assign G[2] = in1[123] & in2[123];
    assign P[2] = in1[123] ^ in2[123];
    assign G[3] = in1[122] & in2[122];
    assign P[3] = in1[122] ^ in2[122];
    assign G[4] = in1[121] & in2[121];
    assign P[4] = in1[121] ^ in2[121];
    assign G[5] = in1[120] & in2[120];
    assign P[5] = in1[120] ^ in2[120];
    assign G[6] = in1[119] & in2[119];
    assign P[6] = in1[119] ^ in2[119];
    assign G[7] = in1[118] & in2[118];
    assign P[7] = in1[118] ^ in2[118];
    assign G[8] = in1[117] & in2[117];
    assign P[8] = in1[117] ^ in2[117];
    assign G[9] = in1[116] & in2[116];
    assign P[9] = in1[116] ^ in2[116];
    assign G[10] = in1[115] & in2[115];
    assign P[10] = in1[115] ^ in2[115];
    assign G[11] = in1[114] & in2[114];
    assign P[11] = in1[114] ^ in2[114];
    assign G[12] = in1[113] & in2[113];
    assign P[12] = in1[113] ^ in2[113];
    assign G[13] = in1[112] & in2[112];
    assign P[13] = in1[112] ^ in2[112];
    assign G[14] = in1[111] & in2[111];
    assign P[14] = in1[111] ^ in2[111];
    assign G[15] = in1[110] & in2[110];
    assign P[15] = in1[110] ^ in2[110];
    assign G[16] = in1[109] & in2[109];
    assign P[16] = in1[109] ^ in2[109];
    assign G[17] = in1[108] & in2[108];
    assign P[17] = in1[108] ^ in2[108];
    assign G[18] = in1[107] & in2[107];
    assign P[18] = in1[107] ^ in2[107];
    assign G[19] = in1[106] & in2[106];
    assign P[19] = in1[106] ^ in2[106];
    assign G[20] = in1[105] & in2[105];
    assign P[20] = in1[105] ^ in2[105];
    assign G[21] = in1[104] & in2[104];
    assign P[21] = in1[104] ^ in2[104];
    assign G[22] = in1[103] & in2[103];
    assign P[22] = in1[103] ^ in2[103];
    assign G[23] = in1[102] & in2[102];
    assign P[23] = in1[102] ^ in2[102];
    assign G[24] = in1[101] & in2[101];
    assign P[24] = in1[101] ^ in2[101];
    assign G[25] = in1[100] & in2[100];
    assign P[25] = in1[100] ^ in2[100];
    assign G[26] = in1[99] & in2[99];
    assign P[26] = in1[99] ^ in2[99];
    assign G[27] = in1[98] & in2[98];
    assign P[27] = in1[98] ^ in2[98];
    assign G[28] = in1[97] & in2[97];
    assign P[28] = in1[97] ^ in2[97];
    assign G[29] = in1[96] & in2[96];
    assign P[29] = in1[96] ^ in2[96];
    assign G[30] = in1[95] & in2[95];
    assign P[30] = in1[95] ^ in2[95];
    assign G[31] = in1[94] & in2[94];
    assign P[31] = in1[94] ^ in2[94];
    assign G[32] = in1[93] & in2[93];
    assign P[32] = in1[93] ^ in2[93];
    assign G[33] = in1[92] & in2[92];
    assign P[33] = in1[92] ^ in2[92];
    assign G[34] = in1[91] & in2[91];
    assign P[34] = in1[91] ^ in2[91];
    assign G[35] = in1[90] & in2[90];
    assign P[35] = in1[90] ^ in2[90];
    assign G[36] = in1[89] & in2[89];
    assign P[36] = in1[89] ^ in2[89];
    assign G[37] = in1[88] & in2[88];
    assign P[37] = in1[88] ^ in2[88];
    assign G[38] = in1[87] & in2[87];
    assign P[38] = in1[87] ^ in2[87];
    assign G[39] = in1[86] & in2[86];
    assign P[39] = in1[86] ^ in2[86];
    assign G[40] = in1[85] & in2[85];
    assign P[40] = in1[85] ^ in2[85];
    assign G[41] = in1[84] & in2[84];
    assign P[41] = in1[84] ^ in2[84];
    assign G[42] = in1[83] & in2[83];
    assign P[42] = in1[83] ^ in2[83];
    assign G[43] = in1[82] & in2[82];
    assign P[43] = in1[82] ^ in2[82];
    assign G[44] = in1[81] & in2[81];
    assign P[44] = in1[81] ^ in2[81];
    assign G[45] = in1[80] & in2[80];
    assign P[45] = in1[80] ^ in2[80];
    assign G[46] = in1[79] & in2[79];
    assign P[46] = in1[79] ^ in2[79];
    assign G[47] = in1[78] & in2[78];
    assign P[47] = in1[78] ^ in2[78];
    assign G[48] = in1[77] & in2[77];
    assign P[48] = in1[77] ^ in2[77];
    assign G[49] = in1[76] & in2[76];
    assign P[49] = in1[76] ^ in2[76];
    assign G[50] = in1[75] & in2[75];
    assign P[50] = in1[75] ^ in2[75];
    assign G[51] = in1[74] & in2[74];
    assign P[51] = in1[74] ^ in2[74];
    assign G[52] = in1[73] & in2[73];
    assign P[52] = in1[73] ^ in2[73];
    assign G[53] = in1[72] & in2[72];
    assign P[53] = in1[72] ^ in2[72];
    assign G[54] = in1[71] & in2[71];
    assign P[54] = in1[71] ^ in2[71];
    assign G[55] = in1[70] & in2[70];
    assign P[55] = in1[70] ^ in2[70];
    assign G[56] = in1[69] & in2[69];
    assign P[56] = in1[69] ^ in2[69];
    assign G[57] = in1[68] & in2[68];
    assign P[57] = in1[68] ^ in2[68];
    assign G[58] = in1[67] & in2[67];
    assign P[58] = in1[67] ^ in2[67];
    assign G[59] = in1[66] & in2[66];
    assign P[59] = in1[66] ^ in2[66];
    assign G[60] = in1[65] & in2[65];
    assign P[60] = in1[65] ^ in2[65];
    assign G[61] = in1[64] & in2[64];
    assign P[61] = in1[64] ^ in2[64];
    assign G[62] = in1[63] & in2[63];
    assign P[62] = in1[63] ^ in2[63];
    assign G[63] = in1[62] & in2[62];
    assign P[63] = in1[62] ^ in2[62];
    assign G[64] = in1[61] & in2[61];
    assign P[64] = in1[61] ^ in2[61];
    assign G[65] = in1[60] & in2[60];
    assign P[65] = in1[60] ^ in2[60];
    assign G[66] = in1[59] & in2[59];
    assign P[66] = in1[59] ^ in2[59];
    assign G[67] = in1[58] & in2[58];
    assign P[67] = in1[58] ^ in2[58];
    assign G[68] = in1[57] & in2[57];
    assign P[68] = in1[57] ^ in2[57];
    assign G[69] = in1[56] & in2[56];
    assign P[69] = in1[56] ^ in2[56];
    assign G[70] = in1[55] & in2[55];
    assign P[70] = in1[55] ^ in2[55];
    assign G[71] = in1[54] & in2[54];
    assign P[71] = in1[54] ^ in2[54];
    assign G[72] = in1[53] & in2[53];
    assign P[72] = in1[53] ^ in2[53];
    assign G[73] = in1[52] & in2[52];
    assign P[73] = in1[52] ^ in2[52];
    assign G[74] = in1[51] & in2[51];
    assign P[74] = in1[51] ^ in2[51];
    assign G[75] = in1[50] & in2[50];
    assign P[75] = in1[50] ^ in2[50];
    assign G[76] = in1[49] & in2[49];
    assign P[76] = in1[49] ^ in2[49];
    assign G[77] = in1[48] & in2[48];
    assign P[77] = in1[48] ^ in2[48];
    assign G[78] = in1[47] & in2[47];
    assign P[78] = in1[47] ^ in2[47];
    assign G[79] = in1[46] & in2[46];
    assign P[79] = in1[46] ^ in2[46];
    assign G[80] = in1[45] & in2[45];
    assign P[80] = in1[45] ^ in2[45];
    assign G[81] = in1[44] & in2[44];
    assign P[81] = in1[44] ^ in2[44];
    assign G[82] = in1[43] & in2[43];
    assign P[82] = in1[43] ^ in2[43];
    assign G[83] = in1[42] & in2[42];
    assign P[83] = in1[42] ^ in2[42];
    assign G[84] = in1[41] & in2[41];
    assign P[84] = in1[41] ^ in2[41];
    assign G[85] = in1[40] & in2[40];
    assign P[85] = in1[40] ^ in2[40];
    assign G[86] = in1[39] & in2[39];
    assign P[86] = in1[39] ^ in2[39];
    assign G[87] = in1[38] & in2[38];
    assign P[87] = in1[38] ^ in2[38];
    assign G[88] = in1[37] & in2[37];
    assign P[88] = in1[37] ^ in2[37];
    assign G[89] = in1[36] & in2[36];
    assign P[89] = in1[36] ^ in2[36];
    assign G[90] = in1[35] & in2[35];
    assign P[90] = in1[35] ^ in2[35];
    assign G[91] = in1[34] & in2[34];
    assign P[91] = in1[34] ^ in2[34];
    assign G[92] = in1[33] & in2[33];
    assign P[92] = in1[33] ^ in2[33];
    assign G[93] = in1[32] & in2[32];
    assign P[93] = in1[32] ^ in2[32];
    assign G[94] = in1[31] & in2[31];
    assign P[94] = in1[31] ^ in2[31];
    assign G[95] = in1[30] & in2[30];
    assign P[95] = in1[30] ^ in2[30];
    assign G[96] = in1[29] & in2[29];
    assign P[96] = in1[29] ^ in2[29];
    assign G[97] = in1[28] & in2[28];
    assign P[97] = in1[28] ^ in2[28];
    assign G[98] = in1[27] & in2[27];
    assign P[98] = in1[27] ^ in2[27];
    assign G[99] = in1[26] & in2[26];
    assign P[99] = in1[26] ^ in2[26];
    assign G[100] = in1[25] & in2[25];
    assign P[100] = in1[25] ^ in2[25];
    assign G[101] = in1[24] & in2[24];
    assign P[101] = in1[24] ^ in2[24];
    assign G[102] = in1[23] & in2[23];
    assign P[102] = in1[23] ^ in2[23];
    assign G[103] = in1[22] & in2[22];
    assign P[103] = in1[22] ^ in2[22];
    assign G[104] = in1[21] & in2[21];
    assign P[104] = in1[21] ^ in2[21];
    assign G[105] = in1[20] & in2[20];
    assign P[105] = in1[20] ^ in2[20];
    assign G[106] = in1[19] & in2[19];
    assign P[106] = in1[19] ^ in2[19];
    assign G[107] = in1[18] & in2[18];
    assign P[107] = in1[18] ^ in2[18];
    assign G[108] = in1[17] & in2[17];
    assign P[108] = in1[17] ^ in2[17];
    assign G[109] = in1[16] & in2[16];
    assign P[109] = in1[16] ^ in2[16];
    assign G[110] = in1[15] & in2[15];
    assign P[110] = in1[15] ^ in2[15];
    assign G[111] = in1[14] & in2[14];
    assign P[111] = in1[14] ^ in2[14];
    assign G[112] = in1[13] & in2[13];
    assign P[112] = in1[13] ^ in2[13];
    assign G[113] = in1[12] & in2[12];
    assign P[113] = in1[12] ^ in2[12];
    assign G[114] = in1[11] & in2[11];
    assign P[114] = in1[11] ^ in2[11];
    assign G[115] = in1[10] & in2[10];
    assign P[115] = in1[10] ^ in2[10];
    assign G[116] = in1[9] & in2[9];
    assign P[116] = in1[9] ^ in2[9];
    assign G[117] = in1[8] & in2[8];
    assign P[117] = in1[8] ^ in2[8];
    assign G[118] = in1[7] & in2[7];
    assign P[118] = in1[7] ^ in2[7];
    assign G[119] = in1[6] & in2[6];
    assign P[119] = in1[6] ^ in2[6];
    assign G[120] = in1[5] & in2[5];
    assign P[120] = in1[5] ^ in2[5];
    assign G[121] = in1[4] & in2[4];
    assign P[121] = in1[4] ^ in2[4];
    assign G[122] = in1[3] & in2[3];
    assign P[122] = in1[3] ^ in2[3];
    assign G[123] = in1[2] & in2[2];
    assign P[123] = in1[2] ^ in2[2];
    assign G[124] = in1[1] & in2[1];
    assign P[124] = in1[1] ^ in2[1];
    assign G[125] = in1[0] & in2[0];
    assign P[125] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign cout = G[125] | (P[125] & C[125]);
    assign sum = P ^ C;
endmodule

