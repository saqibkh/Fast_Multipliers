module reduced_multiplier_8(output wire [15:0] product,
                            input wire [7:0] A, B);

    assign product[0]  = 
    assign product[1]  =
    assign product[2]  =
    assign product[3]  =
    assign product[4]  =
    assign product[5]  =
    assign product[6]  =
    assign product[7]  =
    assign product[8]  =
    assign product[9]  =
    assign product[10] =
    assign product[11] =
    assign product[12] =
    assign product[13] =
    assign product[14] =
    assign product[15] =

endmodule
