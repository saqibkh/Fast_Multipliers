module multiplier_8bits_version14(product, A, B);

    output [15:0] product;
    input [7:0] A, B;

    /*
     * Area: 1192.491263
     * Power: 0.5894mW
     * Timing: 1.17ns
     */

    wire [7:0] pp0;
    wire [7:0] pp1;
    wire [7:0] pp2;
    wire [7:0] pp3;
    wire [7:0] pp4;
    wire [7:0] pp5;
    wire [7:0] pp6;
    wire [7:0] pp7;


    assign pp0 = A[0] ? B: 8'b00000000;
    assign pp1 = A[1] ? B: 8'b00000000;
    assign pp2 = A[2] ? B: 8'b00000000;
    assign pp3 = A[3] ? B: 8'b00000000;
    assign pp4 = A[4] ? B: 8'b00000000;
    assign pp5 = A[5] ? B: 8'b00000000;
    assign pp6 = A[6] ? B: 8'b00000000;
    assign pp7 = A[7] ? B: 8'b00000000;


    /*Stage 1*/
    wire[0:0] s1, in1_1, in1_2;
    wire c1;
    assign in1_1 = {pp0[6]};
    assign in1_2 = {pp1[5]};
    Half_Adder HA_1(s1, c1, in1_1, in1_2);
    wire[0:0] s2, in2_1, in2_2;
    wire c2;
    assign in2_1 = {pp0[7]};
    assign in2_2 = {pp1[6]};
    Half_Adder HA_2(s2, c2, in2_1, in2_2);
    wire[0:0] s3, in3_1, in3_2;
    wire c3;
    assign in3_1 = {pp3[4]};
    assign in3_2 = {pp4[3]};
    Full_Adder FA_3(s3, c3, in3_1, in3_2, pp2[5]);
    wire[0:0] s4, in4_1, in4_2;
    wire c4;
    assign in4_1 = {pp1[7]};
    assign in4_2 = {pp2[6]};
    Half_Adder HA_4(s4, c4, in4_1, in4_2);
    wire[0:0] s5, in5_1, in5_2;
    wire c5;
    assign in5_1 = {pp4[4]};
    assign in5_2 = {pp5[3]};
    Full_Adder FA_5(s5, c5, in5_1, in5_2, pp3[5]);
    wire[0:0] s6, in6_1, in6_2;
    wire c6;
    assign in6_1 = {pp3[6]};
    assign in6_2 = {pp4[5]};
    Full_Adder FA_6(s6, c6, in6_1, in6_2, pp2[7]);

    /*Stage 2*/
    wire[0:0] s7, in7_1, in7_2;
    wire c7;
    assign in7_1 = {pp0[4]};
    assign in7_2 = {pp1[3]};
    Half_Adder HA_7(s7, c7, in7_1, in7_2);
    wire[0:0] s8, in8_1, in8_2;
    wire c8;
    assign in8_1 = {pp0[5]};
    assign in8_2 = {pp1[4]};
    Half_Adder HA_8(s8, c8, in8_1, in8_2);
    wire[0:0] s9, in9_1, in9_2;
    wire c9;
    assign in9_1 = {pp3[2]};
    assign in9_2 = {pp4[1]};
    Full_Adder FA_9(s9, c9, in9_1, in9_2, pp2[3]);
    wire[0:0] s10, in10_1, in10_2;
    wire c10;
    assign in10_1 = {pp2[4]};
    assign in10_2 = {pp3[3]};
    Half_Adder HA_10(s10, c10, in10_1, in10_2);
    wire[0:0] s11, in11_1, in11_2;
    wire c11;
    assign in11_1 = {pp4[2]};
    assign in11_2 = {pp5[1]};
    Half_Adder HA_11(s11, c11, in11_1, in11_2);
    wire[0:0] s12, in12_1, in12_2;
    wire c12;
    assign in12_1 = {s1[0]};
    assign in12_2 = {c8};
    Full_Adder FA_12(s12, c12, in12_1, in12_2, pp6[0]);
    wire[0:0] s13, in13_1, in13_2;
    wire c13;
    assign in13_1 = {pp5[2]};
    assign in13_2 = {pp6[1]};
    Half_Adder HA_13(s13, c13, in13_1, in13_2);
    wire[0:0] s14, in14_1, in14_2;
    wire c14;
    assign in14_1 = {pp7[0]};
    assign in14_2 = {c1};
    Half_Adder HA_14(s14, c14, in14_1, in14_2);
    wire[0:0] s15, in15_1, in15_2;
    wire c15;
    assign in15_1 = {s2[0]};
    assign in15_2 = {s3[0]};
    Half_Adder HA_15(s15, c15, in15_1, in15_2);
    wire[0:0] s16, in16_1, in16_2;
    wire c16;
    assign in16_1 = {c11};
    assign in16_2 = {c12};
    Full_Adder FA_16(s16, c16, in16_1, in16_2, c10);
    wire[0:0] s17, in17_1, in17_2;
    wire c17;
    assign in17_1 = {pp6[2]};
    assign in17_2 = {pp7[1]};
    Half_Adder HA_17(s17, c17, in17_1, in17_2);
    wire[0:0] s18, in18_1, in18_2;
    wire c18;
    assign in18_1 = {c2};
    assign in18_2 = {c3};
    Half_Adder HA_18(s18, c18, in18_1, in18_2);
    wire[0:0] s19, in19_1, in19_2;
    wire c19;
    assign in19_1 = {s4[0]};
    assign in19_2 = {s5[0]};
    Half_Adder HA_19(s19, c19, in19_1, in19_2);
    wire[0:0] s20, in20_1, in20_2;
    wire c20;
    assign in20_1 = {c13};
    assign in20_2 = {c14};
    Half_Adder HA_20(s20, c20, in20_1, in20_2);
    wire[0:0] s21, in21_1, in21_2;
    wire c21;
    assign in21_1 = {c16};
    assign in21_2 = {s17[0]};
    Full_Adder FA_21(s21, c21, in21_1, in21_2, c15);
    wire[0:0] s22, in22_1, in22_2;
    wire c22;
    assign in22_1 = {pp5[4]};
    assign in22_2 = {pp6[3]};
    Half_Adder HA_22(s22, c22, in22_1, in22_2);
    wire[0:0] s23, in23_1, in23_2;
    wire c23;
    assign in23_1 = {pp7[2]};
    assign in23_2 = {c4};
    Half_Adder HA_23(s23, c23, in23_1, in23_2);
    wire[0:0] s24, in24_1, in24_2;
    wire c24;
    assign in24_1 = {c5};
    assign in24_2 = {s6[0]};
    Half_Adder HA_24(s24, c24, in24_1, in24_2);
    wire[0:0] s25, in25_1, in25_2;
    wire c25;
    assign in25_1 = {c17};
    assign in25_2 = {c18};
    Half_Adder HA_25(s25, c25, in25_1, in25_2);
    wire[0:0] s26, in26_1, in26_2;
    wire c26;
    assign in26_1 = {c19};
    assign in26_2 = {c20};
    Half_Adder HA_26(s26, c26, in26_1, in26_2);
    wire[0:0] s27, in27_1, in27_2;
    wire c27;
    assign in27_1 = {s22[0]};
    assign in27_2 = {s23[0]};
    Full_Adder FA_27(s27, c27, in27_1, in27_2, c21);
    wire[0:0] s28, in28_1, in28_2;
    wire c28;
    assign in28_1 = {pp3[7]};
    assign in28_2 = {pp4[6]};
    Half_Adder HA_28(s28, c28, in28_1, in28_2);
    wire[0:0] s29, in29_1, in29_2;
    wire c29;
    assign in29_1 = {pp5[5]};
    assign in29_2 = {pp6[4]};
    Half_Adder HA_29(s29, c29, in29_1, in29_2);
    wire[0:0] s30, in30_1, in30_2;
    wire c30;
    assign in30_1 = {pp7[3]};
    assign in30_2 = {c6};
    Half_Adder HA_30(s30, c30, in30_1, in30_2);
    wire[0:0] s31, in31_1, in31_2;
    wire c31;
    assign in31_1 = {c22};
    assign in31_2 = {c23};
    Half_Adder HA_31(s31, c31, in31_1, in31_2);
    wire[0:0] s32, in32_1, in32_2;
    wire c32;
    assign in32_1 = {c24};
    assign in32_2 = {c25};
    Half_Adder HA_32(s32, c32, in32_1, in32_2);
    wire[0:0] s33, in33_1, in33_2;
    wire c33;
    assign in33_1 = {c26};
    assign in33_2 = {c27};
    Half_Adder HA_33(s33, c33, in33_1, in33_2);
    wire[0:0] s34, in34_1, in34_2;
    wire c34;
    assign in34_1 = {s29[0]};
    assign in34_2 = {s30[0]};
    Full_Adder FA_34(s34, c34, in34_1, in34_2, s28[0]);
    wire[0:0] s35, in35_1, in35_2;
    wire c35;
    assign in35_1 = {pp4[7]};
    assign in35_2 = {pp5[6]};
    Half_Adder HA_35(s35, c35, in35_1, in35_2);
    wire[0:0] s36, in36_1, in36_2;
    wire c36;
    assign in36_1 = {pp6[5]};
    assign in36_2 = {pp7[4]};
    Half_Adder HA_36(s36, c36, in36_1, in36_2);
    wire[0:0] s37, in37_1, in37_2;
    wire c37;
    assign in37_1 = {c28};
    assign in37_2 = {c29};
    Half_Adder HA_37(s37, c37, in37_1, in37_2);
    wire[0:0] s38, in38_1, in38_2;
    wire c38;
    assign in38_1 = {c30};
    assign in38_2 = {c31};
    Half_Adder HA_38(s38, c38, in38_1, in38_2);
    wire[0:0] s39, in39_1, in39_2;
    wire c39;
    assign in39_1 = {c32};
    assign in39_2 = {c33};
    Half_Adder HA_39(s39, c39, in39_1, in39_2);
    wire[0:0] s40, in40_1, in40_2;
    wire c40;
    assign in40_1 = {s35[0]};
    assign in40_2 = {s36[0]};
    Full_Adder FA_40(s40, c40, in40_1, in40_2, c34);
    wire[0:0] s41, in41_1, in41_2;
    wire c41;
    assign in41_1 = {pp5[7]};
    assign in41_2 = {pp6[6]};
    Half_Adder HA_41(s41, c41, in41_1, in41_2);
    wire[0:0] s42, in42_1, in42_2;
    wire c42;
    assign in42_1 = {pp7[5]};
    assign in42_2 = {c35};
    Half_Adder HA_42(s42, c42, in42_1, in42_2);
    wire[0:0] s43, in43_1, in43_2;
    wire c43;
    assign in43_1 = {c36};
    assign in43_2 = {c37};
    Half_Adder HA_43(s43, c43, in43_1, in43_2);
    wire[0:0] s44, in44_1, in44_2;
    wire c44;
    assign in44_1 = {c39};
    assign in44_2 = {c40};
    Full_Adder FA_44(s44, c44, in44_1, in44_2, c38);
    wire[0:0] s45, in45_1, in45_2;
    wire c45;
    assign in45_1 = {pp7[6]};
    assign in45_2 = {c41};
    Full_Adder FA_45(s45, c45, in45_1, in45_2, pp6[7]);

    /*Stage 3*/
    wire[0:0] s46, in46_1, in46_2;
    wire c46;
    assign in46_1 = {pp0[3]};
    assign in46_2 = {pp1[2]};
    Half_Adder HA_46(s46, c46, in46_1, in46_2);
    wire[0:0] s47, in47_1, in47_2;
    wire c47;
    assign in47_1 = {pp3[1]};
    assign in47_2 = {pp4[0]};
    Full_Adder FA_47(s47, c47, in47_1, in47_2, pp2[2]);
    wire[0:0] s48, in48_1, in48_2;
    wire c48;
    assign in48_1 = {c7};
    assign in48_2 = {s8[0]};
    Full_Adder FA_48(s48, c48, in48_1, in48_2, pp5[0]);
    wire[0:0] s49, in49_1, in49_2;
    wire c49;
    assign in49_1 = {s10[0]};
    assign in49_2 = {s11[0]};
    Full_Adder FA_49(s49, c49, in49_1, in49_2, c9);
    wire[0:0] s50, in50_1, in50_2;
    wire c50;
    assign in50_1 = {s14[0]};
    assign in50_2 = {s15[0]};
    Full_Adder FA_50(s50, c50, in50_1, in50_2, s13[0]);
    wire[0:0] s51, in51_1, in51_2;
    wire c51;
    assign in51_1 = {s19[0]};
    assign in51_2 = {s20[0]};
    Full_Adder FA_51(s51, c51, in51_1, in51_2, s18[0]);
    wire[0:0] s52, in52_1, in52_2;
    wire c52;
    assign in52_1 = {s25[0]};
    assign in52_2 = {s26[0]};
    Full_Adder FA_52(s52, c52, in52_1, in52_2, s24[0]);
    wire[0:0] s53, in53_1, in53_2;
    wire c53;
    assign in53_1 = {s32[0]};
    assign in53_2 = {s33[0]};
    Full_Adder FA_53(s53, c53, in53_1, in53_2, s31[0]);
    wire[0:0] s54, in54_1, in54_2;
    wire c54;
    assign in54_1 = {s38[0]};
    assign in54_2 = {s39[0]};
    Full_Adder FA_54(s54, c54, in54_1, in54_2, s37[0]);
    wire[0:0] s55, in55_1, in55_2;
    wire c55;
    assign in55_1 = {s42[0]};
    assign in55_2 = {s43[0]};
    Full_Adder FA_55(s55, c55, in55_1, in55_2, s41[0]);
    wire[0:0] s56, in56_1, in56_2;
    wire c56;
    assign in56_1 = {c43};
    assign in56_2 = {c44};
    Full_Adder FA_56(s56, c56, in56_1, in56_2, c42);

    /*Stage 4*/
    wire[0:0] s57, in57_1, in57_2;
    wire c57;
    assign in57_1 = {pp0[2]};
    assign in57_2 = {pp1[1]};
    Half_Adder HA_57(s57, c57, in57_1, in57_2);
    wire[0:0] s58, in58_1, in58_2;
    wire c58;
    assign in58_1 = {pp3[0]};
    assign in58_2 = {s46[0]};
    Full_Adder FA_58(s58, c58, in58_1, in58_2, pp2[1]);
    wire[0:0] s59, in59_1, in59_2;
    wire c59;
    assign in59_1 = {c46};
    assign in59_2 = {s47[0]};
    Full_Adder FA_59(s59, c59, in59_1, in59_2, s7[0]);
    wire[0:0] s60, in60_1, in60_2;
    wire c60;
    assign in60_1 = {c47};
    assign in60_2 = {s48[0]};
    Full_Adder FA_60(s60, c60, in60_1, in60_2, s9[0]);
    wire[0:0] s61, in61_1, in61_2;
    wire c61;
    assign in61_1 = {c48};
    assign in61_2 = {s49[0]};
    Full_Adder FA_61(s61, c61, in61_1, in61_2, s12[0]);
    wire[0:0] s62, in62_1, in62_2;
    wire c62;
    assign in62_1 = {c49};
    assign in62_2 = {s50[0]};
    Full_Adder FA_62(s62, c62, in62_1, in62_2, s16[0]);
    wire[0:0] s63, in63_1, in63_2;
    wire c63;
    assign in63_1 = {c50};
    assign in63_2 = {s51[0]};
    Full_Adder FA_63(s63, c63, in63_1, in63_2, s21[0]);
    wire[0:0] s64, in64_1, in64_2;
    wire c64;
    assign in64_1 = {c51};
    assign in64_2 = {s52[0]};
    Full_Adder FA_64(s64, c64, in64_1, in64_2, s27[0]);
    wire[0:0] s65, in65_1, in65_2;
    wire c65;
    assign in65_1 = {c52};
    assign in65_2 = {s53[0]};
    Full_Adder FA_65(s65, c65, in65_1, in65_2, s34[0]);
    wire[0:0] s66, in66_1, in66_2;
    wire c66;
    assign in66_1 = {c53};
    assign in66_2 = {s54[0]};
    Full_Adder FA_66(s66, c66, in66_1, in66_2, s40[0]);
    wire[0:0] s67, in67_1, in67_2;
    wire c67;
    assign in67_1 = {c54};
    assign in67_2 = {s55[0]};
    Full_Adder FA_67(s67, c67, in67_1, in67_2, s44[0]);
    wire[0:0] s68, in68_1, in68_2;
    wire c68;
    assign in68_1 = {c55};
    assign in68_2 = {s56[0]};
    Full_Adder FA_68(s68, c68, in68_1, in68_2, s45[0]);


    /*Final Stage 4*/
    wire[13:0] s, in_1, in_2;
    wire c;
    assign in_1 = {pp0[1],pp2[0],c57,c58,c59,c60,c61,c62,c63,c64,c65,c66,c67,c68};
    assign in_2 = {pp1[0],s57[0],s58[0],s59[0],s60[0],s61[0],s62[0],s63[0],s64[0],s65[0],s66[0],s67[0],s68[0],1'b0};
    CLA_14(s, c, in_1, in_2);

    assign product[0] = pp0[0];
    assign product[1] = s[0];
    assign product[2] = s[1];
    assign product[3] = s[2];
    assign product[4] = s[3];
    assign product[5] = s[4];
    assign product[6] = s[5];
    assign product[7] = s[6];
    assign product[8] = s[7];
    assign product[9] = s[8];
    assign product[10] = s[9];
    assign product[11] = s[10];
    assign product[12] = s[11];
    assign product[13] = s[12];
    assign product[14] = s[13];
    assign product[15] = c;
endmodule


module CLA_14(output [13:0] sum, output cout, input [13:0] in1, input [13:0] in2);

    wire[13:0] G;
    wire[13:0] C;
    wire[13:0] P;

    assign G[0] = in1[13] & in2[13];
    assign P[0] = in1[13] ^ in2[13];
    assign G[1] = in1[12] & in2[12];
    assign P[1] = in1[12] ^ in2[12];
    assign G[2] = in1[11] & in2[11];
    assign P[2] = in1[11] ^ in2[11];
    assign G[3] = in1[10] & in2[10];
    assign P[3] = in1[10] ^ in2[10];
    assign G[4] = in1[9] & in2[9];
    assign P[4] = in1[9] ^ in2[9];
    assign G[5] = in1[8] & in2[8];
    assign P[5] = in1[8] ^ in2[8];
    assign G[6] = in1[7] & in2[7];
    assign P[6] = in1[7] ^ in2[7];
    assign G[7] = in1[6] & in2[6];
    assign P[7] = in1[6] ^ in2[6];
    assign G[8] = in1[5] & in2[5];
    assign P[8] = in1[5] ^ in2[5];
    assign G[9] = in1[4] & in2[4];
    assign P[9] = in1[4] ^ in2[4];
    assign G[10] = in1[3] & in2[3];
    assign P[10] = in1[3] ^ in2[3];
    assign G[11] = in1[2] & in2[2];
    assign P[11] = in1[2] ^ in2[2];
    assign G[12] = in1[1] & in2[1];
    assign P[12] = in1[1] ^ in2[1];
    assign G[13] = in1[0] & in2[0];
    assign P[13] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign cout = G[13] | (P[13] & C[13]);
    assign sum = P ^ C;
endmodule

module Half_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2);
    xor(sum, in1, in2);
    and(cout, in1, in2);
endmodule

module Full_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2,
                  input wire cin);
    wire temp1;
    wire temp2;
    wire temp3;
    xor(sum, in1, in2, cin);
    and(temp1,in1,in2);
    and(temp2,in1,cin);
    and(temp3,in2,cin);
    or(cout,temp1,temp2,temp3);
endmodule
