module kogge_stone_64(output [63:0] sum,
        output cout,
        input [63:0] in1,
        input [63:0] in2);

    /* 
     * Area: 3520.688503
     * Power: 1.1894mW
     * Timing: 0.68ns
     */

    assign cin = 0;
    wire[63:0] G_0;
    wire[63:0] P_0;
    wire[63:0] G_1;
    wire[63:0] P_1;
    wire[63:0] G_2;
    wire[63:0] P_2;
    wire[63:0] G_3;
    wire[63:0] P_3;
    wire[63:0] G_4;
    wire[63:0] P_4;
    wire[63:0] G_5;
    wire[63:0] P_5;
    wire[63:0] G_6;
    wire[63:0] P_6;
    wire[63:0] G_7;
    wire[63:0] P_7;

    assign G_0[0] = in1[63] & in2[63];
    assign P_0[0] = in1[63] ^ in2[63];
    assign G_0[1] = in1[62] & in2[62];
    assign P_0[1] = in1[62] ^ in2[62];
    assign G_0[2] = in1[61] & in2[61];
    assign P_0[2] = in1[61] ^ in2[61];
    assign G_0[3] = in1[60] & in2[60];
    assign P_0[3] = in1[60] ^ in2[60];
    assign G_0[4] = in1[59] & in2[59];
    assign P_0[4] = in1[59] ^ in2[59];
    assign G_0[5] = in1[58] & in2[58];
    assign P_0[5] = in1[58] ^ in2[58];
    assign G_0[6] = in1[57] & in2[57];
    assign P_0[6] = in1[57] ^ in2[57];
    assign G_0[7] = in1[56] & in2[56];
    assign P_0[7] = in1[56] ^ in2[56];
    assign G_0[8] = in1[55] & in2[55];
    assign P_0[8] = in1[55] ^ in2[55];
    assign G_0[9] = in1[54] & in2[54];
    assign P_0[9] = in1[54] ^ in2[54];
    assign G_0[10] = in1[53] & in2[53];
    assign P_0[10] = in1[53] ^ in2[53];
    assign G_0[11] = in1[52] & in2[52];
    assign P_0[11] = in1[52] ^ in2[52];
    assign G_0[12] = in1[51] & in2[51];
    assign P_0[12] = in1[51] ^ in2[51];
    assign G_0[13] = in1[50] & in2[50];
    assign P_0[13] = in1[50] ^ in2[50];
    assign G_0[14] = in1[49] & in2[49];
    assign P_0[14] = in1[49] ^ in2[49];
    assign G_0[15] = in1[48] & in2[48];
    assign P_0[15] = in1[48] ^ in2[48];
    assign G_0[16] = in1[47] & in2[47];
    assign P_0[16] = in1[47] ^ in2[47];
    assign G_0[17] = in1[46] & in2[46];
    assign P_0[17] = in1[46] ^ in2[46];
    assign G_0[18] = in1[45] & in2[45];
    assign P_0[18] = in1[45] ^ in2[45];
    assign G_0[19] = in1[44] & in2[44];
    assign P_0[19] = in1[44] ^ in2[44];
    assign G_0[20] = in1[43] & in2[43];
    assign P_0[20] = in1[43] ^ in2[43];
    assign G_0[21] = in1[42] & in2[42];
    assign P_0[21] = in1[42] ^ in2[42];
    assign G_0[22] = in1[41] & in2[41];
    assign P_0[22] = in1[41] ^ in2[41];
    assign G_0[23] = in1[40] & in2[40];
    assign P_0[23] = in1[40] ^ in2[40];
    assign G_0[24] = in1[39] & in2[39];
    assign P_0[24] = in1[39] ^ in2[39];
    assign G_0[25] = in1[38] & in2[38];
    assign P_0[25] = in1[38] ^ in2[38];
    assign G_0[26] = in1[37] & in2[37];
    assign P_0[26] = in1[37] ^ in2[37];
    assign G_0[27] = in1[36] & in2[36];
    assign P_0[27] = in1[36] ^ in2[36];
    assign G_0[28] = in1[35] & in2[35];
    assign P_0[28] = in1[35] ^ in2[35];
    assign G_0[29] = in1[34] & in2[34];
    assign P_0[29] = in1[34] ^ in2[34];
    assign G_0[30] = in1[33] & in2[33];
    assign P_0[30] = in1[33] ^ in2[33];
    assign G_0[31] = in1[32] & in2[32];
    assign P_0[31] = in1[32] ^ in2[32];
    assign G_0[32] = in1[31] & in2[31];
    assign P_0[32] = in1[31] ^ in2[31];
    assign G_0[33] = in1[30] & in2[30];
    assign P_0[33] = in1[30] ^ in2[30];
    assign G_0[34] = in1[29] & in2[29];
    assign P_0[34] = in1[29] ^ in2[29];
    assign G_0[35] = in1[28] & in2[28];
    assign P_0[35] = in1[28] ^ in2[28];
    assign G_0[36] = in1[27] & in2[27];
    assign P_0[36] = in1[27] ^ in2[27];
    assign G_0[37] = in1[26] & in2[26];
    assign P_0[37] = in1[26] ^ in2[26];
    assign G_0[38] = in1[25] & in2[25];
    assign P_0[38] = in1[25] ^ in2[25];
    assign G_0[39] = in1[24] & in2[24];
    assign P_0[39] = in1[24] ^ in2[24];
    assign G_0[40] = in1[23] & in2[23];
    assign P_0[40] = in1[23] ^ in2[23];
    assign G_0[41] = in1[22] & in2[22];
    assign P_0[41] = in1[22] ^ in2[22];
    assign G_0[42] = in1[21] & in2[21];
    assign P_0[42] = in1[21] ^ in2[21];
    assign G_0[43] = in1[20] & in2[20];
    assign P_0[43] = in1[20] ^ in2[20];
    assign G_0[44] = in1[19] & in2[19];
    assign P_0[44] = in1[19] ^ in2[19];
    assign G_0[45] = in1[18] & in2[18];
    assign P_0[45] = in1[18] ^ in2[18];
    assign G_0[46] = in1[17] & in2[17];
    assign P_0[46] = in1[17] ^ in2[17];
    assign G_0[47] = in1[16] & in2[16];
    assign P_0[47] = in1[16] ^ in2[16];
    assign G_0[48] = in1[15] & in2[15];
    assign P_0[48] = in1[15] ^ in2[15];
    assign G_0[49] = in1[14] & in2[14];
    assign P_0[49] = in1[14] ^ in2[14];
    assign G_0[50] = in1[13] & in2[13];
    assign P_0[50] = in1[13] ^ in2[13];
    assign G_0[51] = in1[12] & in2[12];
    assign P_0[51] = in1[12] ^ in2[12];
    assign G_0[52] = in1[11] & in2[11];
    assign P_0[52] = in1[11] ^ in2[11];
    assign G_0[53] = in1[10] & in2[10];
    assign P_0[53] = in1[10] ^ in2[10];
    assign G_0[54] = in1[9] & in2[9];
    assign P_0[54] = in1[9] ^ in2[9];
    assign G_0[55] = in1[8] & in2[8];
    assign P_0[55] = in1[8] ^ in2[8];
    assign G_0[56] = in1[7] & in2[7];
    assign P_0[56] = in1[7] ^ in2[7];
    assign G_0[57] = in1[6] & in2[6];
    assign P_0[57] = in1[6] ^ in2[6];
    assign G_0[58] = in1[5] & in2[5];
    assign P_0[58] = in1[5] ^ in2[5];
    assign G_0[59] = in1[4] & in2[4];
    assign P_0[59] = in1[4] ^ in2[4];
    assign G_0[60] = in1[3] & in2[3];
    assign P_0[60] = in1[3] ^ in2[3];
    assign G_0[61] = in1[2] & in2[2];
    assign P_0[61] = in1[2] ^ in2[2];
    assign G_0[62] = in1[1] & in2[1];
    assign P_0[62] = in1[1] ^ in2[1];
    assign G_0[63] = in1[0] & in2[0];
    assign P_0[63] = in1[0] ^ in2[0];



    /*Stage 1*/
    gray_cell level_1_0(cin, P_0[0], G_0[0], G_1[0]);
    black_cell level_0_1(G_0[0], P_0[1], G_0[1], P_0[0], G_1[1], P_1[1]);
    black_cell level_0_2(G_0[1], P_0[2], G_0[2], P_0[1], G_1[2], P_1[2]);
    black_cell level_0_3(G_0[2], P_0[3], G_0[3], P_0[2], G_1[3], P_1[3]);
    black_cell level_0_4(G_0[3], P_0[4], G_0[4], P_0[3], G_1[4], P_1[4]);
    black_cell level_0_5(G_0[4], P_0[5], G_0[5], P_0[4], G_1[5], P_1[5]);
    black_cell level_0_6(G_0[5], P_0[6], G_0[6], P_0[5], G_1[6], P_1[6]);
    black_cell level_0_7(G_0[6], P_0[7], G_0[7], P_0[6], G_1[7], P_1[7]);
    black_cell level_0_8(G_0[7], P_0[8], G_0[8], P_0[7], G_1[8], P_1[8]);
    black_cell level_0_9(G_0[8], P_0[9], G_0[9], P_0[8], G_1[9], P_1[9]);
    black_cell level_0_10(G_0[9], P_0[10], G_0[10], P_0[9], G_1[10], P_1[10]);
    black_cell level_0_11(G_0[10], P_0[11], G_0[11], P_0[10], G_1[11], P_1[11]);
    black_cell level_0_12(G_0[11], P_0[12], G_0[12], P_0[11], G_1[12], P_1[12]);
    black_cell level_0_13(G_0[12], P_0[13], G_0[13], P_0[12], G_1[13], P_1[13]);
    black_cell level_0_14(G_0[13], P_0[14], G_0[14], P_0[13], G_1[14], P_1[14]);
    black_cell level_0_15(G_0[14], P_0[15], G_0[15], P_0[14], G_1[15], P_1[15]);
    black_cell level_0_16(G_0[15], P_0[16], G_0[16], P_0[15], G_1[16], P_1[16]);
    black_cell level_0_17(G_0[16], P_0[17], G_0[17], P_0[16], G_1[17], P_1[17]);
    black_cell level_0_18(G_0[17], P_0[18], G_0[18], P_0[17], G_1[18], P_1[18]);
    black_cell level_0_19(G_0[18], P_0[19], G_0[19], P_0[18], G_1[19], P_1[19]);
    black_cell level_0_20(G_0[19], P_0[20], G_0[20], P_0[19], G_1[20], P_1[20]);
    black_cell level_0_21(G_0[20], P_0[21], G_0[21], P_0[20], G_1[21], P_1[21]);
    black_cell level_0_22(G_0[21], P_0[22], G_0[22], P_0[21], G_1[22], P_1[22]);
    black_cell level_0_23(G_0[22], P_0[23], G_0[23], P_0[22], G_1[23], P_1[23]);
    black_cell level_0_24(G_0[23], P_0[24], G_0[24], P_0[23], G_1[24], P_1[24]);
    black_cell level_0_25(G_0[24], P_0[25], G_0[25], P_0[24], G_1[25], P_1[25]);
    black_cell level_0_26(G_0[25], P_0[26], G_0[26], P_0[25], G_1[26], P_1[26]);
    black_cell level_0_27(G_0[26], P_0[27], G_0[27], P_0[26], G_1[27], P_1[27]);
    black_cell level_0_28(G_0[27], P_0[28], G_0[28], P_0[27], G_1[28], P_1[28]);
    black_cell level_0_29(G_0[28], P_0[29], G_0[29], P_0[28], G_1[29], P_1[29]);
    black_cell level_0_30(G_0[29], P_0[30], G_0[30], P_0[29], G_1[30], P_1[30]);
    black_cell level_0_31(G_0[30], P_0[31], G_0[31], P_0[30], G_1[31], P_1[31]);
    black_cell level_0_32(G_0[31], P_0[32], G_0[32], P_0[31], G_1[32], P_1[32]);
    black_cell level_0_33(G_0[32], P_0[33], G_0[33], P_0[32], G_1[33], P_1[33]);
    black_cell level_0_34(G_0[33], P_0[34], G_0[34], P_0[33], G_1[34], P_1[34]);
    black_cell level_0_35(G_0[34], P_0[35], G_0[35], P_0[34], G_1[35], P_1[35]);
    black_cell level_0_36(G_0[35], P_0[36], G_0[36], P_0[35], G_1[36], P_1[36]);
    black_cell level_0_37(G_0[36], P_0[37], G_0[37], P_0[36], G_1[37], P_1[37]);
    black_cell level_0_38(G_0[37], P_0[38], G_0[38], P_0[37], G_1[38], P_1[38]);
    black_cell level_0_39(G_0[38], P_0[39], G_0[39], P_0[38], G_1[39], P_1[39]);
    black_cell level_0_40(G_0[39], P_0[40], G_0[40], P_0[39], G_1[40], P_1[40]);
    black_cell level_0_41(G_0[40], P_0[41], G_0[41], P_0[40], G_1[41], P_1[41]);
    black_cell level_0_42(G_0[41], P_0[42], G_0[42], P_0[41], G_1[42], P_1[42]);
    black_cell level_0_43(G_0[42], P_0[43], G_0[43], P_0[42], G_1[43], P_1[43]);
    black_cell level_0_44(G_0[43], P_0[44], G_0[44], P_0[43], G_1[44], P_1[44]);
    black_cell level_0_45(G_0[44], P_0[45], G_0[45], P_0[44], G_1[45], P_1[45]);
    black_cell level_0_46(G_0[45], P_0[46], G_0[46], P_0[45], G_1[46], P_1[46]);
    black_cell level_0_47(G_0[46], P_0[47], G_0[47], P_0[46], G_1[47], P_1[47]);
    black_cell level_0_48(G_0[47], P_0[48], G_0[48], P_0[47], G_1[48], P_1[48]);
    black_cell level_0_49(G_0[48], P_0[49], G_0[49], P_0[48], G_1[49], P_1[49]);
    black_cell level_0_50(G_0[49], P_0[50], G_0[50], P_0[49], G_1[50], P_1[50]);
    black_cell level_0_51(G_0[50], P_0[51], G_0[51], P_0[50], G_1[51], P_1[51]);
    black_cell level_0_52(G_0[51], P_0[52], G_0[52], P_0[51], G_1[52], P_1[52]);
    black_cell level_0_53(G_0[52], P_0[53], G_0[53], P_0[52], G_1[53], P_1[53]);
    black_cell level_0_54(G_0[53], P_0[54], G_0[54], P_0[53], G_1[54], P_1[54]);
    black_cell level_0_55(G_0[54], P_0[55], G_0[55], P_0[54], G_1[55], P_1[55]);
    black_cell level_0_56(G_0[55], P_0[56], G_0[56], P_0[55], G_1[56], P_1[56]);
    black_cell level_0_57(G_0[56], P_0[57], G_0[57], P_0[56], G_1[57], P_1[57]);
    black_cell level_0_58(G_0[57], P_0[58], G_0[58], P_0[57], G_1[58], P_1[58]);
    black_cell level_0_59(G_0[58], P_0[59], G_0[59], P_0[58], G_1[59], P_1[59]);
    black_cell level_0_60(G_0[59], P_0[60], G_0[60], P_0[59], G_1[60], P_1[60]);
    black_cell level_0_61(G_0[60], P_0[61], G_0[61], P_0[60], G_1[61], P_1[61]);
    black_cell level_0_62(G_0[61], P_0[62], G_0[62], P_0[61], G_1[62], P_1[62]);
    black_cell level_0_63(G_0[62], P_0[63], G_0[63], P_0[62], G_1[63], P_1[63]);

    /*Stage 2*/
    gray_cell level_2_1(cin, P_1[1], G_1[1], G_2[1]);
    gray_cell level_2_2(G_1[0], P_1[2], G_1[2], G_2[2]);
    black_cell level_1_3(G_1[1], P_1[3], G_1[3], P_1[1], G_2[3], P_2[3]);
    black_cell level_1_4(G_1[2], P_1[4], G_1[4], P_1[2], G_2[4], P_2[4]);
    black_cell level_1_5(G_1[3], P_1[5], G_1[5], P_1[3], G_2[5], P_2[5]);
    black_cell level_1_6(G_1[4], P_1[6], G_1[6], P_1[4], G_2[6], P_2[6]);
    black_cell level_1_7(G_1[5], P_1[7], G_1[7], P_1[5], G_2[7], P_2[7]);
    black_cell level_1_8(G_1[6], P_1[8], G_1[8], P_1[6], G_2[8], P_2[8]);
    black_cell level_1_9(G_1[7], P_1[9], G_1[9], P_1[7], G_2[9], P_2[9]);
    black_cell level_1_10(G_1[8], P_1[10], G_1[10], P_1[8], G_2[10], P_2[10]);
    black_cell level_1_11(G_1[9], P_1[11], G_1[11], P_1[9], G_2[11], P_2[11]);
    black_cell level_1_12(G_1[10], P_1[12], G_1[12], P_1[10], G_2[12], P_2[12]);
    black_cell level_1_13(G_1[11], P_1[13], G_1[13], P_1[11], G_2[13], P_2[13]);
    black_cell level_1_14(G_1[12], P_1[14], G_1[14], P_1[12], G_2[14], P_2[14]);
    black_cell level_1_15(G_1[13], P_1[15], G_1[15], P_1[13], G_2[15], P_2[15]);
    black_cell level_1_16(G_1[14], P_1[16], G_1[16], P_1[14], G_2[16], P_2[16]);
    black_cell level_1_17(G_1[15], P_1[17], G_1[17], P_1[15], G_2[17], P_2[17]);
    black_cell level_1_18(G_1[16], P_1[18], G_1[18], P_1[16], G_2[18], P_2[18]);
    black_cell level_1_19(G_1[17], P_1[19], G_1[19], P_1[17], G_2[19], P_2[19]);
    black_cell level_1_20(G_1[18], P_1[20], G_1[20], P_1[18], G_2[20], P_2[20]);
    black_cell level_1_21(G_1[19], P_1[21], G_1[21], P_1[19], G_2[21], P_2[21]);
    black_cell level_1_22(G_1[20], P_1[22], G_1[22], P_1[20], G_2[22], P_2[22]);
    black_cell level_1_23(G_1[21], P_1[23], G_1[23], P_1[21], G_2[23], P_2[23]);
    black_cell level_1_24(G_1[22], P_1[24], G_1[24], P_1[22], G_2[24], P_2[24]);
    black_cell level_1_25(G_1[23], P_1[25], G_1[25], P_1[23], G_2[25], P_2[25]);
    black_cell level_1_26(G_1[24], P_1[26], G_1[26], P_1[24], G_2[26], P_2[26]);
    black_cell level_1_27(G_1[25], P_1[27], G_1[27], P_1[25], G_2[27], P_2[27]);
    black_cell level_1_28(G_1[26], P_1[28], G_1[28], P_1[26], G_2[28], P_2[28]);
    black_cell level_1_29(G_1[27], P_1[29], G_1[29], P_1[27], G_2[29], P_2[29]);
    black_cell level_1_30(G_1[28], P_1[30], G_1[30], P_1[28], G_2[30], P_2[30]);
    black_cell level_1_31(G_1[29], P_1[31], G_1[31], P_1[29], G_2[31], P_2[31]);
    black_cell level_1_32(G_1[30], P_1[32], G_1[32], P_1[30], G_2[32], P_2[32]);
    black_cell level_1_33(G_1[31], P_1[33], G_1[33], P_1[31], G_2[33], P_2[33]);
    black_cell level_1_34(G_1[32], P_1[34], G_1[34], P_1[32], G_2[34], P_2[34]);
    black_cell level_1_35(G_1[33], P_1[35], G_1[35], P_1[33], G_2[35], P_2[35]);
    black_cell level_1_36(G_1[34], P_1[36], G_1[36], P_1[34], G_2[36], P_2[36]);
    black_cell level_1_37(G_1[35], P_1[37], G_1[37], P_1[35], G_2[37], P_2[37]);
    black_cell level_1_38(G_1[36], P_1[38], G_1[38], P_1[36], G_2[38], P_2[38]);
    black_cell level_1_39(G_1[37], P_1[39], G_1[39], P_1[37], G_2[39], P_2[39]);
    black_cell level_1_40(G_1[38], P_1[40], G_1[40], P_1[38], G_2[40], P_2[40]);
    black_cell level_1_41(G_1[39], P_1[41], G_1[41], P_1[39], G_2[41], P_2[41]);
    black_cell level_1_42(G_1[40], P_1[42], G_1[42], P_1[40], G_2[42], P_2[42]);
    black_cell level_1_43(G_1[41], P_1[43], G_1[43], P_1[41], G_2[43], P_2[43]);
    black_cell level_1_44(G_1[42], P_1[44], G_1[44], P_1[42], G_2[44], P_2[44]);
    black_cell level_1_45(G_1[43], P_1[45], G_1[45], P_1[43], G_2[45], P_2[45]);
    black_cell level_1_46(G_1[44], P_1[46], G_1[46], P_1[44], G_2[46], P_2[46]);
    black_cell level_1_47(G_1[45], P_1[47], G_1[47], P_1[45], G_2[47], P_2[47]);
    black_cell level_1_48(G_1[46], P_1[48], G_1[48], P_1[46], G_2[48], P_2[48]);
    black_cell level_1_49(G_1[47], P_1[49], G_1[49], P_1[47], G_2[49], P_2[49]);
    black_cell level_1_50(G_1[48], P_1[50], G_1[50], P_1[48], G_2[50], P_2[50]);
    black_cell level_1_51(G_1[49], P_1[51], G_1[51], P_1[49], G_2[51], P_2[51]);
    black_cell level_1_52(G_1[50], P_1[52], G_1[52], P_1[50], G_2[52], P_2[52]);
    black_cell level_1_53(G_1[51], P_1[53], G_1[53], P_1[51], G_2[53], P_2[53]);
    black_cell level_1_54(G_1[52], P_1[54], G_1[54], P_1[52], G_2[54], P_2[54]);
    black_cell level_1_55(G_1[53], P_1[55], G_1[55], P_1[53], G_2[55], P_2[55]);
    black_cell level_1_56(G_1[54], P_1[56], G_1[56], P_1[54], G_2[56], P_2[56]);
    black_cell level_1_57(G_1[55], P_1[57], G_1[57], P_1[55], G_2[57], P_2[57]);
    black_cell level_1_58(G_1[56], P_1[58], G_1[58], P_1[56], G_2[58], P_2[58]);
    black_cell level_1_59(G_1[57], P_1[59], G_1[59], P_1[57], G_2[59], P_2[59]);
    black_cell level_1_60(G_1[58], P_1[60], G_1[60], P_1[58], G_2[60], P_2[60]);
    black_cell level_1_61(G_1[59], P_1[61], G_1[61], P_1[59], G_2[61], P_2[61]);
    black_cell level_1_62(G_1[60], P_1[62], G_1[62], P_1[60], G_2[62], P_2[62]);
    black_cell level_1_63(G_1[61], P_1[63], G_1[63], P_1[61], G_2[63], P_2[63]);

    /*Stage 3*/
    gray_cell level_3_3(cin, P_2[3], G_2[3], G_3[3]);
    gray_cell level_3_4(G_1[0], P_2[4], G_2[4], G_3[4]);
    gray_cell level_3_5(G_2[1], P_2[5], G_2[5], G_3[5]);
    gray_cell level_3_6(G_2[2], P_2[6], G_2[6], G_3[6]);
    black_cell level_2_7(G_2[3], P_2[7], G_2[7], P_2[3], G_3[7], P_3[7]);
    black_cell level_2_8(G_2[4], P_2[8], G_2[8], P_2[4], G_3[8], P_3[8]);
    black_cell level_2_9(G_2[5], P_2[9], G_2[9], P_2[5], G_3[9], P_3[9]);
    black_cell level_2_10(G_2[6], P_2[10], G_2[10], P_2[6], G_3[10], P_3[10]);
    black_cell level_2_11(G_2[7], P_2[11], G_2[11], P_2[7], G_3[11], P_3[11]);
    black_cell level_2_12(G_2[8], P_2[12], G_2[12], P_2[8], G_3[12], P_3[12]);
    black_cell level_2_13(G_2[9], P_2[13], G_2[13], P_2[9], G_3[13], P_3[13]);
    black_cell level_2_14(G_2[10], P_2[14], G_2[14], P_2[10], G_3[14], P_3[14]);
    black_cell level_2_15(G_2[11], P_2[15], G_2[15], P_2[11], G_3[15], P_3[15]);
    black_cell level_2_16(G_2[12], P_2[16], G_2[16], P_2[12], G_3[16], P_3[16]);
    black_cell level_2_17(G_2[13], P_2[17], G_2[17], P_2[13], G_3[17], P_3[17]);
    black_cell level_2_18(G_2[14], P_2[18], G_2[18], P_2[14], G_3[18], P_3[18]);
    black_cell level_2_19(G_2[15], P_2[19], G_2[19], P_2[15], G_3[19], P_3[19]);
    black_cell level_2_20(G_2[16], P_2[20], G_2[20], P_2[16], G_3[20], P_3[20]);
    black_cell level_2_21(G_2[17], P_2[21], G_2[21], P_2[17], G_3[21], P_3[21]);
    black_cell level_2_22(G_2[18], P_2[22], G_2[22], P_2[18], G_3[22], P_3[22]);
    black_cell level_2_23(G_2[19], P_2[23], G_2[23], P_2[19], G_3[23], P_3[23]);
    black_cell level_2_24(G_2[20], P_2[24], G_2[24], P_2[20], G_3[24], P_3[24]);
    black_cell level_2_25(G_2[21], P_2[25], G_2[25], P_2[21], G_3[25], P_3[25]);
    black_cell level_2_26(G_2[22], P_2[26], G_2[26], P_2[22], G_3[26], P_3[26]);
    black_cell level_2_27(G_2[23], P_2[27], G_2[27], P_2[23], G_3[27], P_3[27]);
    black_cell level_2_28(G_2[24], P_2[28], G_2[28], P_2[24], G_3[28], P_3[28]);
    black_cell level_2_29(G_2[25], P_2[29], G_2[29], P_2[25], G_3[29], P_3[29]);
    black_cell level_2_30(G_2[26], P_2[30], G_2[30], P_2[26], G_3[30], P_3[30]);
    black_cell level_2_31(G_2[27], P_2[31], G_2[31], P_2[27], G_3[31], P_3[31]);
    black_cell level_2_32(G_2[28], P_2[32], G_2[32], P_2[28], G_3[32], P_3[32]);
    black_cell level_2_33(G_2[29], P_2[33], G_2[33], P_2[29], G_3[33], P_3[33]);
    black_cell level_2_34(G_2[30], P_2[34], G_2[34], P_2[30], G_3[34], P_3[34]);
    black_cell level_2_35(G_2[31], P_2[35], G_2[35], P_2[31], G_3[35], P_3[35]);
    black_cell level_2_36(G_2[32], P_2[36], G_2[36], P_2[32], G_3[36], P_3[36]);
    black_cell level_2_37(G_2[33], P_2[37], G_2[37], P_2[33], G_3[37], P_3[37]);
    black_cell level_2_38(G_2[34], P_2[38], G_2[38], P_2[34], G_3[38], P_3[38]);
    black_cell level_2_39(G_2[35], P_2[39], G_2[39], P_2[35], G_3[39], P_3[39]);
    black_cell level_2_40(G_2[36], P_2[40], G_2[40], P_2[36], G_3[40], P_3[40]);
    black_cell level_2_41(G_2[37], P_2[41], G_2[41], P_2[37], G_3[41], P_3[41]);
    black_cell level_2_42(G_2[38], P_2[42], G_2[42], P_2[38], G_3[42], P_3[42]);
    black_cell level_2_43(G_2[39], P_2[43], G_2[43], P_2[39], G_3[43], P_3[43]);
    black_cell level_2_44(G_2[40], P_2[44], G_2[44], P_2[40], G_3[44], P_3[44]);
    black_cell level_2_45(G_2[41], P_2[45], G_2[45], P_2[41], G_3[45], P_3[45]);
    black_cell level_2_46(G_2[42], P_2[46], G_2[46], P_2[42], G_3[46], P_3[46]);
    black_cell level_2_47(G_2[43], P_2[47], G_2[47], P_2[43], G_3[47], P_3[47]);
    black_cell level_2_48(G_2[44], P_2[48], G_2[48], P_2[44], G_3[48], P_3[48]);
    black_cell level_2_49(G_2[45], P_2[49], G_2[49], P_2[45], G_3[49], P_3[49]);
    black_cell level_2_50(G_2[46], P_2[50], G_2[50], P_2[46], G_3[50], P_3[50]);
    black_cell level_2_51(G_2[47], P_2[51], G_2[51], P_2[47], G_3[51], P_3[51]);
    black_cell level_2_52(G_2[48], P_2[52], G_2[52], P_2[48], G_3[52], P_3[52]);
    black_cell level_2_53(G_2[49], P_2[53], G_2[53], P_2[49], G_3[53], P_3[53]);
    black_cell level_2_54(G_2[50], P_2[54], G_2[54], P_2[50], G_3[54], P_3[54]);
    black_cell level_2_55(G_2[51], P_2[55], G_2[55], P_2[51], G_3[55], P_3[55]);
    black_cell level_2_56(G_2[52], P_2[56], G_2[56], P_2[52], G_3[56], P_3[56]);
    black_cell level_2_57(G_2[53], P_2[57], G_2[57], P_2[53], G_3[57], P_3[57]);
    black_cell level_2_58(G_2[54], P_2[58], G_2[58], P_2[54], G_3[58], P_3[58]);
    black_cell level_2_59(G_2[55], P_2[59], G_2[59], P_2[55], G_3[59], P_3[59]);
    black_cell level_2_60(G_2[56], P_2[60], G_2[60], P_2[56], G_3[60], P_3[60]);
    black_cell level_2_61(G_2[57], P_2[61], G_2[61], P_2[57], G_3[61], P_3[61]);
    black_cell level_2_62(G_2[58], P_2[62], G_2[62], P_2[58], G_3[62], P_3[62]);
    black_cell level_2_63(G_2[59], P_2[63], G_2[63], P_2[59], G_3[63], P_3[63]);

    /*Stage 4*/
    gray_cell level_4_7(cin, P_3[7], G_3[7], G_4[7]);
    gray_cell level_4_8(G_1[0], P_3[8], G_3[8], G_4[8]);
    gray_cell level_4_9(G_2[1], P_3[9], G_3[9], G_4[9]);
    gray_cell level_4_10(G_2[2], P_3[10], G_3[10], G_4[10]);
    gray_cell level_4_11(G_3[3], P_3[11], G_3[11], G_4[11]);
    gray_cell level_4_12(G_3[4], P_3[12], G_3[12], G_4[12]);
    gray_cell level_4_13(G_3[5], P_3[13], G_3[13], G_4[13]);
    gray_cell level_4_14(G_3[6], P_3[14], G_3[14], G_4[14]);
    black_cell level_3_15(G_3[7], P_3[15], G_3[15], P_3[7], G_4[15], P_4[15]);
    black_cell level_3_16(G_3[8], P_3[16], G_3[16], P_3[8], G_4[16], P_4[16]);
    black_cell level_3_17(G_3[9], P_3[17], G_3[17], P_3[9], G_4[17], P_4[17]);
    black_cell level_3_18(G_3[10], P_3[18], G_3[18], P_3[10], G_4[18], P_4[18]);
    black_cell level_3_19(G_3[11], P_3[19], G_3[19], P_3[11], G_4[19], P_4[19]);
    black_cell level_3_20(G_3[12], P_3[20], G_3[20], P_3[12], G_4[20], P_4[20]);
    black_cell level_3_21(G_3[13], P_3[21], G_3[21], P_3[13], G_4[21], P_4[21]);
    black_cell level_3_22(G_3[14], P_3[22], G_3[22], P_3[14], G_4[22], P_4[22]);
    black_cell level_3_23(G_3[15], P_3[23], G_3[23], P_3[15], G_4[23], P_4[23]);
    black_cell level_3_24(G_3[16], P_3[24], G_3[24], P_3[16], G_4[24], P_4[24]);
    black_cell level_3_25(G_3[17], P_3[25], G_3[25], P_3[17], G_4[25], P_4[25]);
    black_cell level_3_26(G_3[18], P_3[26], G_3[26], P_3[18], G_4[26], P_4[26]);
    black_cell level_3_27(G_3[19], P_3[27], G_3[27], P_3[19], G_4[27], P_4[27]);
    black_cell level_3_28(G_3[20], P_3[28], G_3[28], P_3[20], G_4[28], P_4[28]);
    black_cell level_3_29(G_3[21], P_3[29], G_3[29], P_3[21], G_4[29], P_4[29]);
    black_cell level_3_30(G_3[22], P_3[30], G_3[30], P_3[22], G_4[30], P_4[30]);
    black_cell level_3_31(G_3[23], P_3[31], G_3[31], P_3[23], G_4[31], P_4[31]);
    black_cell level_3_32(G_3[24], P_3[32], G_3[32], P_3[24], G_4[32], P_4[32]);
    black_cell level_3_33(G_3[25], P_3[33], G_3[33], P_3[25], G_4[33], P_4[33]);
    black_cell level_3_34(G_3[26], P_3[34], G_3[34], P_3[26], G_4[34], P_4[34]);
    black_cell level_3_35(G_3[27], P_3[35], G_3[35], P_3[27], G_4[35], P_4[35]);
    black_cell level_3_36(G_3[28], P_3[36], G_3[36], P_3[28], G_4[36], P_4[36]);
    black_cell level_3_37(G_3[29], P_3[37], G_3[37], P_3[29], G_4[37], P_4[37]);
    black_cell level_3_38(G_3[30], P_3[38], G_3[38], P_3[30], G_4[38], P_4[38]);
    black_cell level_3_39(G_3[31], P_3[39], G_3[39], P_3[31], G_4[39], P_4[39]);
    black_cell level_3_40(G_3[32], P_3[40], G_3[40], P_3[32], G_4[40], P_4[40]);
    black_cell level_3_41(G_3[33], P_3[41], G_3[41], P_3[33], G_4[41], P_4[41]);
    black_cell level_3_42(G_3[34], P_3[42], G_3[42], P_3[34], G_4[42], P_4[42]);
    black_cell level_3_43(G_3[35], P_3[43], G_3[43], P_3[35], G_4[43], P_4[43]);
    black_cell level_3_44(G_3[36], P_3[44], G_3[44], P_3[36], G_4[44], P_4[44]);
    black_cell level_3_45(G_3[37], P_3[45], G_3[45], P_3[37], G_4[45], P_4[45]);
    black_cell level_3_46(G_3[38], P_3[46], G_3[46], P_3[38], G_4[46], P_4[46]);
    black_cell level_3_47(G_3[39], P_3[47], G_3[47], P_3[39], G_4[47], P_4[47]);
    black_cell level_3_48(G_3[40], P_3[48], G_3[48], P_3[40], G_4[48], P_4[48]);
    black_cell level_3_49(G_3[41], P_3[49], G_3[49], P_3[41], G_4[49], P_4[49]);
    black_cell level_3_50(G_3[42], P_3[50], G_3[50], P_3[42], G_4[50], P_4[50]);
    black_cell level_3_51(G_3[43], P_3[51], G_3[51], P_3[43], G_4[51], P_4[51]);
    black_cell level_3_52(G_3[44], P_3[52], G_3[52], P_3[44], G_4[52], P_4[52]);
    black_cell level_3_53(G_3[45], P_3[53], G_3[53], P_3[45], G_4[53], P_4[53]);
    black_cell level_3_54(G_3[46], P_3[54], G_3[54], P_3[46], G_4[54], P_4[54]);
    black_cell level_3_55(G_3[47], P_3[55], G_3[55], P_3[47], G_4[55], P_4[55]);
    black_cell level_3_56(G_3[48], P_3[56], G_3[56], P_3[48], G_4[56], P_4[56]);
    black_cell level_3_57(G_3[49], P_3[57], G_3[57], P_3[49], G_4[57], P_4[57]);
    black_cell level_3_58(G_3[50], P_3[58], G_3[58], P_3[50], G_4[58], P_4[58]);
    black_cell level_3_59(G_3[51], P_3[59], G_3[59], P_3[51], G_4[59], P_4[59]);
    black_cell level_3_60(G_3[52], P_3[60], G_3[60], P_3[52], G_4[60], P_4[60]);
    black_cell level_3_61(G_3[53], P_3[61], G_3[61], P_3[53], G_4[61], P_4[61]);
    black_cell level_3_62(G_3[54], P_3[62], G_3[62], P_3[54], G_4[62], P_4[62]);
    black_cell level_3_63(G_3[55], P_3[63], G_3[63], P_3[55], G_4[63], P_4[63]);

    /*Stage 5*/
    gray_cell level_5_15(cin, P_4[15], G_4[15], G_5[15]);
    gray_cell level_5_16(G_1[0], P_4[16], G_4[16], G_5[16]);
    gray_cell level_5_17(G_2[1], P_4[17], G_4[17], G_5[17]);
    gray_cell level_5_18(G_2[2], P_4[18], G_4[18], G_5[18]);
    gray_cell level_5_19(G_3[3], P_4[19], G_4[19], G_5[19]);
    gray_cell level_5_20(G_3[4], P_4[20], G_4[20], G_5[20]);
    gray_cell level_5_21(G_3[5], P_4[21], G_4[21], G_5[21]);
    gray_cell level_5_22(G_3[6], P_4[22], G_4[22], G_5[22]);
    gray_cell level_5_23(G_4[7], P_4[23], G_4[23], G_5[23]);
    gray_cell level_5_24(G_4[8], P_4[24], G_4[24], G_5[24]);
    gray_cell level_5_25(G_4[9], P_4[25], G_4[25], G_5[25]);
    gray_cell level_5_26(G_4[10], P_4[26], G_4[26], G_5[26]);
    gray_cell level_5_27(G_4[11], P_4[27], G_4[27], G_5[27]);
    gray_cell level_5_28(G_4[12], P_4[28], G_4[28], G_5[28]);
    gray_cell level_5_29(G_4[13], P_4[29], G_4[29], G_5[29]);
    gray_cell level_5_30(G_4[14], P_4[30], G_4[30], G_5[30]);
    black_cell level_4_31(G_4[15], P_4[31], G_4[31], P_4[15], G_5[31], P_5[31]);
    black_cell level_4_32(G_4[16], P_4[32], G_4[32], P_4[16], G_5[32], P_5[32]);
    black_cell level_4_33(G_4[17], P_4[33], G_4[33], P_4[17], G_5[33], P_5[33]);
    black_cell level_4_34(G_4[18], P_4[34], G_4[34], P_4[18], G_5[34], P_5[34]);
    black_cell level_4_35(G_4[19], P_4[35], G_4[35], P_4[19], G_5[35], P_5[35]);
    black_cell level_4_36(G_4[20], P_4[36], G_4[36], P_4[20], G_5[36], P_5[36]);
    black_cell level_4_37(G_4[21], P_4[37], G_4[37], P_4[21], G_5[37], P_5[37]);
    black_cell level_4_38(G_4[22], P_4[38], G_4[38], P_4[22], G_5[38], P_5[38]);
    black_cell level_4_39(G_4[23], P_4[39], G_4[39], P_4[23], G_5[39], P_5[39]);
    black_cell level_4_40(G_4[24], P_4[40], G_4[40], P_4[24], G_5[40], P_5[40]);
    black_cell level_4_41(G_4[25], P_4[41], G_4[41], P_4[25], G_5[41], P_5[41]);
    black_cell level_4_42(G_4[26], P_4[42], G_4[42], P_4[26], G_5[42], P_5[42]);
    black_cell level_4_43(G_4[27], P_4[43], G_4[43], P_4[27], G_5[43], P_5[43]);
    black_cell level_4_44(G_4[28], P_4[44], G_4[44], P_4[28], G_5[44], P_5[44]);
    black_cell level_4_45(G_4[29], P_4[45], G_4[45], P_4[29], G_5[45], P_5[45]);
    black_cell level_4_46(G_4[30], P_4[46], G_4[46], P_4[30], G_5[46], P_5[46]);
    black_cell level_4_47(G_4[31], P_4[47], G_4[47], P_4[31], G_5[47], P_5[47]);
    black_cell level_4_48(G_4[32], P_4[48], G_4[48], P_4[32], G_5[48], P_5[48]);
    black_cell level_4_49(G_4[33], P_4[49], G_4[49], P_4[33], G_5[49], P_5[49]);
    black_cell level_4_50(G_4[34], P_4[50], G_4[50], P_4[34], G_5[50], P_5[50]);
    black_cell level_4_51(G_4[35], P_4[51], G_4[51], P_4[35], G_5[51], P_5[51]);
    black_cell level_4_52(G_4[36], P_4[52], G_4[52], P_4[36], G_5[52], P_5[52]);
    black_cell level_4_53(G_4[37], P_4[53], G_4[53], P_4[37], G_5[53], P_5[53]);
    black_cell level_4_54(G_4[38], P_4[54], G_4[54], P_4[38], G_5[54], P_5[54]);
    black_cell level_4_55(G_4[39], P_4[55], G_4[55], P_4[39], G_5[55], P_5[55]);
    black_cell level_4_56(G_4[40], P_4[56], G_4[56], P_4[40], G_5[56], P_5[56]);
    black_cell level_4_57(G_4[41], P_4[57], G_4[57], P_4[41], G_5[57], P_5[57]);
    black_cell level_4_58(G_4[42], P_4[58], G_4[58], P_4[42], G_5[58], P_5[58]);
    black_cell level_4_59(G_4[43], P_4[59], G_4[59], P_4[43], G_5[59], P_5[59]);
    black_cell level_4_60(G_4[44], P_4[60], G_4[60], P_4[44], G_5[60], P_5[60]);
    black_cell level_4_61(G_4[45], P_4[61], G_4[61], P_4[45], G_5[61], P_5[61]);
    black_cell level_4_62(G_4[46], P_4[62], G_4[62], P_4[46], G_5[62], P_5[62]);
    black_cell level_4_63(G_4[47], P_4[63], G_4[63], P_4[47], G_5[63], P_5[63]);

    /*Stage 6*/
    gray_cell level_6_31(cin, P_5[31], G_5[31], G_6[31]);
    gray_cell level_6_32(G_1[0], P_5[32], G_5[32], G_6[32]);
    gray_cell level_6_33(G_2[1], P_5[33], G_5[33], G_6[33]);
    gray_cell level_6_34(G_2[2], P_5[34], G_5[34], G_6[34]);
    gray_cell level_6_35(G_3[3], P_5[35], G_5[35], G_6[35]);
    gray_cell level_6_36(G_3[4], P_5[36], G_5[36], G_6[36]);
    gray_cell level_6_37(G_3[5], P_5[37], G_5[37], G_6[37]);
    gray_cell level_6_38(G_3[6], P_5[38], G_5[38], G_6[38]);
    gray_cell level_6_39(G_4[7], P_5[39], G_5[39], G_6[39]);
    gray_cell level_6_40(G_4[8], P_5[40], G_5[40], G_6[40]);
    gray_cell level_6_41(G_4[9], P_5[41], G_5[41], G_6[41]);
    gray_cell level_6_42(G_4[10], P_5[42], G_5[42], G_6[42]);
    gray_cell level_6_43(G_4[11], P_5[43], G_5[43], G_6[43]);
    gray_cell level_6_44(G_4[12], P_5[44], G_5[44], G_6[44]);
    gray_cell level_6_45(G_4[13], P_5[45], G_5[45], G_6[45]);
    gray_cell level_6_46(G_4[14], P_5[46], G_5[46], G_6[46]);
    gray_cell level_6_47(G_5[15], P_5[47], G_5[47], G_6[47]);
    gray_cell level_6_48(G_5[16], P_5[48], G_5[48], G_6[48]);
    gray_cell level_6_49(G_5[17], P_5[49], G_5[49], G_6[49]);
    gray_cell level_6_50(G_5[18], P_5[50], G_5[50], G_6[50]);
    gray_cell level_6_51(G_5[19], P_5[51], G_5[51], G_6[51]);
    gray_cell level_6_52(G_5[20], P_5[52], G_5[52], G_6[52]);
    gray_cell level_6_53(G_5[21], P_5[53], G_5[53], G_6[53]);
    gray_cell level_6_54(G_5[22], P_5[54], G_5[54], G_6[54]);
    gray_cell level_6_55(G_5[23], P_5[55], G_5[55], G_6[55]);
    gray_cell level_6_56(G_5[24], P_5[56], G_5[56], G_6[56]);
    gray_cell level_6_57(G_5[25], P_5[57], G_5[57], G_6[57]);
    gray_cell level_6_58(G_5[26], P_5[58], G_5[58], G_6[58]);
    gray_cell level_6_59(G_5[27], P_5[59], G_5[59], G_6[59]);
    gray_cell level_6_60(G_5[28], P_5[60], G_5[60], G_6[60]);
    gray_cell level_6_61(G_5[29], P_5[61], G_5[61], G_6[61]);
    gray_cell level_6_62(G_5[30], P_5[62], G_5[62], G_6[62]);
    black_cell level_5_63(G_5[31], P_5[63], G_5[63], P_5[31], G_6[63], P_6[63]);

    /*Stage 7*/
    gray_cell level_7_63(cin, P_6[63], G_6[63], cout);

    assign sum[0] = cin    ^ P_0[0];
    assign sum[1] = G_1[0] ^ P_0[1];
    assign sum[2] = G_2[1] ^ P_0[2];
    assign sum[3] = G_2[2] ^ P_0[3];
    assign sum[4] = G_3[3] ^ P_0[4];
    assign sum[5] = G_3[4] ^ P_0[5];
    assign sum[6] = G_3[5] ^ P_0[6];
    assign sum[7] = G_3[6] ^ P_0[7];
    assign sum[8] = G_4[7] ^ P_0[8];
    assign sum[9] = G_4[8] ^ P_0[9];
    assign sum[10] = G_4[9] ^ P_0[10];
    assign sum[11] = G_4[10] ^ P_0[11];
    assign sum[12] = G_4[11] ^ P_0[12];
    assign sum[13] = G_4[12] ^ P_0[13];
    assign sum[14] = G_4[13] ^ P_0[14];
    assign sum[15] = G_4[14] ^ P_0[15];
    assign sum[16] = G_5[15] ^ P_0[16];
    assign sum[17] = G_5[16] ^ P_0[17];
    assign sum[18] = G_5[17] ^ P_0[18];
    assign sum[19] = G_5[18] ^ P_0[19];
    assign sum[20] = G_5[19] ^ P_0[20];
    assign sum[21] = G_5[20] ^ P_0[21];
    assign sum[22] = G_5[21] ^ P_0[22];
    assign sum[23] = G_5[22] ^ P_0[23];
    assign sum[24] = G_5[23] ^ P_0[24];
    assign sum[25] = G_5[24] ^ P_0[25];
    assign sum[26] = G_5[25] ^ P_0[26];
    assign sum[27] = G_5[26] ^ P_0[27];
    assign sum[28] = G_5[27] ^ P_0[28];
    assign sum[29] = G_5[28] ^ P_0[29];
    assign sum[30] = G_5[29] ^ P_0[30];
    assign sum[31] = G_5[30] ^ P_0[31];
    assign sum[32] = G_6[31] ^ P_0[32];
    assign sum[33] = G_6[32] ^ P_0[33];
    assign sum[34] = G_6[33] ^ P_0[34];
    assign sum[35] = G_6[34] ^ P_0[35];
    assign sum[36] = G_6[35] ^ P_0[36];
    assign sum[37] = G_6[36] ^ P_0[37];
    assign sum[38] = G_6[37] ^ P_0[38];
    assign sum[39] = G_6[38] ^ P_0[39];
    assign sum[40] = G_6[39] ^ P_0[40];
    assign sum[41] = G_6[40] ^ P_0[41];
    assign sum[42] = G_6[41] ^ P_0[42];
    assign sum[43] = G_6[42] ^ P_0[43];
    assign sum[44] = G_6[43] ^ P_0[44];
    assign sum[45] = G_6[44] ^ P_0[45];
    assign sum[46] = G_6[45] ^ P_0[46];
    assign sum[47] = G_6[46] ^ P_0[47];
    assign sum[48] = G_6[47] ^ P_0[48];
    assign sum[49] = G_6[48] ^ P_0[49];
    assign sum[50] = G_6[49] ^ P_0[50];
    assign sum[51] = G_6[50] ^ P_0[51];
    assign sum[52] = G_6[51] ^ P_0[52];
    assign sum[53] = G_6[52] ^ P_0[53];
    assign sum[54] = G_6[53] ^ P_0[54];
    assign sum[55] = G_6[54] ^ P_0[55];
    assign sum[56] = G_6[55] ^ P_0[56];
    assign sum[57] = G_6[56] ^ P_0[57];
    assign sum[58] = G_6[57] ^ P_0[58];
    assign sum[59] = G_6[58] ^ P_0[59];
    assign sum[60] = G_6[59] ^ P_0[60];
    assign sum[61] = G_6[60] ^ P_0[61];
    assign sum[62] = G_6[61] ^ P_0[62];
    assign sum[63] = G_6[62] ^ P_0[63];
endmodule

module gray_cell(Gk_j, Pi_k, Gi_k, G);
    input Gk_j, Pi_k, Gi_k;
    output G;
    wire Y;
    and(Y, Gk_j, Pi_k);
    or(G, Y, Gi_k);
endmodule

module black_cell(Gk_j, Pi_k, Gi_k, Pk_j, G, P);
    input Gk_j, Pi_k, Gi_k, Pk_j;
    output G, P;
    wire Y;
    and(Y, Gk_j, Pi_k);
    or(G, Gi_k, Y);
    and(P, Pk_j, Pi_k);
endmodule
