module multiplier_32bits_version13(product, A, B);

    /*
     * Area: 
     * Power: mW
     * Timing: ns
     */

    output [63:0] product;
    input [31:0] A, B;

    wire [31:0] pp0;
    wire [31:0] pp1;
    wire [31:0] pp2;
    wire [31:0] pp3;
    wire [31:0] pp4;
    wire [31:0] pp5;
    wire [31:0] pp6;
    wire [31:0] pp7;
    wire [31:0] pp8;
    wire [31:0] pp9;
    wire [31:0] pp10;
    wire [31:0] pp11;
    wire [31:0] pp12;
    wire [31:0] pp13;
    wire [31:0] pp14;
    wire [31:0] pp15;
    wire [31:0] pp16;
    wire [31:0] pp17;
    wire [31:0] pp18;
    wire [31:0] pp19;
    wire [31:0] pp20;
    wire [31:0] pp21;
    wire [31:0] pp22;
    wire [31:0] pp23;
    wire [31:0] pp24;
    wire [31:0] pp25;
    wire [31:0] pp26;
    wire [31:0] pp27;
    wire [31:0] pp28;
    wire [31:0] pp29;
    wire [31:0] pp30;
    wire [31:0] pp31;


    assign pp0 = A[0] ? B: 32'b00000000000000000000000000000000;
    assign pp1 = A[1] ? B: 32'b00000000000000000000000000000000;
    assign pp2 = A[2] ? B: 32'b00000000000000000000000000000000;
    assign pp3 = A[3] ? B: 32'b00000000000000000000000000000000;
    assign pp4 = A[4] ? B: 32'b00000000000000000000000000000000;
    assign pp5 = A[5] ? B: 32'b00000000000000000000000000000000;
    assign pp6 = A[6] ? B: 32'b00000000000000000000000000000000;
    assign pp7 = A[7] ? B: 32'b00000000000000000000000000000000;
    assign pp8 = A[8] ? B: 32'b00000000000000000000000000000000;
    assign pp9 = A[9] ? B: 32'b00000000000000000000000000000000;
    assign pp10 = A[10] ? B: 32'b00000000000000000000000000000000;
    assign pp11 = A[11] ? B: 32'b00000000000000000000000000000000;
    assign pp12 = A[12] ? B: 32'b00000000000000000000000000000000;
    assign pp13 = A[13] ? B: 32'b00000000000000000000000000000000;
    assign pp14 = A[14] ? B: 32'b00000000000000000000000000000000;
    assign pp15 = A[15] ? B: 32'b00000000000000000000000000000000;
    assign pp16 = A[16] ? B: 32'b00000000000000000000000000000000;
    assign pp17 = A[17] ? B: 32'b00000000000000000000000000000000;
    assign pp18 = A[18] ? B: 32'b00000000000000000000000000000000;
    assign pp19 = A[19] ? B: 32'b00000000000000000000000000000000;
    assign pp20 = A[20] ? B: 32'b00000000000000000000000000000000;
    assign pp21 = A[21] ? B: 32'b00000000000000000000000000000000;
    assign pp22 = A[22] ? B: 32'b00000000000000000000000000000000;
    assign pp23 = A[23] ? B: 32'b00000000000000000000000000000000;
    assign pp24 = A[24] ? B: 32'b00000000000000000000000000000000;
    assign pp25 = A[25] ? B: 32'b00000000000000000000000000000000;
    assign pp26 = A[26] ? B: 32'b00000000000000000000000000000000;
    assign pp27 = A[27] ? B: 32'b00000000000000000000000000000000;
    assign pp28 = A[28] ? B: 32'b00000000000000000000000000000000;
    assign pp29 = A[29] ? B: 32'b00000000000000000000000000000000;
    assign pp30 = A[30] ? B: 32'b00000000000000000000000000000000;
    assign pp31 = A[31] ? B: 32'b00000000000000000000000000000000;


    /*Stage 1*/
    wire[3:0] s1, in1_1, in1_2;
    wire c1;
    assign in1_1 = {pp0[19],pp0[20],pp0[21],pp0[22]};
    assign in1_2 = {pp1[18],pp1[19],pp1[20],pp1[21]};
    CLA_4 KS_1(s1, c1, in1_1, in1_2);
    wire[3:0] s2, in2_1, in2_2;
    wire c2;
    assign in2_1 = {pp2[18],pp2[19],pp2[20],pp0[23]};
    assign in2_2 = {pp3[17],pp3[18],pp3[19],pp1[22]};
    CLA_4 KS_2(s2, c2, in2_1, in2_2);
    wire[3:0] s3, in3_1, in3_2;
    wire c3;
    assign in3_1 = {pp4[17],pp4[18],pp2[21],pp0[24]};
    assign in3_2 = {pp5[16],pp5[17],pp3[20],pp1[23]};
    CLA_4 KS_3(s3, c3, in3_1, in3_2);
    wire[3:0] s4, in4_1, in4_2;
    wire c4;
    assign in4_1 = {pp6[16],pp4[19],pp2[22],pp0[25]};
    assign in4_2 = {pp7[15],pp5[18],pp3[21],pp1[24]};
    CLA_4 KS_4(s4, c4, in4_1, in4_2);
    wire[3:0] s5, in5_1, in5_2;
    wire c5;
    assign in5_1 = {pp6[17],pp4[20],pp2[23],pp0[26]};
    assign in5_2 = {pp7[16],pp5[19],pp3[22],pp1[25]};
    CLA_4 KS_5(s5, c5, in5_1, in5_2);
    wire[3:0] s6, in6_1, in6_2;
    wire c6;
    assign in6_1 = {pp9[14],pp6[18],pp4[21],pp2[24]};
    assign in6_2 = {pp10[13],pp7[17],pp5[20],pp3[23]};
    CLA_4_c KS_6(s6, c6, in6_1, in6_2, pp8[15]);
    wire[3:0] s7, in7_1, in7_2;
    wire c7;
    assign in7_1 = {pp8[16],pp6[19],pp4[22],pp0[27]};
    assign in7_2 = {pp9[15],pp7[18],pp5[21],pp1[26]};
    CLA_4 KS_7(s7, c7, in7_1, in7_2);
    wire[3:0] s8, in8_1, in8_2;
    wire c8;
    assign in8_1 = {pp11[13],pp8[17],pp6[20],pp2[25]};
    assign in8_2 = {pp12[12],pp9[16],pp7[19],pp3[24]};
    CLA_4_c KS_8(s8, c8, in8_1, in8_2, pp10[14]);
    wire[3:0] s9, in9_1, in9_2;
    wire c9;
    assign in9_1 = {pp10[15],pp8[18],pp4[23],pp0[28]};
    assign in9_2 = {pp11[14],pp9[17],pp5[22],pp1[27]};
    CLA_4 KS_9(s9, c9, in9_1, in9_2);
    wire[3:0] s10, in10_1, in10_2;
    wire c10;
    assign in10_1 = {pp13[12],pp10[16],pp6[21],pp2[26]};
    assign in10_2 = {pp14[11],pp11[15],pp7[20],pp3[25]};
    CLA_4_c KS_10(s10, c10, in10_1, in10_2, pp12[13]);
    wire[3:0] s11, in11_1, in11_2;
    wire c11;
    assign in11_1 = {pp12[14],pp8[19],pp4[24],pp0[29]};
    assign in11_2 = {pp13[13],pp9[18],pp5[23],pp1[28]};
    CLA_4 KS_11(s11, c11, in11_1, in11_2);
    wire[3:0] s12, in12_1, in12_2;
    wire c12;
    assign in12_1 = {pp15[11],pp10[17],pp6[22],pp2[27]};
    assign in12_2 = {pp16[10],pp11[16],pp7[21],pp3[26]};
    CLA_4_c KS_12(s12, c12, in12_1, in12_2, pp14[12]);
    wire[3:0] s13, in13_1, in13_2;
    wire c13;
    assign in13_1 = {pp12[15],pp8[20],pp4[25],pp0[30]};
    assign in13_2 = {pp13[14],pp9[19],pp5[24],pp1[29]};
    CLA_4 KS_13(s13, c13, in13_1, in13_2);
    wire[3:0] s14, in14_1, in14_2;
    wire c14;
    assign in14_1 = {pp14[13],pp10[18],pp6[23],pp2[28]};
    assign in14_2 = {pp15[12],pp11[17],pp7[22],pp3[27]};
    CLA_4 KS_14(s14, c14, in14_1, in14_2);
    wire[3:0] s15, in15_1, in15_2;
    wire c15;
    assign in15_1 = {pp16[11],pp12[16],pp8[21],pp4[26]};
    assign in15_2 = {pp17[10],pp13[15],pp9[20],pp5[25]};
    CLA_4 KS_15(s15, c15, in15_1, in15_2);
    wire[3:0] s16, in16_1, in16_2;
    wire c16;
    assign in16_1 = {pp19[8],pp14[14],pp10[19],pp6[24]};
    assign in16_2 = {pp20[7],pp15[13],pp11[18],pp7[23]};
    CLA_4_c KS_16(s16, c16, in16_1, in16_2, pp18[9]);
    wire[3:0] s17, in17_1, in17_2;
    wire c17;
    assign in17_1 = {pp16[12],pp12[17],pp8[22],pp0[31]};
    assign in17_2 = {pp17[11],pp13[16],pp9[21],pp1[30]};
    CLA_4 KS_17(s17, c17, in17_1, in17_2);
    wire[3:0] s18, in18_1, in18_2;
    wire c18;
    assign in18_1 = {pp18[10],pp14[15],pp10[20],pp2[29]};
    assign in18_2 = {pp19[9],pp15[14],pp11[19],pp3[28]};
    CLA_4 KS_18(s18, c18, in18_1, in18_2);
    wire[3:0] s19, in19_1, in19_2;
    wire c19;
    assign in19_1 = {pp21[7],pp16[13],pp12[18],pp4[27]};
    assign in19_2 = {pp22[6],pp17[12],pp13[17],pp5[26]};
    CLA_4_c KS_19(s19, c19, in19_1, in19_2, pp20[8]);
    wire[3:0] s20, in20_1, in20_2;
    wire c20;
    assign in20_1 = {pp18[11],pp14[16],pp6[25],pp1[31]};
    assign in20_2 = {pp19[10],pp15[15],pp7[24],pp2[30]};
    CLA_4 KS_20(s20, c20, in20_1, in20_2);
    wire[3:0] s21, in21_1, in21_2;
    wire c21;
    assign in21_1 = {pp20[9],pp16[14],pp8[23],pp3[29]};
    assign in21_2 = {pp21[8],pp17[13],pp9[22],pp4[28]};
    CLA_4 KS_21(s21, c21, in21_1, in21_2);
    wire[3:0] s22, in22_1, in22_2;
    wire c22;
    assign in22_1 = {pp23[6],pp18[12],pp10[21],pp5[27]};
    assign in22_2 = {pp24[5],pp19[11],pp11[20],pp6[26]};
    CLA_4_c KS_22(s22, c22, in22_1, in22_2, pp22[7]);
    wire[3:0] s23, in23_1, in23_2;
    wire c23;
    assign in23_1 = {pp20[10],pp12[19],pp7[25],pp2[31]};
    assign in23_2 = {pp21[9],pp13[18],pp8[24],pp3[30]};
    CLA_4 KS_23(s23, c23, in23_1, in23_2);
    wire[3:0] s24, in24_1, in24_2;
    wire c24;
    assign in24_1 = {pp22[8],pp14[17],pp9[23],pp4[29]};
    assign in24_2 = {pp23[7],pp15[16],pp10[22],pp5[28]};
    CLA_4 KS_24(s24, c24, in24_1, in24_2);
    wire[3:0] s25, in25_1, in25_2;
    wire c25;
    assign in25_1 = {pp25[5],pp16[15],pp11[21],pp6[27]};
    assign in25_2 = {pp26[4],pp17[14],pp12[20],pp7[26]};
    CLA_4_c KS_25(s25, c25, in25_1, in25_2, pp24[6]);
    wire[3:0] s26, in26_1, in26_2;
    wire c26;
    assign in26_1 = {pp18[13],pp13[19],pp8[25],pp3[31]};
    assign in26_2 = {pp19[12],pp14[18],pp9[24],pp4[30]};
    CLA_4 KS_26(s26, c26, in26_1, in26_2);
    wire[3:0] s27, in27_1, in27_2;
    wire c27;
    assign in27_1 = {pp20[11],pp15[17],pp10[23],pp5[29]};
    assign in27_2 = {pp21[10],pp16[16],pp11[22],pp6[28]};
    CLA_4 KS_27(s27, c27, in27_1, in27_2);
    wire[3:0] s28, in28_1, in28_2;
    wire c28;
    assign in28_1 = {pp22[9],pp17[15],pp12[21],pp7[27]};
    assign in28_2 = {pp23[8],pp18[14],pp13[20],pp8[26]};
    CLA_4 KS_28(s28, c28, in28_1, in28_2);
    wire[3:0] s29, in29_1, in29_2;
    wire c29;
    assign in29_1 = {pp24[7],pp19[13],pp14[19],pp9[25]};
    assign in29_2 = {pp25[6],pp20[12],pp15[18],pp10[24]};
    CLA_4 KS_29(s29, c29, in29_1, in29_2);
    wire[3:0] s30, in30_1, in30_2;
    wire c30;
    assign in30_1 = {pp26[5],pp21[11],pp16[17],pp11[23]};
    assign in30_2 = {pp27[4],pp22[10],pp17[16],pp12[22]};
    CLA_4 KS_30(s30, c30, in30_1, in30_2);
    wire[3:0] s31, in31_1, in31_2;
    wire c31;
    assign in31_1 = {pp28[3],pp23[9],pp18[15],pp13[21]};
    assign in31_2 = {pp29[2],pp24[8],pp19[14],pp14[20]};
    CLA_4 KS_31(s31, c31, in31_1, in31_2);
    wire[3:0] s32, in32_1, in32_2;
    wire c32;
    assign in32_1 = {pp31[0],pp25[7],pp20[13],pp15[19]};
    assign in32_2 = {c13,pp26[6],pp21[12],pp16[18]};
    CLA_4_c KS_32(s32, c32, in32_1, in32_2, pp30[1]);
    wire[3:0] s33, in33_1, in33_2;
    wire c33;
    assign in33_1 = {pp27[5],pp22[11],pp17[17],pp4[31]};
    assign in33_2 = {pp28[4],pp23[10],pp18[16],pp5[30]};
    CLA_4 KS_33(s33, c33, in33_1, in33_2);
    wire[3:0] s34, in34_1, in34_2;
    wire c34;
    assign in34_1 = {pp30[2],pp24[9],pp19[15],pp6[29]};
    assign in34_2 = {pp31[1],pp25[8],pp20[14],pp7[28]};
    CLA_4_c KS_34(s34, c34, in34_1, in34_2, pp29[3]);
    wire[3:0] s35, in35_1, in35_2;
    wire c35;
    assign in35_1 = {pp27[6],pp21[13],pp8[27],pp5[31]};
    assign in35_2 = {pp28[5],pp22[12],pp9[26],pp6[30]};
    CLA_4_c KS_35(s35, c35, in35_1, in35_2, pp26[7]);
    wire[3:0] s36, in36_1, in36_2;
    wire c36;
    assign in36_1 = {pp23[11],pp10[25],pp7[29],pp6[31]};
    assign in36_2 = {pp24[10],pp11[24],pp8[28],pp7[30]};
    CLA_4 KS_36(s36, c36, in36_1, in36_2);
    wire[3:0] s37, in37_1, in37_2;
    wire c37;
    assign in37_1 = {pp26[8],pp12[23],pp9[27],pp8[29]};
    assign in37_2 = {pp27[7],pp13[22],pp10[26],pp9[28]};
    CLA_4_c KS_37(s37, c37, in37_1, in37_2, pp25[9]);
    wire[3:0] s38, in38_1, in38_2;
    wire c38;
    assign in38_1 = {pp14[21],pp11[25],pp10[27],pp7[31]};
    assign in38_2 = {pp15[20],pp12[24],pp11[26],pp8[30]};
    CLA_4 KS_38(s38, c38, in38_1, in38_2);
    wire[3:0] s39, in39_1, in39_2;
    wire c39;
    assign in39_1 = {pp16[19],pp13[23],pp12[25],pp9[29]};
    assign in39_2 = {pp17[18],pp14[22],pp13[24],pp10[28]};
    CLA_4 KS_39(s39, c39, in39_1, in39_2);
    wire[3:0] s40, in40_1, in40_2;
    wire c40;
    assign in40_1 = {pp18[17],pp15[21],pp14[23],pp11[27]};
    assign in40_2 = {pp19[16],pp16[20],pp15[22],pp12[26]};
    CLA_4 KS_40(s40, c40, in40_1, in40_2);
    wire[3:0] s41, in41_1, in41_2;
    wire c41;
    assign in41_1 = {pp20[15],pp17[19],pp16[21],pp13[25]};
    assign in41_2 = {pp21[14],pp18[18],pp17[20],pp14[24]};
    CLA_4 KS_41(s41, c41, in41_1, in41_2);
    wire[3:0] s42, in42_1, in42_2;
    wire c42;
    assign in42_1 = {pp22[13],pp19[17],pp18[19],pp15[23]};
    assign in42_2 = {pp23[12],pp20[16],pp19[18],pp16[22]};
    CLA_4 KS_42(s42, c42, in42_1, in42_2);
    wire[3:0] s43, in43_1, in43_2;
    wire c43;
    assign in43_1 = {pp24[11],pp21[15],pp20[17],pp17[21]};
    assign in43_2 = {pp25[10],pp22[14],pp21[16],pp18[20]};
    CLA_4 KS_43(s43, c43, in43_1, in43_2);
    wire[3:0] s44, in44_1, in44_2;
    wire c44;
    assign in44_1 = {pp26[9],pp23[13],pp22[15],pp19[19]};
    assign in44_2 = {pp27[8],pp24[12],pp23[14],pp20[18]};
    CLA_4 KS_44(s44, c44, in44_1, in44_2);
    wire[1:0] s45, in45_1, in45_2;
    wire c45;
    assign in45_1 = {pp28[7],pp25[11]};
    assign in45_2 = {pp29[6],pp26[10]};
    CLA_2 KS_45(s45, c45, in45_1, in45_2);
    wire[0:0] s46, in46_1, in46_2;
    wire c46;
    assign in46_1 = {pp30[5]};
    assign in46_2 = {pp31[4]};
    Half_Adder KS_46(s46, c46, in46_1, in46_2);
    wire[3:0] s47, in47_1, in47_2;
    wire c47;
    assign in47_1 = {c27,pp27[9],pp24[13],pp21[17]};
    assign in47_2 = {c28,pp28[8],pp25[12],pp22[16]};
    CLA_4_c KS_47(s47, c47, in47_1, in47_2, c26);
    wire[3:0] s48, in48_1, in48_2;
    wire c48;
    assign in48_1 = {pp8[31],pp9[31],pp10[31],pp11[31]};
    assign in48_2 = {pp9[30],pp10[30],pp11[30],pp12[30]};
    CLA_4 KS_48(s48, c48, in48_1, in48_2);
    wire[3:0] s49, in49_1, in49_2;
    wire c49;
    assign in49_1 = {pp10[29],pp11[29],pp12[29],pp13[29]};
    assign in49_2 = {pp11[28],pp12[28],pp13[28],pp14[28]};
    CLA_4 KS_49(s49, c49, in49_1, in49_2);
    wire[3:0] s50, in50_1, in50_2;
    wire c50;
    assign in50_1 = {pp12[27],pp13[27],pp14[27],pp15[27]};
    assign in50_2 = {pp13[26],pp14[26],pp15[26],pp16[26]};
    CLA_4 KS_50(s50, c50, in50_1, in50_2);
    wire[2:0] s51, in51_1, in51_2;
    wire c51;
    assign in51_1 = {pp14[25],pp15[25],pp16[25]};
    assign in51_2 = {pp15[24],pp16[24],pp17[24]};
    CLA_3 KS_51(s51, c51, in51_1, in51_2);
    wire[1:0] s52, in52_1, in52_2;
    wire c52;
    assign in52_1 = {pp16[23],pp17[23]};
    assign in52_2 = {pp17[22],pp18[22]};
    CLA_2 KS_52(s52, c52, in52_1, in52_2);
    wire[0:0] s53, in53_1, in53_2;
    wire c53;
    assign in53_1 = {pp18[21]};
    assign in53_2 = {pp19[20]};
    Half_Adder KS_53(s53, c53, in53_1, in53_2);
    wire[3:0] s54, in54_1, in54_2;
    wire c54;
    assign in54_1 = {pp20[19],pp19[21],pp18[23],pp17[25]};
    assign in54_2 = {pp21[18],pp20[20],pp19[22],pp18[24]};
    CLA_4 KS_54(s54, c54, in54_1, in54_2);
    wire[0:0] s55, in55_1, in55_2;
    wire c55;
    assign in55_1 = {pp22[17]};
    assign in55_2 = {pp23[16]};
    Half_Adder KS_55(s55, c55, in55_1, in55_2);
    wire[1:0] s56, in56_1, in56_2;
    wire c56;
    assign in56_1 = {pp24[15],pp21[19]};
    assign in56_2 = {pp25[14],pp22[18]};
    CLA_2 KS_56(s56, c56, in56_1, in56_2);
    wire[0:0] s57, in57_1, in57_2;
    wire c57;
    assign in57_1 = {pp26[13]};
    assign in57_2 = {pp27[12]};
    Half_Adder KS_57(s57, c57, in57_1, in57_2);
    wire[2:0] s58, in58_1, in58_2;
    wire c58;
    assign in58_1 = {pp28[11],pp23[17],pp20[21]};
    assign in58_2 = {pp29[10],pp24[16],pp21[20]};
    CLA_3 KS_58(s58, c58, in58_1, in58_2);
    wire[0:0] s59, in59_1, in59_2;
    wire c59;
    assign in59_1 = {pp31[8]};
    assign in59_2 = {c38};
    Full_Adder KS_59(s59, c59, in59_1, in59_2, pp30[9]);
    wire[1:0] s60, in60_1, in60_2;
    wire c60;
    assign in60_1 = {pp12[31],pp13[31]};
    assign in60_2 = {pp13[30],pp14[30]};
    CLA_2 KS_60(s60, c60, in60_1, in60_2);
    wire[0:0] s61, in61_1, in61_2;
    wire c61;
    assign in61_1 = {pp14[29]};
    assign in61_2 = {pp15[28]};
    Half_Adder KS_61(s61, c61, in61_1, in61_2);
    wire[2:0] s62, in62_1, in62_2;
    wire c62;
    assign in62_1 = {pp16[27],pp15[29],pp14[31]};
    assign in62_2 = {pp17[26],pp16[28],pp15[30]};
    CLA_3 KS_62(s62, c62, in62_1, in62_2);
    wire[0:0] s63, in63_1, in63_2;
    wire c63;
    assign in63_1 = {pp19[24]};
    assign in63_2 = {pp20[23]};
    Full_Adder KS_63(s63, c63, in63_1, in63_2, pp18[25]);

    /*Stage 2*/
    wire[3:0] s64, in64_1, in64_2;
    wire c64;
    assign in64_1 = {pp0[12],pp0[13],pp0[14],pp0[15]};
    assign in64_2 = {pp1[11],pp1[12],pp1[13],pp1[14]};
    CLA_4 KS_64(s64, c64, in64_1, in64_2);
    wire[3:0] s65, in65_1, in65_2;
    wire c65;
    assign in65_1 = {pp2[11],pp2[12],pp2[13],pp0[16]};
    assign in65_2 = {pp3[10],pp3[11],pp3[12],pp1[15]};
    CLA_4 KS_65(s65, c65, in65_1, in65_2);
    wire[3:0] s66, in66_1, in66_2;
    wire c66;
    assign in66_1 = {pp4[10],pp4[11],pp2[14],pp0[17]};
    assign in66_2 = {pp5[9],pp5[10],pp3[13],pp1[16]};
    CLA_4 KS_66(s66, c66, in66_1, in66_2);
    wire[3:0] s67, in67_1, in67_2;
    wire c67;
    assign in67_1 = {pp6[9],pp4[12],pp2[15],pp0[18]};
    assign in67_2 = {pp7[8],pp5[11],pp3[14],pp1[17]};
    CLA_4 KS_67(s67, c67, in67_1, in67_2);
    wire[3:0] s68, in68_1, in68_2;
    wire c68;
    assign in68_1 = {pp6[10],pp4[13],pp2[16],pp2[17]};
    assign in68_2 = {pp7[9],pp5[12],pp3[15],pp3[16]};
    CLA_4 KS_68(s68, c68, in68_1, in68_2);
    wire[3:0] s69, in69_1, in69_2;
    wire c69;
    assign in69_1 = {pp9[7],pp6[11],pp4[14],pp4[15]};
    assign in69_2 = {pp10[6],pp7[10],pp5[13],pp5[14]};
    CLA_4_c KS_69(s69, c69, in69_1, in69_2, pp8[8]);
    wire[3:0] s70, in70_1, in70_2;
    wire c70;
    assign in70_1 = {pp8[9],pp6[12],pp6[13],pp4[16]};
    assign in70_2 = {pp9[8],pp7[11],pp7[12],pp5[15]};
    CLA_4 KS_70(s70, c70, in70_1, in70_2);
    wire[3:0] s71, in71_1, in71_2;
    wire c71;
    assign in71_1 = {pp11[6],pp8[10],pp8[11],pp6[14]};
    assign in71_2 = {pp12[5],pp9[9],pp9[10],pp7[13]};
    CLA_4_c KS_71(s71, c71, in71_1, in71_2, pp10[7]);
    wire[3:0] s72, in72_1, in72_2;
    wire c72;
    assign in72_1 = {pp10[8],pp10[9],pp8[12],pp6[15]};
    assign in72_2 = {pp11[7],pp11[8],pp9[11],pp7[14]};
    CLA_4 KS_72(s72, c72, in72_1, in72_2);
    wire[3:0] s73, in73_1, in73_2;
    wire c73;
    assign in73_1 = {pp13[5],pp12[7],pp10[10],pp8[13]};
    assign in73_2 = {pp14[4],pp13[6],pp11[9],pp9[12]};
    CLA_4_c KS_73(s73, c73, in73_1, in73_2, pp12[6]);
    wire[3:0] s74, in74_1, in74_2;
    wire c74;
    assign in74_1 = {pp15[4],pp12[8],pp10[11],pp8[14]};
    assign in74_2 = {pp16[3],pp13[7],pp11[10],pp9[13]};
    CLA_4_c KS_74(s74, c74, in74_1, in74_2, pp14[5]);
    wire[3:0] s75, in75_1, in75_2;
    wire c75;
    assign in75_1 = {pp14[6],pp12[9],pp10[12],pp11[12]};
    assign in75_2 = {pp15[5],pp13[8],pp11[11],pp12[11]};
    CLA_4 KS_75(s75, c75, in75_1, in75_2);
    wire[3:0] s76, in76_1, in76_2;
    wire c76;
    assign in76_1 = {pp16[4],pp14[7],pp12[10],pp13[10]};
    assign in76_2 = {pp17[3],pp15[6],pp13[9],pp14[9]};
    CLA_4 KS_76(s76, c76, in76_1, in76_2);
    wire[3:0] s77, in77_1, in77_2;
    wire c77;
    assign in77_1 = {pp19[1],pp16[5],pp14[8],pp15[8]};
    assign in77_2 = {pp20[0],pp17[4],pp15[7],pp16[7]};
    CLA_4_c KS_77(s77, c77, in77_1, in77_2, pp18[2]);
    wire[3:0] s78, in78_1, in78_2;
    wire c78;
    assign in78_1 = {pp18[3],pp16[6],pp17[6],pp13[11]};
    assign in78_2 = {pp19[2],pp17[5],pp18[5],pp14[10]};
    CLA_4 KS_78(s78, c78, in78_1, in78_2);
    wire[3:0] s79, in79_1, in79_2;
    wire c79;
    assign in79_1 = {pp21[0],pp18[4],pp19[4],pp15[9]};
    assign in79_2 = {s1[2],pp19[3],pp20[3],pp16[8]};
    CLA_4_c KS_79(s79, c79, in79_1, in79_2, pp20[1]);
    wire[3:0] s80, in80_1, in80_2;
    wire c80;
    assign in80_1 = {pp20[2],pp21[2],pp17[7],pp15[10]};
    assign in80_2 = {pp21[1],pp22[1],pp18[6],pp16[9]};
    CLA_4 KS_80(s80, c80, in80_1, in80_2);
    wire[3:0] s81, in81_1, in81_2;
    wire c81;
    assign in81_1 = {s1[3],pp23[0],pp19[5],pp17[8]};
    assign in81_2 = {s2[2],c1,pp20[4],pp18[7]};
    CLA_4_c KS_81(s81, c81, in81_1, in81_2, pp22[0]);
    wire[3:0] s82, in82_1, in82_2;
    wire c82;
    assign in82_1 = {s2[3],pp21[3],pp19[6],pp17[9]};
    assign in82_2 = {s3[2],pp22[2],pp20[5],pp18[8]};
    CLA_4 KS_82(s82, c82, in82_1, in82_2);
    wire[3:0] s83, in83_1, in83_2;
    wire c83;
    assign in83_1 = {pp23[1],pp21[4],pp19[7],pp21[6]};
    assign in83_2 = {pp24[0],pp22[3],pp20[6],pp22[5]};
    CLA_4 KS_83(s83, c83, in83_1, in83_2);
    wire[3:0] s84, in84_1, in84_2;
    wire c84;
    assign in84_1 = {c2,pp23[2],pp21[5],pp23[4]};
    assign in84_2 = {s3[3],pp24[1],pp22[4],pp24[3]};
    CLA_4 KS_84(s84, c84, in84_1, in84_2);
    wire[3:0] s85, in85_1, in85_2;
    wire c85;
    assign in85_1 = {s4[2],pp25[0],pp23[3],pp25[2]};
    assign in85_2 = {s5[1],c3,pp24[2],pp26[1]};
    CLA_4 KS_85(s85, c85, in85_1, in85_2);
    wire[3:0] s86, in86_1, in86_2;
    wire c86;
    assign in86_1 = {s7[0],s4[3],pp25[1],pp27[0]};
    assign in86_2 = {s8[0],s5[2],pp26[0],c5};
    CLA_4_c KS_86(s86, c86, in86_1, in86_2, s6[1]);
    wire[3:0] s87, in87_1, in87_2;
    wire c87;
    assign in87_1 = {s7[1],c4,c6,pp23[5]};
    assign in87_2 = {s8[1],s5[3],s7[3],pp24[4]};
    CLA_4_c KS_87(s87, c87, in87_1, in87_2, s6[2]);
    wire[3:0] s88, in88_1, in88_2;
    wire c88;
    assign in88_1 = {s6[3],s8[3],pp25[3],pp25[4]};
    assign in88_2 = {s7[2],s9[2],pp26[2],pp26[3]};
    CLA_4 KS_88(s88, c88, in88_1, in88_2);
    wire[3:0] s89, in89_1, in89_2;
    wire c89;
    assign in89_1 = {s9[1],s10[2],pp27[1],pp27[2]};
    assign in89_2 = {s10[1],s11[1],pp28[0],pp28[1]};
    CLA_4_c KS_89(s89, c89, in89_1, in89_2, s8[2]);
    wire[3:0] s90, in90_1, in90_2;
    wire c90;
    assign in90_1 = {s12[1],c7,pp29[0],pp27[3]};
    assign in90_2 = {s13[0],c8,c9,pp28[2]};
    CLA_4 KS_90(s90, c90, in90_1, in90_2);
    wire[3:0] s91, in91_1, in91_2;
    wire c91;
    assign in91_1 = {s9[3],c10,pp29[1],c14};
    assign in91_2 = {s10[3],s11[3],pp30[0],c15};
    CLA_4 KS_91(s91, c91, in91_1, in91_2);
    wire[3:0] s92, in92_1, in92_2;
    wire c92;
    assign in92_1 = {s11[2],s12[3],c11,c16};
    assign in92_2 = {s12[2],s13[2],c12,s17[3]};
    CLA_4 KS_92(s92, c92, in92_1, in92_2);
    wire[3:0] s93, in93_1, in93_2;
    wire c93;
    assign in93_1 = {s13[1],s14[2],s13[3],s18[3]};
    assign in93_2 = {s14[1],s15[2],s14[3],s19[3]};
    CLA_4 KS_93(s93, c93, in93_1, in93_2);
    wire[3:0] s94, in94_1, in94_2;
    wire c94;
    assign in94_1 = {s15[1],s16[2],s15[3],s20[2]};
    assign in94_2 = {s16[1],s17[1],s16[3],s21[2]};
    CLA_4 KS_94(s94, c94, in94_1, in94_2);
    wire[3:0] s95, in95_1, in95_2;
    wire c95;
    assign in95_1 = {s17[0],s18[1],s17[2],s22[2]};
    assign in95_2 = {s18[0],s19[1],s18[2],s23[1]};
    CLA_4 KS_95(s95, c95, in95_1, in95_2);
    wire[3:0] s96, in96_1, in96_2;
    wire c96;
    assign in96_1 = {c83,s20[0],s19[2],s24[1]};
    assign in96_2 = {c84,s21[0],s20[1],s25[1]};
    CLA_4_c KS_96(s96, c96, in96_1, in96_2, s19[0]);
    wire[3:0] s97, in97_1, in97_2;
    wire c97;
    assign in97_1 = {s22[1],s26[0],1'b0,pp29[4]};
    assign in97_2 = {s23[0],s27[0],c17,pp30[3]};
    CLA_4_c KS_97(s97, c97, in97_1, in97_2, s21[1]);
    wire[3:0] s98, in98_1, in98_2;
    wire c98;
    assign in98_1 = {s28[0],c18,pp31[2],pp28[6]};
    assign in98_2 = {s29[0],c19,c20,pp29[5]};
    CLA_4 KS_98(s98, c98, in98_1, in98_2);
    wire[3:0] s99, in99_1, in99_2;
    wire c99;
    assign in99_1 = {s20[3],c21,pp30[4],c29};
    assign in99_2 = {s21[3],c22,pp31[3],c30};
    CLA_4 KS_99(s99, c99, in99_1, in99_2);
    wire[3:0] s100, in100_1, in100_2;
    wire c100;
    assign in100_1 = {s22[3],s23[3],c23,c31};
    assign in100_2 = {s23[2],s24[3],c24,c32};
    CLA_4 KS_100(s100, c100, in100_1, in100_2);
    wire[3:0] s101, in101_1, in101_2;
    wire c101;
    assign in101_1 = {s24[2],s25[3],c25,s33[3]};
    assign in101_2 = {s25[2],s26[2],s26[3],s34[3]};
    CLA_4 KS_101(s101, c101, in101_1, in101_2);
    wire[3:0] s102, in102_1, in102_2;
    wire c102;
    assign in102_1 = {s26[1],s27[2],s27[3],s35[2]};
    assign in102_2 = {s27[1],s28[2],s28[3],s36[1]};
    CLA_4 KS_102(s102, c102, in102_1, in102_2);
    wire[3:0] s103, in103_1, in103_2;
    wire c103;
    assign in103_1 = {s28[1],s29[2],s29[3],s37[1]};
    assign in103_2 = {s29[1],s30[2],s30[3],s38[0]};
    CLA_4 KS_103(s103, c103, in103_1, in103_2);
    wire[3:0] s104, in104_1, in104_2;
    wire c104;
    assign in104_1 = {s30[1],s31[2],s31[3],s39[0]};
    assign in104_2 = {s31[1],s32[2],s32[3],s40[0]};
    CLA_4 KS_104(s104, c104, in104_1, in104_2);
    wire[0:0] s105, in105_1, in105_2;
    wire c105;
    assign in105_1 = {s32[1]};
    assign in105_2 = {s33[0]};
    Half_Adder KS_105(s105, c105, in105_1, in105_2);
    wire[3:0] s106, in106_1, in106_2;
    wire c106;
    assign in106_1 = {s34[0],s33[1],s33[2],s41[0]};
    assign in106_2 = {c91,s34[1],s34[2],s42[0]};
    CLA_4 KS_106(s106, c106, in106_1, in106_2);
    wire[0:0] s107, in107_1, in107_2;
    wire c107;
    assign in107_1 = {c92};
    assign in107_2 = {c93};
    Half_Adder KS_107(s107, c107, in107_1, in107_2);
    wire[3:0] s108, in108_1, in108_2;
    wire c108;
    assign in108_1 = {c95,s35[0],s35[1],s43[0]};
    assign in108_2 = {c96,s97[3],s36[0],s44[0]};
    CLA_4_c KS_108(s108, c108, in108_1, in108_2, c94);
    wire[3:0] s109, in109_1, in109_2;
    wire c109;
    assign in109_1 = {pp29[7],pp26[11],pp23[15],c39};
    assign in109_2 = {pp30[6],pp27[10],pp24[14],c40};
    CLA_4 KS_109(s109, c109, in109_1, in109_2);
    wire[3:0] s110, in110_1, in110_2;
    wire c110;
    assign in110_1 = {pp31[5],pp28[9],pp25[13],c41};
    assign in110_2 = {c33,pp29[8],pp26[12],c42};
    CLA_4 KS_110(s110, c110, in110_1, in110_2);
    wire[3:0] s111, in111_1, in111_2;
    wire c111;
    assign in111_1 = {c34,pp30[7],pp27[11],c43};
    assign in111_2 = {s35[3],pp31[6],pp28[10],c44};
    CLA_4 KS_111(s111, c111, in111_1, in111_2);
    wire[3:0] s112, in112_1, in112_2;
    wire c112;
    assign in112_1 = {s36[2],c35,pp29[9],c47};
    assign in112_2 = {s37[2],s36[3],pp30[8],s48[0]};
    CLA_4 KS_112(s112, c112, in112_1, in112_2);
    wire[3:0] s113, in113_1, in113_2;
    wire c113;
    assign in113_1 = {s38[1],s37[3],pp31[7],s49[0]};
    assign in113_2 = {s39[1],s38[2],c36,s50[0]};
    CLA_4 KS_113(s113, c113, in113_1, in113_2);
    wire[3:0] s114, in114_1, in114_2;
    wire c114;
    assign in114_1 = {s40[1],s39[2],c37,s51[0]};
    assign in114_2 = {s41[1],s40[2],s38[3],s52[0]};
    CLA_4 KS_114(s114, c114, in114_1, in114_2);
    wire[3:0] s115, in115_1, in115_2;
    wire c115;
    assign in115_1 = {s42[1],s41[2],s39[3],s53[0]};
    assign in115_2 = {s43[1],s42[2],s40[3],s54[0]};
    CLA_4 KS_115(s115, c115, in115_1, in115_2);
    wire[0:0] s116, in116_1, in116_2;
    wire c116;
    assign in116_1 = {s44[1]};
    assign in116_2 = {s45[1]};
    Half_Adder KS_116(s116, c116, in116_1, in116_2);
    wire[3:0] s117, in117_1, in117_2;
    wire c117;
    assign in117_1 = {c46,s43[2],s41[3],s55[0]};
    assign in117_2 = {s47[1],s44[2],s42[3],s56[0]};
    CLA_4 KS_117(s117, c117, in117_1, in117_2);
    wire[0:0] s118, in118_1, in118_2;
    wire c118;
    assign in118_1 = {c99};
    assign in118_2 = {c100};
    Half_Adder KS_118(s118, c118, in118_1, in118_2);
    wire[1:0] s119, in119_1, in119_2;
    wire c119;
    assign in119_1 = {c101,c45};
    assign in119_2 = {c102,s47[2]};
    CLA_2 KS_119(s119, c119, in119_1, in119_2);
    wire[0:0] s120, in120_1, in120_2;
    wire c120;
    assign in120_1 = {c103};
    assign in120_2 = {c104};
    Half_Adder KS_120(s120, c120, in120_1, in120_2);
    wire[2:0] s121, in121_1, in121_2;
    wire c121;
    assign in121_1 = {c108,s109[1],s43[3]};
    assign in121_2 = {s109[0],s110[1],s44[3]};
    CLA_3_c KS_121(s121, c121, in121_1, in121_2, c106);
    wire[3:0] s122, in122_1, in122_2;
    wire c122;
    assign in122_1 = {pp25[15],pp22[19],pp19[23],pp21[22]};
    assign in122_2 = {pp26[14],pp23[18],pp20[22],pp22[21]};
    CLA_4 KS_122(s122, c122, in122_1, in122_2);
    wire[3:0] s123, in123_1, in123_2;
    wire c123;
    assign in123_1 = {pp27[13],pp24[17],pp21[21],pp23[20]};
    assign in123_2 = {pp28[12],pp25[16],pp22[20],pp24[19]};
    CLA_4 KS_123(s123, c123, in123_1, in123_2);
    wire[3:0] s124, in124_1, in124_2;
    wire c124;
    assign in124_1 = {pp29[11],pp26[15],pp23[19],pp25[18]};
    assign in124_2 = {pp30[10],pp27[14],pp24[18],pp26[17]};
    CLA_4 KS_124(s124, c124, in124_1, in124_2);
    wire[3:0] s125, in125_1, in125_2;
    wire c125;
    assign in125_1 = {pp31[9],pp28[13],pp25[17],pp27[16]};
    assign in125_2 = {s48[1],pp29[12],pp26[16],pp28[15]};
    CLA_4 KS_125(s125, c125, in125_1, in125_2);
    wire[3:0] s126, in126_1, in126_2;
    wire c126;
    assign in126_1 = {s49[1],pp30[11],pp27[15],pp29[14]};
    assign in126_2 = {s50[1],pp31[10],pp28[14],pp30[13]};
    CLA_4 KS_126(s126, c126, in126_1, in126_2);
    wire[3:0] s127, in127_1, in127_2;
    wire c127;
    assign in127_1 = {s51[1],s48[2],pp29[13],pp31[12]};
    assign in127_2 = {s52[1],s49[2],pp30[12],c48};
    CLA_4 KS_127(s127, c127, in127_1, in127_2);
    wire[3:0] s128, in128_1, in128_2;
    wire c128;
    assign in128_1 = {c53,s50[2],pp31[11],c49};
    assign in128_2 = {s54[1],s51[2],s48[3],c50};
    CLA_4 KS_128(s128, c128, in128_1, in128_2);
    wire[0:0] s129, in129_1, in129_2;
    wire c129;
    assign in129_1 = {c55};
    assign in129_2 = {s56[1]};
    Half_Adder KS_129(s129, c129, in129_1, in129_2);
    wire[3:0] s130, in130_1, in130_2;
    wire c130;
    assign in130_1 = {c57,c52,s49[3],c54};
    assign in130_2 = {s58[1],s54[2],s50[3],s60[0]};
    CLA_4 KS_130(s130, c130, in130_1, in130_2);
    wire[0:0] s131, in131_1, in131_2;
    wire c131;
    assign in131_1 = {c59};
    assign in131_2 = {c109};
    Half_Adder KS_131(s131, c131, in131_1, in131_2);
    wire[1:0] s132, in132_1, in132_2;
    wire c132;
    assign in132_1 = {c110,c56};
    assign in132_2 = {c111,s58[2]};
    CLA_2 KS_132(s132, c132, in132_1, in132_2);
    wire[0:0] s133, in133_1, in133_2;
    wire c133;
    assign in133_1 = {c112};
    assign in133_2 = {c113};
    Half_Adder KS_133(s133, c133, in133_1, in133_2);
    wire[2:0] s134, in134_1, in134_2;
    wire c134;
    assign in134_1 = {c114,s122[1],c51};
    assign in134_2 = {c115,s123[1],s54[3]};
    CLA_3 KS_134(s134, c134, in134_1, in134_2);
    wire[0:0] s135, in135_1, in135_2;
    wire c135;
    assign in135_1 = {s122[0]};
    assign in135_2 = {s123[0]};
    Full_Adder KS_135(s135, c135, in135_1, in135_2, c117);
    wire[3:0] s136, in136_1, in136_2;
    wire c136;
    assign in136_1 = {pp17[27],pp16[29],pp15[31],pp16[31]};
    assign in136_2 = {pp18[26],pp17[28],pp16[30],pp17[30]};
    CLA_4 KS_136(s136, c136, in136_1, in136_2);
    wire[3:0] s137, in137_1, in137_2;
    wire c137;
    assign in137_1 = {pp19[25],pp18[27],pp17[29],pp18[29]};
    assign in137_2 = {pp20[24],pp19[26],pp18[28],pp19[28]};
    CLA_4 KS_137(s137, c137, in137_1, in137_2);
    wire[3:0] s138, in138_1, in138_2;
    wire c138;
    assign in138_1 = {pp21[23],pp20[25],pp19[27],pp20[27]};
    assign in138_2 = {pp22[22],pp21[24],pp20[26],pp21[26]};
    CLA_4 KS_138(s138, c138, in138_1, in138_2);
    wire[3:0] s139, in139_1, in139_2;
    wire c139;
    assign in139_1 = {pp23[21],pp22[23],pp21[25],pp22[25]};
    assign in139_2 = {pp24[20],pp23[22],pp22[24],pp23[24]};
    CLA_4 KS_139(s139, c139, in139_1, in139_2);
    wire[3:0] s140, in140_1, in140_2;
    wire c140;
    assign in140_1 = {pp25[19],pp24[21],pp23[23],pp24[23]};
    assign in140_2 = {pp26[18],pp25[20],pp24[22],pp25[22]};
    CLA_4 KS_140(s140, c140, in140_1, in140_2);
    wire[2:0] s141, in141_1, in141_2;
    wire c141;
    assign in141_1 = {pp27[17],pp26[19],pp25[21]};
    assign in141_2 = {pp28[16],pp27[18],pp26[20]};
    CLA_3 KS_141(s141, c141, in141_1, in141_2);
    wire[3:0] s142, in142_1, in142_2;
    wire c142;
    assign in142_1 = {pp29[15],pp28[17],pp27[19],pp26[21]};
    assign in142_2 = {pp30[14],pp29[16],pp28[18],pp27[20]};
    CLA_4 KS_142(s142, c142, in142_1, in142_2);
    wire[0:0] s143, in143_1, in143_2;
    wire c143;
    assign in143_1 = {pp31[13]};
    assign in143_2 = {s60[1]};
    Half_Adder KS_143(s143, c143, in143_1, in143_2);
    wire[1:0] s144, in144_1, in144_2;
    wire c144;
    assign in144_1 = {c61,pp30[15]};
    assign in144_2 = {s62[1],pp31[14]};
    CLA_2 KS_144(s144, c144, in144_1, in144_2);
    wire[0:0] s145, in145_1, in145_2;
    wire c145;
    assign in145_1 = {c63};
    assign in145_2 = {c122};
    Half_Adder KS_145(s145, c145, in145_1, in145_2);
    wire[2:0] s146, in146_1, in146_2;
    wire c146;
    assign in146_1 = {c123,c60,pp29[17]};
    assign in146_2 = {c124,s62[2],pp30[16]};
    CLA_3 KS_146(s146, c146, in146_1, in146_2);
    wire[0:0] s147, in147_1, in147_2;
    wire c147;
    assign in147_1 = {c125};
    assign in147_2 = {c126};
    Half_Adder KS_147(s147, c147, in147_1, in147_2);
    wire[1:0] s148, in148_1, in148_2;
    wire c148;
    assign in148_1 = {c127,s136[1]};
    assign in148_2 = {c128,s137[1]};
    CLA_2 KS_148(s148, c148, in148_1, in148_2);
    wire[0:0] s149, in149_1, in149_2;
    wire c149;
    assign in149_1 = {s136[0]};
    assign in149_2 = {s137[0]};
    Full_Adder KS_149(s149, c149, in149_1, in149_2, c130);
    wire[3:0] s150, in150_1, in150_2;
    wire c150;
    assign in150_1 = {pp17[31],pp18[31],pp19[31],pp20[31]};
    assign in150_2 = {pp18[30],pp19[30],pp20[30],pp21[30]};
    CLA_4 KS_150(s150, c150, in150_1, in150_2);
    wire[2:0] s151, in151_1, in151_2;
    wire c151;
    assign in151_1 = {pp19[29],pp20[29],pp21[29]};
    assign in151_2 = {pp20[28],pp21[28],pp22[28]};
    CLA_3 KS_151(s151, c151, in151_1, in151_2);
    wire[1:0] s152, in152_1, in152_2;
    wire c152;
    assign in152_1 = {pp21[27],pp22[27]};
    assign in152_2 = {pp22[26],pp23[26]};
    CLA_2 KS_152(s152, c152, in152_1, in152_2);
    wire[0:0] s153, in153_1, in153_2;
    wire c153;
    assign in153_1 = {pp23[25]};
    assign in153_2 = {pp24[24]};
    Half_Adder KS_153(s153, c153, in153_1, in153_2);
    wire[3:0] s154, in154_1, in154_2;
    wire c154;
    assign in154_1 = {pp25[23],pp24[25],pp23[27],pp22[29]};
    assign in154_2 = {pp26[22],pp25[24],pp24[26],pp23[28]};
    CLA_4 KS_154(s154, c154, in154_1, in154_2);
    wire[0:0] s155, in155_1, in155_2;
    wire c155;
    assign in155_1 = {pp27[21]};
    assign in155_2 = {pp28[20]};
    Half_Adder KS_155(s155, c155, in155_1, in155_2);
    wire[1:0] s156, in156_1, in156_2;
    wire c156;
    assign in156_1 = {pp29[19],pp26[23]};
    assign in156_2 = {pp30[18],pp27[22]};
    CLA_2 KS_156(s156, c156, in156_1, in156_2);
    wire[0:0] s157, in157_1, in157_2;
    wire c157;
    assign in157_1 = {c136};
    assign in157_2 = {c137};
    Full_Adder KS_157(s157, c157, in157_1, in157_2, pp31[17]);
    wire[0:0] s158, in158_1, in158_2;
    wire c158;
    assign in158_1 = {pp21[31]};
    assign in158_2 = {pp22[30]};
    Half_Adder KS_158(s158, c158, in158_1, in158_2);

    /*Stage 3*/
    wire[3:0] s159, in159_1, in159_2;
    wire c159;
    assign in159_1 = {pp0[8],pp0[9],pp0[10],pp0[11]};
    assign in159_2 = {pp1[7],pp1[8],pp1[9],pp1[10]};
    CLA_4 KS_159(s159, c159, in159_1, in159_2);
    wire[3:0] s160, in160_1, in160_2;
    wire c160;
    assign in160_1 = {pp2[7],pp2[8],pp2[9],pp2[10]};
    assign in160_2 = {pp3[6],pp3[7],pp3[8],pp3[9]};
    CLA_4 KS_160(s160, c160, in160_1, in160_2);
    wire[3:0] s161, in161_1, in161_2;
    wire c161;
    assign in161_1 = {pp4[6],pp4[7],pp4[8],pp4[9]};
    assign in161_2 = {pp5[5],pp5[6],pp5[7],pp5[8]};
    CLA_4 KS_161(s161, c161, in161_1, in161_2);
    wire[3:0] s162, in162_1, in162_2;
    wire c162;
    assign in162_1 = {pp6[5],pp6[6],pp6[7],pp6[8]};
    assign in162_2 = {pp7[4],pp7[5],pp7[6],pp7[7]};
    CLA_4 KS_162(s162, c162, in162_1, in162_2);
    wire[3:0] s163, in163_1, in163_2;
    wire c163;
    assign in163_1 = {pp9[3],pp8[5],pp8[6],pp8[7]};
    assign in163_2 = {pp10[2],pp9[4],pp9[5],pp9[6]};
    CLA_4_c KS_163(s163, c163, in163_1, in163_2, pp8[4]);
    wire[3:0] s164, in164_1, in164_2;
    wire c164;
    assign in164_1 = {pp11[2],pp10[4],pp10[5],pp11[5]};
    assign in164_2 = {pp12[1],pp11[3],pp11[4],pp12[4]};
    CLA_4_c KS_164(s164, c164, in164_1, in164_2, pp10[3]);
    wire[3:0] s165, in165_1, in165_2;
    wire c165;
    assign in165_1 = {pp13[1],pp12[3],pp13[3],pp13[4]};
    assign in165_2 = {pp14[0],pp13[2],pp14[2],pp14[3]};
    CLA_4_c KS_165(s165, c165, in165_1, in165_2, pp12[2]);
    wire[3:0] s166, in166_1, in166_2;
    wire c166;
    assign in166_1 = {pp15[0],pp15[1],pp15[2],pp15[3]};
    assign in166_2 = {s64[3],pp16[0],pp16[1],pp16[2]};
    CLA_4_c KS_166(s166, c166, in166_1, in166_2, pp14[1]);
    wire[3:0] s167, in167_1, in167_2;
    wire c167;
    assign in167_1 = {s65[3],pp17[0],pp17[1],pp17[2]};
    assign in167_2 = {s66[2],c65,pp18[0],pp18[1]};
    CLA_4_c KS_167(s167, c167, in167_1, in167_2, c64);
    wire[3:0] s168, in168_1, in168_2;
    wire c168;
    assign in168_1 = {s67[2],c66,pp19[0],s1[1]};
    assign in168_2 = {s68[1],s67[3],s1[0],s2[0]};
    CLA_4_c KS_168(s168, c168, in168_1, in168_2, s66[3]);
    wire[3:0] s169, in169_1, in169_2;
    wire c169;
    assign in169_1 = {s69[2],c67,c68,s2[1]};
    assign in169_2 = {s70[1],s68[3],c69,s3[0]};
    CLA_4_c KS_169(s169, c169, in169_1, in169_2, s68[2]);
    wire[3:0] s170, in170_1, in170_2;
    wire c170;
    assign in170_1 = {s70[2],s70[3],c70,s3[1]};
    assign in170_2 = {s71[2],s71[3],c71,s4[0]};
    CLA_4_c KS_170(s170, c170, in170_1, in170_2, s69[3]);
    wire[3:0] s171, in171_1, in171_2;
    wire c171;
    assign in171_1 = {s73[2],s72[3],c72,s4[1]};
    assign in171_2 = {s74[1],s73[3],c73,s5[0]};
    CLA_4_c KS_171(s171, c171, in171_1, in171_2, s72[2]);
    wire[3:0] s172, in172_1, in172_2;
    wire c172;
    assign in172_1 = {s75[1],s74[3],s6[0],c75};
    assign in172_2 = {s76[1],s75[2],c74,c76};
    CLA_4_c KS_172(s172, c172, in172_1, in172_2, s74[2]);
    wire[3:0] s173, in173_1, in173_2;
    wire c173;
    assign in173_1 = {s77[2],s75[3],c77,s9[0]};
    assign in173_2 = {s78[1],s76[3],s78[3],s10[0]};
    CLA_4_c KS_173(s173, c173, in173_1, in173_2, s76[2]);
    wire[3:0] s174, in174_1, in174_2;
    wire c174;
    assign in174_1 = {s78[2],s79[3],c78,s11[0]};
    assign in174_2 = {s79[2],s80[2],c79,s12[0]};
    CLA_4_c KS_174(s174, c174, in174_1, in174_2, s77[3]);
    wire[3:0] s175, in175_1, in175_2;
    wire c175;
    assign in175_1 = {s82[1],s80[3],c80,s14[0]};
    assign in175_2 = {s83[0],s81[3],c81,s15[0]};
    CLA_4_c KS_175(s175, c175, in175_1, in175_2, s81[2]);
    wire[3:0] s176, in176_1, in176_2;
    wire c176;
    assign in176_1 = {s83[1],s82[3],s16[0],c85};
    assign in176_2 = {s84[1],s83[2],c82,c86};
    CLA_4_c KS_176(s176, c176, in176_1, in176_2, s82[2]);
    wire[3:0] s177, in177_1, in177_2;
    wire c177;
    assign in177_1 = {s85[2],s83[3],s87[3],s22[0]};
    assign in177_2 = {s86[2],s84[3],s88[2],c87};
    CLA_4_c KS_177(s177, c177, in177_1, in177_2, s84[2]);
    wire[3:0] s178, in178_1, in178_2;
    wire c178;
    assign in178_1 = {s86[3],s89[2],s88[3],s24[0]};
    assign in178_2 = {s87[2],s90[1],s89[3],s25[0]};
    CLA_4_c KS_178(s178, c178, in178_1, in178_2, s85[3]);
    wire[3:0] s179, in179_1, in179_2;
    wire c179;
    assign in179_1 = {s92[0],s90[2],c88,s30[0]};
    assign in179_2 = {s93[0],s91[1],c89,s31[0]};
    CLA_4_c KS_179(s179, c179, in179_1, in179_2, s91[0]);
    wire[3:0] s180, in180_1, in180_2;
    wire c180;
    assign in180_1 = {s92[1],s90[3],s32[0],s97[2]};
    assign in180_2 = {s93[1],s91[2],c90,s98[1]};
    CLA_4 KS_180(s180, c180, in180_1, in180_2);
    wire[3:0] s181, in181_1, in181_2;
    wire c181;
    assign in181_1 = {s93[2],s91[3],s99[0],s98[2]};
    assign in181_2 = {s94[2],s92[3],s100[0],s99[1]};
    CLA_4_c KS_181(s181, c181, in181_1, in181_2, s92[2]);
    wire[3:0] s182, in182_1, in182_2;
    wire c182;
    assign in182_1 = {s94[3],s101[0],s100[1],s37[0]};
    assign in182_2 = {s95[3],s102[0],s101[1],c97};
    CLA_4_c KS_182(s182, c182, in182_1, in182_2, s93[3]);
    wire[3:0] s183, in183_1, in183_2;
    wire c183;
    assign in183_1 = {s104[0],s102[1],s98[3],s45[0]};
    assign in183_2 = {s105[0],s103[1],s99[2],s46[0]};
    CLA_4_c KS_183(s183, c183, in183_1, in183_2, s103[0]);
    wire[3:0] s184, in184_1, in184_2;
    wire c184;
    assign in184_1 = {s104[1],s100[2],s47[0],s110[0]};
    assign in184_2 = {c105,s101[2],c98,s111[0]};
    CLA_4 KS_184(s184, c184, in184_1, in184_2);
    wire[3:0] s185, in185_1, in185_2;
    wire c185;
    assign in185_1 = {s102[2],s99[3],s112[0],s111[1]};
    assign in185_2 = {s103[2],s100[3],s113[0],s112[1]};
    CLA_4 KS_185(s185, c185, in185_1, in185_2);
    wire[3:0] s186, in186_1, in186_2;
    wire c186;
    assign in186_1 = {s102[3],s114[0],s113[1],s47[3]};
    assign in186_2 = {s103[3],s115[0],s114[1],s109[2]};
    CLA_4_c KS_186(s186, c186, in186_1, in186_2, s101[3]);
    wire[3:0] s187, in187_1, in187_2;
    wire c187;
    assign in187_1 = {s117[0],s115[1],s110[2],s57[0]};
    assign in187_2 = {s118[0],c116,s111[2],s58[0]};
    CLA_4_c KS_187(s187, c187, in187_1, in187_2, s116[0]);
    wire[3:0] s188, in188_1, in188_2;
    wire c188;
    assign in188_1 = {s117[1],s112[2],s59[0],s124[0]};
    assign in188_2 = {c118,s113[2],s109[3],s125[0]};
    CLA_4 KS_188(s188, c188, in188_1, in188_2);
    wire[3:0] s189, in189_1, in189_2;
    wire c189;
    assign in189_1 = {s114[2],s110[3],s126[0],s124[1]};
    assign in189_2 = {s115[2],s111[3],s127[0],s125[1]};
    CLA_4 KS_189(s189, c189, in189_1, in189_2);
    wire[3:0] s190, in190_1, in190_2;
    wire c190;
    assign in190_1 = {s113[3],s128[0],s126[1],c58};
    assign in190_2 = {s114[3],s129[0],s127[1],s122[2]};
    CLA_4_c KS_190(s190, c190, in190_1, in190_2, s112[3]);
    wire[3:0] s191, in191_1, in191_2;
    wire c191;
    assign in191_1 = {s131[0],s128[1],s123[2],s61[0]};
    assign in191_2 = {s132[0],c129,s124[2],s62[0]};
    CLA_4_c KS_191(s191, c191, in191_1, in191_2, s130[0]);
    wire[3:0] s192, in192_1, in192_2;
    wire c192;
    assign in192_1 = {c131,s125[2],s63[0],s138[0]};
    assign in192_2 = {s132[1],s126[2],s122[3],s139[0]};
    CLA_4_c KS_192(s192, c192, in192_1, in192_2, s130[1]);
    wire[3:0] s193, in193_1, in193_2;
    wire c193;
    assign in193_1 = {s127[2],s123[3],s140[0],s138[1]};
    assign in193_2 = {s128[2],s124[3],s141[0],s139[1]};
    CLA_4 KS_193(s193, c193, in193_1, in193_2);
    wire[3:0] s194, in194_1, in194_2;
    wire c194;
    assign in194_1 = {s126[3],s142[0],s140[1],pp31[15]};
    assign in194_2 = {s127[3],s143[0],s141[1],c62};
    CLA_4_c KS_194(s194, c194, in194_1, in194_2, s125[3]);
    wire[3:0] s195, in195_1, in195_2;
    wire c195;
    assign in195_1 = {s145[0],s142[1],s136[2],pp28[19]};
    assign in195_2 = {s146[0],c143,s137[2],pp29[18]};
    CLA_4_c KS_195(s195, c195, in195_1, in195_2, s144[0]);
    wire[3:0] s196, in196_1, in196_2;
    wire c196;
    assign in196_1 = {c145,s138[2],pp30[17],c138};
    assign in196_2 = {s146[1],s139[2],pp31[16],c139};
    CLA_4_c KS_196(s196, c196, in196_1, in196_2, s144[1]);
    wire[3:0] s197, in197_1, in197_2;
    wire c197;
    assign in197_1 = {s141[2],s136[3],c140,pp28[21]};
    assign in197_2 = {s142[2],s137[3],c142,pp29[20]};
    CLA_4_c KS_197(s197, c197, in197_1, in197_2, s140[2]);
    wire[3:0] s198, in198_1, in198_2;
    wire c198;
    assign in198_1 = {s139[3],s150[0],pp30[19],pp25[25]};
    assign in198_2 = {s140[3],s151[0],pp31[18],pp26[24]};
    CLA_4_c KS_198(s198, c198, in198_1, in198_2, s138[3]);
    wire[3:0] s199, in199_1, in199_2;
    wire c199;
    assign in199_1 = {s153[0],s150[1],pp27[23],pp24[27]};
    assign in199_2 = {s154[0],s151[1],pp28[22],pp25[26]};
    CLA_4_c KS_199(s199, c199, in199_1, in199_2, s152[0]);
    wire[3:0] s200, in200_1, in200_2;
    wire c200;
    assign in200_1 = {c153,pp29[21],pp26[25],pp23[29]};
    assign in200_2 = {s154[1],pp30[20],pp27[24],pp24[28]};
    CLA_4_c KS_200(s200, c200, in200_1, in200_2, s152[1]);
    wire[3:0] s201, in201_1, in201_2;
    wire c201;
    assign in201_1 = {s150[2],pp28[23],pp25[27],pp22[31]};
    assign in201_2 = {s151[2],pp29[22],pp26[26],pp23[30]};
    CLA_4_c KS_201(s201, c201, in201_1, in201_2, pp31[19]);
    wire[3:0] s202, in202_1, in202_2;
    wire c202;
    assign in202_1 = {pp30[21],pp27[25],pp24[29],pp23[31]};
    assign in202_2 = {pp31[20],pp28[24],pp25[28],pp24[30]};
    CLA_4 KS_202(s202, c202, in202_1, in202_2);
    wire[3:0] s203, in203_1, in203_2;
    wire c203;
    assign in203_1 = {pp30[22],pp26[27],pp25[29],pp24[31]};
    assign in203_2 = {pp31[21],pp27[26],pp26[28],pp25[30]};
    CLA_4_c KS_203(s203, c203, in203_1, in203_2, pp29[23]);
    wire[3:0] s204, in204_1, in204_2;
    wire c204;
    assign in204_1 = {pp28[25],pp27[27],pp26[29],pp25[31]};
    assign in204_2 = {pp29[24],pp28[26],pp27[28],pp26[30]};
    CLA_4 KS_204(s204, c204, in204_1, in204_2);

    /*Stage 4*/
    wire[3:0] s205, in205_1, in205_2;
    wire c205;
    assign in205_1 = {pp0[5],pp0[6],pp0[7],pp2[6]};
    assign in205_2 = {pp1[4],pp1[5],pp1[6],pp3[5]};
    CLA_4 KS_205(s205, c205, in205_1, in205_2);
    wire[3:0] s206, in206_1, in206_2;
    wire c206;
    assign in206_1 = {pp2[4],pp2[5],pp4[4],pp4[5]};
    assign in206_2 = {pp3[3],pp3[4],pp5[3],pp5[4]};
    CLA_4 KS_206(s206, c206, in206_1, in206_2);
    wire[3:0] s207, in207_1, in207_2;
    wire c207;
    assign in207_1 = {pp4[3],pp6[2],pp6[3],pp6[4]};
    assign in207_2 = {pp5[2],pp7[1],pp7[2],pp7[3]};
    CLA_4 KS_207(s207, c207, in207_1, in207_2);
    wire[3:0] s208, in208_1, in208_2;
    wire c208;
    assign in208_1 = {pp9[0],pp8[2],pp8[3],pp11[1]};
    assign in208_2 = {s159[1],pp9[1],pp9[2],pp12[0]};
    CLA_4_c KS_208(s208, c208, in208_1, in208_2, pp8[1]);
    wire[3:0] s209, in209_1, in209_2;
    wire c209;
    assign in209_1 = {s159[2],pp10[1],s64[0],pp13[0]};
    assign in209_2 = {s160[1],pp11[0],c159,s64[1]};
    CLA_4_c KS_209(s209, c209, in209_1, in209_2, pp10[0]);
    wire[3:0] s210, in210_1, in210_2;
    wire c210;
    assign in210_1 = {s160[2],s160[3],s65[0],s64[2]};
    assign in210_2 = {s161[1],s161[2],c160,s65[1]};
    CLA_4_c KS_210(s210, c210, in210_1, in210_2, s159[3]);
    wire[3:0] s211, in211_1, in211_2;
    wire c211;
    assign in211_1 = {s162[2],s66[0],s65[2],s67[1]};
    assign in211_2 = {s163[1],c161,s66[1],s68[0]};
    CLA_4_c KS_211(s211, c211, in211_1, in211_2, s161[3]);
    wire[3:0] s212, in212_1, in212_2;
    wire c212;
    assign in212_1 = {s163[2],s67[0],s69[0],s69[1]};
    assign in212_2 = {s164[1],c162,c163,s70[0]};
    CLA_4_c KS_212(s212, c212, in212_1, in212_2, s162[3]);
    wire[3:0] s213, in213_1, in213_2;
    wire c213;
    assign in213_1 = {s164[2],s164[3],s71[0],s71[1]};
    assign in213_2 = {s165[1],s165[2],c164,s72[0]};
    CLA_4_c KS_213(s213, c213, in213_1, in213_2, s163[3]);
    wire[3:0] s214, in214_1, in214_2;
    wire c214;
    assign in214_1 = {s166[2],s73[0],s72[1],s75[0]};
    assign in214_2 = {s167[1],c165,s73[1],s76[0]};
    CLA_4_c KS_214(s214, c214, in214_1, in214_2, s165[3]);
    wire[3:0] s215, in215_1, in215_2;
    wire c215;
    assign in215_1 = {s167[2],s74[0],s77[0],s77[1]};
    assign in215_2 = {s168[1],c166,c167,s78[0]};
    CLA_4_c KS_215(s215, c215, in215_1, in215_2, s166[3]);
    wire[3:0] s216, in216_1, in216_2;
    wire c216;
    assign in216_1 = {s168[2],s168[3],s79[0],s79[1]};
    assign in216_2 = {s169[1],s169[2],c168,s80[0]};
    CLA_4_c KS_216(s216, c216, in216_1, in216_2, s167[3]);
    wire[3:0] s217, in217_1, in217_2;
    wire c217;
    assign in217_1 = {s170[2],s81[0],s80[1],s84[0]};
    assign in217_2 = {s171[1],c169,s81[1],s85[0]};
    CLA_4_c KS_217(s217, c217, in217_1, in217_2, s169[3]);
    wire[3:0] s218, in218_1, in218_2;
    wire c218;
    assign in218_1 = {s171[2],s82[0],s86[0],s85[1]};
    assign in218_2 = {s172[1],c170,c171,s86[1]};
    CLA_4_c KS_218(s218, c218, in218_1, in218_2, s170[3]);
    wire[3:0] s219, in219_1, in219_2;
    wire c219;
    assign in219_1 = {s172[2],s172[3],s87[0],s87[1]};
    assign in219_2 = {s173[1],s173[2],c172,s88[0]};
    CLA_4_c KS_219(s219, c219, in219_1, in219_2, s171[3]);
    wire[3:0] s220, in220_1, in220_2;
    wire c220;
    assign in220_1 = {s174[2],s89[0],s88[1],s94[0]};
    assign in220_2 = {s175[1],c173,s89[1],s95[0]};
    CLA_4_c KS_220(s220, c220, in220_1, in220_2, s173[3]);
    wire[3:0] s221, in221_1, in221_2;
    wire c221;
    assign in221_1 = {s175[2],s90[0],s96[0],s94[1]};
    assign in221_2 = {s176[1],c174,c175,s95[1]};
    CLA_4_c KS_221(s221, c221, in221_1, in221_2, s174[3]);
    wire[3:0] s222, in222_1, in222_2;
    wire c222;
    assign in222_1 = {s176[2],s176[3],s96[1],s95[2]};
    assign in222_2 = {s177[1],s177[2],c176,s96[2]};
    CLA_4_c KS_222(s222, c222, in222_1, in222_2, s175[3]);
    wire[3:0] s223, in223_1, in223_2;
    wire c223;
    assign in223_1 = {s178[2],s97[0],s96[3],s106[0]};
    assign in223_2 = {s179[1],c177,s97[1],s107[0]};
    CLA_4_c KS_223(s223, c223, in223_1, in223_2, s177[3]);
    wire[3:0] s224, in224_1, in224_2;
    wire c224;
    assign in224_1 = {s179[2],s98[0],s108[0],s106[1]};
    assign in224_2 = {s180[1],c178,c179,c107};
    CLA_4_c KS_224(s224, c224, in224_1, in224_2, s178[3]);
    wire[3:0] s225, in225_1, in225_2;
    wire c225;
    assign in225_1 = {s180[2],s180[3],s108[1],s104[2]};
    assign in225_2 = {s181[1],s181[2],c180,s106[2]};
    CLA_4_c KS_225(s225, c225, in225_1, in225_2, s179[3]);
    wire[3:0] s226, in226_1, in226_2;
    wire c226;
    assign in226_1 = {s182[2],s108[2],s104[3],s119[0]};
    assign in226_2 = {s183[1],c181,s106[3],s120[0]};
    CLA_4_c KS_226(s226, c226, in226_1, in226_2, s181[3]);
    wire[3:0] s227, in227_1, in227_2;
    wire c227;
    assign in227_1 = {s183[2],s108[3],s121[0],s119[1]};
    assign in227_2 = {s184[1],c182,c183,c120};
    CLA_4_c KS_227(s227, c227, in227_1, in227_2, s182[3]);
    wire[3:0] s228, in228_1, in228_2;
    wire c228;
    assign in228_1 = {s184[2],s184[3],s121[1],s117[2]};
    assign in228_2 = {s185[1],s185[2],c184,c119};
    CLA_4_c KS_228(s228, c228, in228_1, in228_2, s183[3]);
    wire[3:0] s229, in229_1, in229_2;
    wire c229;
    assign in229_1 = {s186[2],s121[2],s115[3],s133[0]};
    assign in229_2 = {s187[1],c185,s117[3],s134[0]};
    CLA_4_c KS_229(s229, c229, in229_1, in229_2, s185[3]);
    wire[3:0] s230, in230_1, in230_2;
    wire c230;
    assign in230_1 = {s187[2],c121,s135[0],c133};
    assign in230_2 = {s188[1],c186,c187,s134[1]};
    CLA_4_c KS_230(s230, c230, in230_1, in230_2, s186[3]);
    wire[3:0] s231, in231_1, in231_2;
    wire c231;
    assign in231_1 = {s188[2],s188[3],c135,s130[2]};
    assign in231_2 = {s189[1],s189[2],c188,c132};
    CLA_4_c KS_231(s231, c231, in231_1, in231_2, s187[3]);
    wire[3:0] s232, in232_1, in232_2;
    wire c232;
    assign in232_1 = {s190[2],s134[2],s128[3],s147[0]};
    assign in232_2 = {s191[1],c189,s130[3],s148[0]};
    CLA_4_c KS_232(s232, c232, in232_1, in232_2, s189[3]);
    wire[3:0] s233, in233_1, in233_2;
    wire c233;
    assign in233_1 = {s191[2],c134,s149[0],c147};
    assign in233_2 = {s192[1],c190,c191,s148[1]};
    CLA_4_c KS_233(s233, c233, in233_1, in233_2, s190[3]);
    wire[3:0] s234, in234_1, in234_2;
    wire c234;
    assign in234_1 = {s192[2],s192[3],c149,c144};
    assign in234_2 = {s193[1],s193[2],c192,s146[2]};
    CLA_4_c KS_234(s234, c234, in234_1, in234_2, s191[3]);
    wire[3:0] s235, in235_1, in235_2;
    wire c235;
    assign in235_1 = {s194[2],c148,c141,s155[0]};
    assign in235_2 = {s195[1],c193,s142[3],s156[0]};
    CLA_4_c KS_235(s235, c235, in235_1, in235_2, s193[3]);
    wire[3:0] s236, in236_1, in236_2;
    wire c236;
    assign in236_1 = {s195[2],c146,s157[0],c155};
    assign in236_2 = {s196[1],c194,c195,s156[1]};
    CLA_4_c KS_236(s236, c236, in236_1, in236_2, s194[3]);
    wire[3:0] s237, in237_1, in237_2;
    wire c237;
    assign in237_1 = {s196[2],s196[3],c157,c152};
    assign in237_2 = {s197[1],s197[2],c196,s154[2]};
    CLA_4_c KS_237(s237, c237, in237_1, in237_2, s195[3]);
    wire[3:0] s238, in238_1, in238_2;
    wire c238;
    assign in238_1 = {s198[2],c156,s150[3],c150};
    assign in238_2 = {s199[1],c197,c151,c154};
    CLA_4_c KS_238(s238, c238, in238_1, in238_2, s197[3]);
    wire[3:0] s239, in239_1, in239_2;
    wire c239;
    assign in239_1 = {s199[2],s154[3],s158[0],pp30[23]};
    assign in239_2 = {s200[1],c198,c199,pp31[22]};
    CLA_4_c KS_239(s239, c239, in239_1, in239_2, s198[3]);
    wire[3:0] s240, in240_1, in240_2;
    wire c240;
    assign in240_1 = {s200[2],s200[3],c158,pp29[25]};
    assign in240_2 = {s201[1],s201[2],c200,pp30[24]};
    CLA_4_c KS_240(s240, c240, in240_1, in240_2, s199[3]);
    wire[3:0] s241, in241_1, in241_2;
    wire c241;
    assign in241_1 = {s202[2],pp31[23],pp28[27],pp27[29]};
    assign in241_2 = {s203[1],c201,pp29[26],pp28[28]};
    CLA_4_c KS_241(s241, c241, in241_1, in241_2, s201[3]);
    wire[3:0] s242, in242_1, in242_2;
    wire c242;
    assign in242_1 = {s202[3],pp30[25],pp29[27],pp26[31]};
    assign in242_2 = {s203[2],pp31[24],pp30[26],pp27[30]};
    CLA_4 KS_242(s242, c242, in242_1, in242_2);
    wire[3:0] s243, in243_1, in243_2;
    wire c243;
    assign in243_1 = {c202,pp31[25],pp28[29],pp27[31]};
    assign in243_2 = {s203[3],c203,pp29[28],pp28[30]};
    CLA_4 KS_243(s243, c243, in243_1, in243_2);
    wire[2:0] s244, in244_1, in244_2;
    wire c244;
    assign in244_1 = {pp30[27],pp29[29],pp28[31]};
    assign in244_2 = {pp31[26],pp30[28],pp29[30]};
    CLA_3 KS_244(s244, c244, in244_1, in244_2);

    /*Stage 5*/
    wire[3:0] s245, in245_1, in245_2;
    wire c245;
    assign in245_1 = {pp0[3],pp0[4],pp2[3],pp4[2]};
    assign in245_2 = {pp1[2],pp1[3],pp3[2],pp5[1]};
    CLA_4 KS_245(s245, c245, in245_1, in245_2);
    wire[3:0] s246, in246_1, in246_2;
    wire c246;
    assign in246_1 = {pp2[2],pp4[1],pp6[0],pp6[1]};
    assign in246_2 = {pp3[1],pp5[0],s205[1],pp7[0]};
    CLA_4 KS_246(s246, c246, in246_1, in246_2);
    wire[3:0] s247, in247_1, in247_2;
    wire c247;
    assign in247_1 = {s206[1],pp8[0],s160[0],s161[0]};
    assign in247_2 = {s207[0],s159[0],c205,c206};
    CLA_4_c KS_247(s247, c247, in247_1, in247_2, s205[2]);
    wire[3:0] s248, in248_1, in248_2;
    wire c248;
    assign in248_1 = {s206[2],s206[3],s207[3],s162[0]};
    assign in248_2 = {s207[1],s207[2],s208[1],c207};
    CLA_4_c KS_248(s248, c248, in248_1, in248_2, s205[3]);
    wire[3:0] s249, in249_1, in249_2;
    wire c249;
    assign in249_1 = {s209[1],s162[1],s164[0],s165[0]};
    assign in249_2 = {s210[0],s163[0],c208,c209};
    CLA_4_c KS_249(s249, c249, in249_1, in249_2, s208[2]);
    wire[3:0] s250, in250_1, in250_2;
    wire c250;
    assign in250_1 = {s209[2],s209[3],s210[3],s166[0]};
    assign in250_2 = {s210[1],s210[2],s211[1],c210};
    CLA_4_c KS_250(s250, c250, in250_1, in250_2, s208[3]);
    wire[3:0] s251, in251_1, in251_2;
    wire c251;
    assign in251_1 = {s212[1],s166[1],s168[0],s169[0]};
    assign in251_2 = {s213[0],s167[0],c211,c212};
    CLA_4_c KS_251(s251, c251, in251_1, in251_2, s211[2]);
    wire[3:0] s252, in252_1, in252_2;
    wire c252;
    assign in252_1 = {s212[2],s212[3],s213[3],s170[0]};
    assign in252_2 = {s213[1],s213[2],s214[1],c213};
    CLA_4_c KS_252(s252, c252, in252_1, in252_2, s211[3]);
    wire[3:0] s253, in253_1, in253_2;
    wire c253;
    assign in253_1 = {s215[1],s170[1],s172[0],s173[0]};
    assign in253_2 = {s216[0],s171[0],c214,c215};
    CLA_4_c KS_253(s253, c253, in253_1, in253_2, s214[2]);
    wire[3:0] s254, in254_1, in254_2;
    wire c254;
    assign in254_1 = {s215[2],s215[3],s216[3],s174[0]};
    assign in254_2 = {s216[1],s216[2],s217[1],c216};
    CLA_4_c KS_254(s254, c254, in254_1, in254_2, s214[3]);
    wire[3:0] s255, in255_1, in255_2;
    wire c255;
    assign in255_1 = {s218[1],s174[1],s176[0],s177[0]};
    assign in255_2 = {s219[0],s175[0],c217,c218};
    CLA_4_c KS_255(s255, c255, in255_1, in255_2, s217[2]);
    wire[3:0] s256, in256_1, in256_2;
    wire c256;
    assign in256_1 = {s218[2],s218[3],s219[3],s178[0]};
    assign in256_2 = {s219[1],s219[2],s220[1],c219};
    CLA_4_c KS_256(s256, c256, in256_1, in256_2, s217[3]);
    wire[3:0] s257, in257_1, in257_2;
    wire c257;
    assign in257_1 = {s221[1],s178[1],s180[0],s181[0]};
    assign in257_2 = {s222[0],s179[0],c220,c221};
    CLA_4_c KS_257(s257, c257, in257_1, in257_2, s220[2]);
    wire[3:0] s258, in258_1, in258_2;
    wire c258;
    assign in258_1 = {s221[2],s221[3],s222[3],s182[0]};
    assign in258_2 = {s222[1],s222[2],s223[1],c222};
    CLA_4_c KS_258(s258, c258, in258_1, in258_2, s220[3]);
    wire[3:0] s259, in259_1, in259_2;
    wire c259;
    assign in259_1 = {s224[1],s182[1],s184[0],s185[0]};
    assign in259_2 = {s225[0],s183[0],c223,c224};
    CLA_4_c KS_259(s259, c259, in259_1, in259_2, s223[2]);
    wire[3:0] s260, in260_1, in260_2;
    wire c260;
    assign in260_1 = {s224[2],s224[3],s225[3],s186[0]};
    assign in260_2 = {s225[1],s225[2],s226[1],c225};
    CLA_4_c KS_260(s260, c260, in260_1, in260_2, s223[3]);
    wire[3:0] s261, in261_1, in261_2;
    wire c261;
    assign in261_1 = {s227[1],s186[1],s188[0],s189[0]};
    assign in261_2 = {s228[0],s187[0],c226,c227};
    CLA_4_c KS_261(s261, c261, in261_1, in261_2, s226[2]);
    wire[3:0] s262, in262_1, in262_2;
    wire c262;
    assign in262_1 = {s227[2],s227[3],s228[3],s190[0]};
    assign in262_2 = {s228[1],s228[2],s229[1],c228};
    CLA_4_c KS_262(s262, c262, in262_1, in262_2, s226[3]);
    wire[3:0] s263, in263_1, in263_2;
    wire c263;
    assign in263_1 = {s230[1],s190[1],s192[0],s193[0]};
    assign in263_2 = {s231[0],s191[0],c229,c230};
    CLA_4_c KS_263(s263, c263, in263_1, in263_2, s229[2]);
    wire[3:0] s264, in264_1, in264_2;
    wire c264;
    assign in264_1 = {s230[2],s230[3],s231[3],s194[0]};
    assign in264_2 = {s231[1],s231[2],s232[1],c231};
    CLA_4_c KS_264(s264, c264, in264_1, in264_2, s229[3]);
    wire[3:0] s265, in265_1, in265_2;
    wire c265;
    assign in265_1 = {s233[1],s194[1],s196[0],s197[0]};
    assign in265_2 = {s234[0],s195[0],c232,c233};
    CLA_4_c KS_265(s265, c265, in265_1, in265_2, s232[2]);
    wire[3:0] s266, in266_1, in266_2;
    wire c266;
    assign in266_1 = {s233[2],s233[3],s234[3],s198[0]};
    assign in266_2 = {s234[1],s234[2],s235[1],c234};
    CLA_4_c KS_266(s266, c266, in266_1, in266_2, s232[3]);
    wire[3:0] s267, in267_1, in267_2;
    wire c267;
    assign in267_1 = {s236[1],s198[1],s200[0],s201[0]};
    assign in267_2 = {s237[0],s199[0],c235,c236};
    CLA_4_c KS_267(s267, c267, in267_1, in267_2, s235[2]);
    wire[3:0] s268, in268_1, in268_2;
    wire c268;
    assign in268_1 = {s236[2],s236[3],s237[3],s202[0]};
    assign in268_2 = {s237[1],s237[2],s238[1],c237};
    CLA_4_c KS_268(s268, c268, in268_1, in268_2, s235[3]);
    wire[3:0] s269, in269_1, in269_2;
    wire c269;
    assign in269_1 = {s239[1],s202[1],s204[0],s204[1]};
    assign in269_2 = {s240[0],s203[0],c238,c239};
    CLA_4_c KS_269(s269, c269, in269_1, in269_2, s238[2]);
    wire[3:0] s270, in270_1, in270_2;
    wire c270;
    assign in270_1 = {s239[2],s239[3],s240[3],s204[2]};
    assign in270_2 = {s240[1],s240[2],s241[1],c240};
    CLA_4_c KS_270(s270, c270, in270_1, in270_2, s238[3]);
    wire[3:0] s271, in271_1, in271_2;
    wire c271;
    assign in271_1 = {s242[1],s204[3],c204,pp31[27]};
    assign in271_2 = {s243[0],s241[3],c241,c242};
    CLA_4_c KS_271(s271, c271, in271_1, in271_2, s241[2]);
    wire[3:0] s272, in272_1, in272_2;
    wire c272;
    assign in272_1 = {s242[2],s242[3],s243[3],pp30[29]};
    assign in272_2 = {s243[1],s243[2],s244[1],pp31[28]};
    CLA_4 KS_272(s272, c272, in272_1, in272_2);
    wire[1:0] s273, in273_1, in273_2;
    wire c273;
    assign in273_1 = {c243,pp29[31]};
    assign in273_2 = {s244[2],pp30[30]};
    CLA_2 KS_273(s273, c273, in273_1, in273_2);
    wire[1:0] s274, in274_1, in274_2;
    wire c274;
    assign in274_1 = {pp31[29],pp30[31]};
    assign in274_2 = {c244,pp31[30]};
    CLA_2 KS_274(s274, c274, in274_1, in274_2);

    /*Stage 6*/
    wire[3:0] s275, in275_1, in275_2;
    wire c275;
    assign in275_1 = {pp0[2],pp2[1],pp4[0],s205[0]};
    assign in275_2 = {pp1[1],pp3[0],s245[1],s245[2]};
    CLA_4 KS_275(s275, c275, in275_1, in275_2);
    wire[3:0] s276, in276_1, in276_2;
    wire c276;
    assign in276_1 = {s245[3],c245,c246,s208[0]};
    assign in276_2 = {s246[2],s246[3],s247[1],s247[2]};
    CLA_4_c KS_276(s276, c276, in276_1, in276_2, s206[0]);
    wire[3:0] s277, in277_1, in277_2;
    wire c277;
    assign in277_1 = {s247[3],c247,c248,s211[0]};
    assign in277_2 = {s248[2],s248[3],s249[1],s249[2]};
    CLA_4_c KS_277(s277, c277, in277_1, in277_2, s209[0]);
    wire[3:0] s278, in278_1, in278_2;
    wire c278;
    assign in278_1 = {s249[3],c249,c250,s214[0]};
    assign in278_2 = {s250[2],s250[3],s251[1],s251[2]};
    CLA_4_c KS_278(s278, c278, in278_1, in278_2, s212[0]);
    wire[3:0] s279, in279_1, in279_2;
    wire c279;
    assign in279_1 = {s251[3],c251,c252,s217[0]};
    assign in279_2 = {s252[2],s252[3],s253[1],s253[2]};
    CLA_4_c KS_279(s279, c279, in279_1, in279_2, s215[0]);
    wire[3:0] s280, in280_1, in280_2;
    wire c280;
    assign in280_1 = {s253[3],c253,c254,s220[0]};
    assign in280_2 = {s254[2],s254[3],s255[1],s255[2]};
    CLA_4_c KS_280(s280, c280, in280_1, in280_2, s218[0]);
    wire[3:0] s281, in281_1, in281_2;
    wire c281;
    assign in281_1 = {s255[3],c255,c256,s223[0]};
    assign in281_2 = {s256[2],s256[3],s257[1],s257[2]};
    CLA_4_c KS_281(s281, c281, in281_1, in281_2, s221[0]);
    wire[3:0] s282, in282_1, in282_2;
    wire c282;
    assign in282_1 = {s257[3],c257,c258,s226[0]};
    assign in282_2 = {s258[2],s258[3],s259[1],s259[2]};
    CLA_4_c KS_282(s282, c282, in282_1, in282_2, s224[0]);
    wire[3:0] s283, in283_1, in283_2;
    wire c283;
    assign in283_1 = {s259[3],c259,c260,s229[0]};
    assign in283_2 = {s260[2],s260[3],s261[1],s261[2]};
    CLA_4_c KS_283(s283, c283, in283_1, in283_2, s227[0]);
    wire[3:0] s284, in284_1, in284_2;
    wire c284;
    assign in284_1 = {s261[3],c261,c262,s232[0]};
    assign in284_2 = {s262[2],s262[3],s263[1],s263[2]};
    CLA_4_c KS_284(s284, c284, in284_1, in284_2, s230[0]);
    wire[3:0] s285, in285_1, in285_2;
    wire c285;
    assign in285_1 = {s263[3],c263,c264,s235[0]};
    assign in285_2 = {s264[2],s264[3],s265[1],s265[2]};
    CLA_4_c KS_285(s285, c285, in285_1, in285_2, s233[0]);
    wire[3:0] s286, in286_1, in286_2;
    wire c286;
    assign in286_1 = {s265[3],c265,c266,s238[0]};
    assign in286_2 = {s266[2],s266[3],s267[1],s267[2]};
    CLA_4_c KS_286(s286, c286, in286_1, in286_2, s236[0]);
    wire[3:0] s287, in287_1, in287_2;
    wire c287;
    assign in287_1 = {s267[3],c267,c268,s241[0]};
    assign in287_2 = {s268[2],s268[3],s269[1],s269[2]};
    CLA_4_c KS_287(s287, c287, in287_1, in287_2, s239[0]);
    wire[3:0] s288, in288_1, in288_2;
    wire c288;
    assign in288_1 = {s269[3],c269,c270,s244[0]};
    assign in288_2 = {s270[2],s270[3],s271[1],s271[2]};
    CLA_4_c KS_288(s288, c288, in288_1, in288_2, s242[0]);
    wire[3:0] s289, in289_1, in289_2;
    wire c289;
    assign in289_1 = {s271[3],c271,c272,c273};
    assign in289_2 = {s272[2],s272[3],s273[1],s274[1]};
    CLA_4 KS_289(s289, c289, in289_1, in289_2);


    /*Final Stage 6*/
    wire[61:0] s, in_1, in_2;
    wire c;
    assign in_1 = {pp0[1],pp2[0],s245[0],s246[0],s246[1],c275,s247[0],s248[0],s248[1],c276,s249[0],s250[0],s250[1],c277,s251[0],s252[0],s252[1],c278,s253[0],s254[0],s254[1],c279,s255[0],s256[0],s256[1],c280,s257[0],s258[0],s258[1],c281,s259[0],s260[0],s260[1],c282,s261[0],s262[0],s262[1],c283,s263[0],s264[0],s264[1],c284,s265[0],s266[0],s266[1],c285,s267[0],s268[0],s268[1],c286,s269[0],s270[0],s270[1],c287,s271[0],s272[0],s272[1],c288,s273[0],s274[0],s289[3],c289};
    assign in_2 = {pp1[0],s275[0],s275[1],s275[2],s275[3],s276[0],s276[1],s276[2],s276[3],s277[0],s277[1],s277[2],s277[3],s278[0],s278[1],s278[2],s278[3],s279[0],s279[1],s279[2],s279[3],s280[0],s280[1],s280[2],s280[3],s281[0],s281[1],s281[2],s281[3],s282[0],s282[1],s282[2],s282[3],s283[0],s283[1],s283[2],s283[3],s284[0],s284[1],s284[2],s284[3],s285[0],s285[1],s285[2],s285[3],s286[0],s286[1],s286[2],s286[3],s287[0],s287[1],s287[2],s287[3],s288[0],s288[1],s288[2],s288[3],s289[0],s289[1],s289[2],1'b0,1'b0};
    kogge_stone_62(s, c, in_1, in_2);

    assign product[0] = pp0[0];
    assign product[1] = s[0];
    assign product[2] = s[1];
    assign product[3] = s[2];
    assign product[4] = s[3];
    assign product[5] = s[4];
    assign product[6] = s[5];
    assign product[7] = s[6];
    assign product[8] = s[7];
    assign product[9] = s[8];
    assign product[10] = s[9];
    assign product[11] = s[10];
    assign product[12] = s[11];
    assign product[13] = s[12];
    assign product[14] = s[13];
    assign product[15] = s[14];
    assign product[16] = s[15];
    assign product[17] = s[16];
    assign product[18] = s[17];
    assign product[19] = s[18];
    assign product[20] = s[19];
    assign product[21] = s[20];
    assign product[22] = s[21];
    assign product[23] = s[22];
    assign product[24] = s[23];
    assign product[25] = s[24];
    assign product[26] = s[25];
    assign product[27] = s[26];
    assign product[28] = s[27];
    assign product[29] = s[28];
    assign product[30] = s[29];
    assign product[31] = s[30];
    assign product[32] = s[31];
    assign product[33] = s[32];
    assign product[34] = s[33];
    assign product[35] = s[34];
    assign product[36] = s[35];
    assign product[37] = s[36];
    assign product[38] = s[37];
    assign product[39] = s[38];
    assign product[40] = s[39];
    assign product[41] = s[40];
    assign product[42] = s[41];
    assign product[43] = s[42];
    assign product[44] = s[43];
    assign product[45] = s[44];
    assign product[46] = s[45];
    assign product[47] = s[46];
    assign product[48] = s[47];
    assign product[49] = s[48];
    assign product[50] = s[49];
    assign product[51] = s[50];
    assign product[52] = s[51];
    assign product[53] = s[52];
    assign product[54] = s[53];
    assign product[55] = s[54];
    assign product[56] = s[55];
    assign product[57] = s[56];
    assign product[58] = s[57];
    assign product[59] = s[58];
    assign product[60] = s[59];
    assign product[61] = s[60];
    assign product[62] = s[61];
    assign product[63] = c;
endmodule

module CLA_2(output [1:0] sum, output cout, input [1:0] in1, input [1:0] in2);

    wire[1:0] G;
    wire[1:0] C;
    wire[1:0] P;

    assign G[0] = in1[1] & in2[1];
    assign P[0] = in1[1] ^ in2[1];
    assign G[1] = in1[0] & in2[0];
    assign P[1] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign cout = G[1] | (P[1] & C[1]);
    assign sum = P ^ C;
endmodule


module CLA_2_c(output [1:0] sum,
            output cout,
            input [1:0] in1, in2,
            input cin);

    wire [1:0] G; /* Generate */
    wire [1:0] P; /* Propagate */
    wire [1:0] C; /* Carry */

    assign G[0] = in1[1] & in2[1]; /*Generate    Gi = Ai * Bi */
    assign G[1] = in1[0] & in2[0];

    assign P[0] = in1[1] ^ in2[1];
    assign P[1] = in1[0] ^ in2[0];

    assign C[0] = cin;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign cout = G[1] | (P[1] & C[1]);
    assign sum = P ^ C;
endmodule


module CLA_3(output [2:0] sum, output cout, input [2:0] in1, input [2:0] in2);

    wire[2:0] G;
    wire[2:0] C;
    wire[2:0] P;

    assign G[0] = in1[2] & in2[2];
    assign P[0] = in1[2] ^ in2[2];
    assign G[1] = in1[1] & in2[1];
    assign P[1] = in1[1] ^ in2[1];
    assign G[2] = in1[0] & in2[0];
    assign P[2] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign cout = G[2] | (P[2] & C[2]);
    assign sum = P ^ C;
endmodule

module CLA_3_c(output [2:0] sum, output cout, input [2:0] in1, input [2:0] in2, input cin);

    wire[2:0] G;
    wire[2:0] C;
    wire[2:0] P;

    assign G[0] = in1[2] & in2[2];
    assign P[0] = in1[2] ^ in2[2];
    assign G[1] = in1[1] & in2[1];
    assign P[1] = in1[1] ^ in2[1];
    assign G[2] = in1[0] & in2[0];
    assign P[2] = in1[0] ^ in2[0];


    assign C[0] = cin;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign cout = G[2] | (P[2] & C[2]);
    assign sum = P ^ C;
endmodule

module CLA_4(output [3:0] sum,
            output cout,
            input [3:0] in1, in2);

    wire [3:0] G; /* Generate */
    wire [3:0] P; /* Propagate */
    wire [3:0] C; /* Carry */

    assign G[0] = in1[3] & in2[3]; /*Generate    Gi = Ai * Bi */
    assign G[1] = in1[2] & in2[2];
    assign G[2] = in1[1] & in2[1];
    assign G[3] = in1[0] & in2[0];
    assign P[0] = in1[3] ^ in2[3]; /*Propagate   Pi = Ai + Bi */
    assign P[1] = in1[2] ^ in2[2];
    assign P[2] = in1[1] ^ in2[1];
    assign P[3] = in1[0] ^ in2[0];

    assign C[0] = 0;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign cout = G[3] | (P[3] & C[3]);
    assign sum = P ^ C;
endmodule

module CLA_4_c(output [3:0] sum,
            output cout,
            input [3:0] in1, in2,
            input cin);

    wire [3:0] G; /* Generate */
    wire [3:0] P; /* Propagate */
    wire [3:0] C; /* Carry */

    assign G[0] = in1[3] & in2[3]; /*Generate    Gi = Ai * Bi */
    assign G[1] = in1[2] & in2[2];
    assign G[2] = in1[1] & in2[1];
    assign G[3] = in1[0] & in2[0];
    assign P[0] = in1[3] ^ in2[3]; /*Propagate   Pi = Ai + Bi */
    assign P[1] = in1[2] ^ in2[2];
    assign P[2] = in1[1] ^ in2[1];
    assign P[3] = in1[0] ^ in2[0];

    assign C[0] = cin;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign cout = G[3] | (P[3] & C[3]);
    assign sum = P ^ C;
endmodule

module Half_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2);
    xor(sum, in1, in2);
    and(cout, in1, in2);
endmodule

module Full_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2,
                  input wire cin);
    wire temp1;
    wire temp2;
    wire temp3;
    xor(sum, in1, in2, cin);
    and(temp1,in1,in2);
    and(temp2,in1,cin);
    and(temp3,in2,cin);
    or(cout,temp1,temp2,temp3);
endmodule


module CLA_62(output [61:0] sum, output cout, input [61:0] in1, input [61:0] in2);

    wire[61:0] G;
    wire[61:0] C;
    wire[61:0] P;

    assign G[0] = in1[61] & in2[61];
    assign P[0] = in1[61] ^ in2[61];
    assign G[1] = in1[60] & in2[60];
    assign P[1] = in1[60] ^ in2[60];
    assign G[2] = in1[59] & in2[59];
    assign P[2] = in1[59] ^ in2[59];
    assign G[3] = in1[58] & in2[58];
    assign P[3] = in1[58] ^ in2[58];
    assign G[4] = in1[57] & in2[57];
    assign P[4] = in1[57] ^ in2[57];
    assign G[5] = in1[56] & in2[56];
    assign P[5] = in1[56] ^ in2[56];
    assign G[6] = in1[55] & in2[55];
    assign P[6] = in1[55] ^ in2[55];
    assign G[7] = in1[54] & in2[54];
    assign P[7] = in1[54] ^ in2[54];
    assign G[8] = in1[53] & in2[53];
    assign P[8] = in1[53] ^ in2[53];
    assign G[9] = in1[52] & in2[52];
    assign P[9] = in1[52] ^ in2[52];
    assign G[10] = in1[51] & in2[51];
    assign P[10] = in1[51] ^ in2[51];
    assign G[11] = in1[50] & in2[50];
    assign P[11] = in1[50] ^ in2[50];
    assign G[12] = in1[49] & in2[49];
    assign P[12] = in1[49] ^ in2[49];
    assign G[13] = in1[48] & in2[48];
    assign P[13] = in1[48] ^ in2[48];
    assign G[14] = in1[47] & in2[47];
    assign P[14] = in1[47] ^ in2[47];
    assign G[15] = in1[46] & in2[46];
    assign P[15] = in1[46] ^ in2[46];
    assign G[16] = in1[45] & in2[45];
    assign P[16] = in1[45] ^ in2[45];
    assign G[17] = in1[44] & in2[44];
    assign P[17] = in1[44] ^ in2[44];
    assign G[18] = in1[43] & in2[43];
    assign P[18] = in1[43] ^ in2[43];
    assign G[19] = in1[42] & in2[42];
    assign P[19] = in1[42] ^ in2[42];
    assign G[20] = in1[41] & in2[41];
    assign P[20] = in1[41] ^ in2[41];
    assign G[21] = in1[40] & in2[40];
    assign P[21] = in1[40] ^ in2[40];
    assign G[22] = in1[39] & in2[39];
    assign P[22] = in1[39] ^ in2[39];
    assign G[23] = in1[38] & in2[38];
    assign P[23] = in1[38] ^ in2[38];
    assign G[24] = in1[37] & in2[37];
    assign P[24] = in1[37] ^ in2[37];
    assign G[25] = in1[36] & in2[36];
    assign P[25] = in1[36] ^ in2[36];
    assign G[26] = in1[35] & in2[35];
    assign P[26] = in1[35] ^ in2[35];
    assign G[27] = in1[34] & in2[34];
    assign P[27] = in1[34] ^ in2[34];
    assign G[28] = in1[33] & in2[33];
    assign P[28] = in1[33] ^ in2[33];
    assign G[29] = in1[32] & in2[32];
    assign P[29] = in1[32] ^ in2[32];
    assign G[30] = in1[31] & in2[31];
    assign P[30] = in1[31] ^ in2[31];
    assign G[31] = in1[30] & in2[30];
    assign P[31] = in1[30] ^ in2[30];
    assign G[32] = in1[29] & in2[29];
    assign P[32] = in1[29] ^ in2[29];
    assign G[33] = in1[28] & in2[28];
    assign P[33] = in1[28] ^ in2[28];
    assign G[34] = in1[27] & in2[27];
    assign P[34] = in1[27] ^ in2[27];
    assign G[35] = in1[26] & in2[26];
    assign P[35] = in1[26] ^ in2[26];
    assign G[36] = in1[25] & in2[25];
    assign P[36] = in1[25] ^ in2[25];
    assign G[37] = in1[24] & in2[24];
    assign P[37] = in1[24] ^ in2[24];
    assign G[38] = in1[23] & in2[23];
    assign P[38] = in1[23] ^ in2[23];
    assign G[39] = in1[22] & in2[22];
    assign P[39] = in1[22] ^ in2[22];
    assign G[40] = in1[21] & in2[21];
    assign P[40] = in1[21] ^ in2[21];
    assign G[41] = in1[20] & in2[20];
    assign P[41] = in1[20] ^ in2[20];
    assign G[42] = in1[19] & in2[19];
    assign P[42] = in1[19] ^ in2[19];
    assign G[43] = in1[18] & in2[18];
    assign P[43] = in1[18] ^ in2[18];
    assign G[44] = in1[17] & in2[17];
    assign P[44] = in1[17] ^ in2[17];
    assign G[45] = in1[16] & in2[16];
    assign P[45] = in1[16] ^ in2[16];
    assign G[46] = in1[15] & in2[15];
    assign P[46] = in1[15] ^ in2[15];
    assign G[47] = in1[14] & in2[14];
    assign P[47] = in1[14] ^ in2[14];
    assign G[48] = in1[13] & in2[13];
    assign P[48] = in1[13] ^ in2[13];
    assign G[49] = in1[12] & in2[12];
    assign P[49] = in1[12] ^ in2[12];
    assign G[50] = in1[11] & in2[11];
    assign P[50] = in1[11] ^ in2[11];
    assign G[51] = in1[10] & in2[10];
    assign P[51] = in1[10] ^ in2[10];
    assign G[52] = in1[9] & in2[9];
    assign P[52] = in1[9] ^ in2[9];
    assign G[53] = in1[8] & in2[8];
    assign P[53] = in1[8] ^ in2[8];
    assign G[54] = in1[7] & in2[7];
    assign P[54] = in1[7] ^ in2[7];
    assign G[55] = in1[6] & in2[6];
    assign P[55] = in1[6] ^ in2[6];
    assign G[56] = in1[5] & in2[5];
    assign P[56] = in1[5] ^ in2[5];
    assign G[57] = in1[4] & in2[4];
    assign P[57] = in1[4] ^ in2[4];
    assign G[58] = in1[3] & in2[3];
    assign P[58] = in1[3] ^ in2[3];
    assign G[59] = in1[2] & in2[2];
    assign P[59] = in1[2] ^ in2[2];
    assign G[60] = in1[1] & in2[1];
    assign P[60] = in1[1] ^ in2[1];
    assign G[61] = in1[0] & in2[0];
    assign P[61] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign cout = G[61] | (P[61] & C[61]);
    assign sum = P ^ C;
endmodule

