module dadda_unsigned_multiplier_CLA_64(product, A, B);
    input [63:0] A, B;
    output [127:0] product;

    wire [63:0] pp0;
    wire [63:0] pp1;
    wire [63:0] pp2;
    wire [63:0] pp3;
    wire [63:0] pp4;
    wire [63:0] pp5;
    wire [63:0] pp6;
    wire [63:0] pp7;
    wire [63:0] pp8;
    wire [63:0] pp9;
    wire [63:0] pp10;
    wire [63:0] pp11;
    wire [63:0] pp12;
    wire [63:0] pp13;
    wire [63:0] pp14;
    wire [63:0] pp15;
    wire [63:0] pp16;
    wire [63:0] pp17;
    wire [63:0] pp18;
    wire [63:0] pp19;
    wire [63:0] pp20;
    wire [63:0] pp21;
    wire [63:0] pp22;
    wire [63:0] pp23;
    wire [63:0] pp24;
    wire [63:0] pp25;
    wire [63:0] pp26;
    wire [63:0] pp27;
    wire [63:0] pp28;
    wire [63:0] pp29;
    wire [63:0] pp30;
    wire [63:0] pp31;
    wire [63:0] pp32;
    wire [63:0] pp33;
    wire [63:0] pp34;
    wire [63:0] pp35;
    wire [63:0] pp36;
    wire [63:0] pp37;
    wire [63:0] pp38;
    wire [63:0] pp39;
    wire [63:0] pp40;
    wire [63:0] pp41;
    wire [63:0] pp42;
    wire [63:0] pp43;
    wire [63:0] pp44;
    wire [63:0] pp45;
    wire [63:0] pp46;
    wire [63:0] pp47;
    wire [63:0] pp48;
    wire [63:0] pp49;
    wire [63:0] pp50;
    wire [63:0] pp51;
    wire [63:0] pp52;
    wire [63:0] pp53;
    wire [63:0] pp54;
    wire [63:0] pp55;
    wire [63:0] pp56;
    wire [63:0] pp57;
    wire [63:0] pp58;
    wire [63:0] pp59;
    wire [63:0] pp60;
    wire [63:0] pp61;
    wire [63:0] pp62;
    wire [63:0] pp63;
	
	wire [127:0] product;

    assign pp0 = A[0] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp1 = A[1] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp2 = A[2] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp3 = A[3] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp4 = A[4] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp5 = A[5] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp6 = A[6] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp7 = A[7] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp8 = A[8] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp9 = A[9] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp10 = A[10] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp11 = A[11] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp12 = A[12] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp13 = A[13] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp14 = A[14] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp15 = A[15] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp16 = A[16] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp17 = A[17] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp18 = A[18] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp19 = A[19] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp20 = A[20] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp21 = A[21] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp22 = A[22] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp23 = A[23] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp24 = A[24] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp25 = A[25] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp26 = A[26] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp27 = A[27] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp28 = A[28] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp29 = A[29] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp30 = A[30] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp31 = A[31] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp32 = A[32] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp33 = A[33] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp34 = A[34] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp35 = A[35] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp36 = A[36] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp37 = A[37] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp38 = A[38] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp39 = A[39] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp40 = A[40] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp41 = A[41] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp42 = A[42] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp43 = A[43] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp44 = A[44] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp45 = A[45] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp46 = A[46] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp47 = A[47] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp48 = A[48] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp49 = A[49] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp50 = A[50] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp51 = A[51] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp52 = A[52] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp53 = A[53] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp54 = A[54] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp55 = A[55] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp56 = A[56] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp57 = A[57] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp58 = A[58] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp59 = A[59] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp60 = A[60] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp61 = A[61] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp62 = A[62] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp63 = A[63] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
	
	wire [4032:0] S;
	wire [4032:0] Cout;
	Half_Adder HA1 (pp0[63], pp1[62], S[1], Cout[1]);
	Half_Adder HA2 (pp1[63], pp2[62], S[2], Cout[2]);
	Half_Adder HA3 (pp0[42], pp1[41], S[3], Cout[3]);
	Full_Adder FA1 (pp0[43], pp1[42], pp2[41], S[4], Cout[4]);
	Half_Adder HA4 (pp3[40], pp4[39], S[5], Cout[5]);
	Full_Adder FA2 (pp0[44], pp1[43], pp2[42], S[6], Cout[6]);
	Full_Adder FA3 (pp3[41], pp4[40], pp5[39], S[7], Cout[7]);
	Half_Adder HA5 (pp6[38], pp7[37], S[8], Cout[8]);
	Full_Adder FA4 (pp0[45], pp1[44], pp2[43], S[9], Cout[9]);
	Full_Adder FA5 (pp3[42], pp4[41], pp5[40], S[10], Cout[10]);
	Full_Adder FA6 (pp6[39], pp7[38], pp8[37], S[11], Cout[11]);
	Half_Adder HA6 (pp9[36], pp10[35], S[12], Cout[12]);
	Full_Adder FA7 (pp0[46], pp1[45], pp2[44], S[13], Cout[13]);
	Full_Adder FA8 (pp3[43], pp4[42], pp5[41], S[14], Cout[14]);
	Full_Adder FA9 (pp6[40], pp7[39], pp8[38], S[15], Cout[15]);
	Full_Adder FA10 (pp9[37], pp10[36], pp11[35], S[16], Cout[16]);
	Half_Adder HA7 (pp12[34], pp13[33], S[17], Cout[17]);
	Full_Adder FA11 (pp0[47], pp1[46], pp2[45], S[18], Cout[18]);
	Full_Adder FA12 (pp3[44], pp4[43], pp5[42], S[19], Cout[19]);
	Full_Adder FA13 (pp6[41], pp7[40], pp8[39], S[20], Cout[20]);
	Full_Adder FA14 (pp9[38], pp10[37], pp11[36], S[21], Cout[21]);
	Full_Adder FA15 (pp12[35], pp13[34], pp14[33], S[22], Cout[22]);
	Half_Adder HA8 (pp15[32], pp16[31], S[23], Cout[23]);
	Full_Adder FA16 (pp0[48], pp1[47], pp2[46], S[24], Cout[24]);
	Full_Adder FA17 (pp3[45], pp4[44], pp5[43], S[25], Cout[25]);
	Full_Adder FA18 (pp6[42], pp7[41], pp8[40], S[26], Cout[26]);
	Full_Adder FA19 (pp9[39], pp10[38], pp11[37], S[27], Cout[27]);
	Full_Adder FA20 (pp12[36], pp13[35], pp14[34], S[28], Cout[28]);
	Full_Adder FA21 (pp15[33], pp16[32], pp17[31], S[29], Cout[29]);
	Half_Adder HA9 (pp18[30], pp19[29], S[30], Cout[30]);
	Full_Adder FA22 (pp0[49], pp1[48], pp2[47], S[31], Cout[31]);
	Full_Adder FA23 (pp3[46], pp4[45], pp5[44], S[32], Cout[32]);
	Full_Adder FA24 (pp6[43], pp7[42], pp8[41], S[33], Cout[33]);
	Full_Adder FA25 (pp9[40], pp10[39], pp11[38], S[34], Cout[34]);
	Full_Adder FA26 (pp12[37], pp13[36], pp14[35], S[35], Cout[35]);
	Full_Adder FA27 (pp15[34], pp16[33], pp17[32], S[36], Cout[36]);
	Full_Adder FA28 (pp18[31], pp19[30], pp20[29], S[37], Cout[37]);
	Half_Adder HA10 (pp21[28], pp22[27], S[38], Cout[38]);
	Full_Adder FA29 (pp0[50], pp1[49], pp2[48], S[39], Cout[39]);
	Full_Adder FA30 (pp3[47], pp4[46], pp5[45], S[40], Cout[40]);
	Full_Adder FA31 (pp6[44], pp7[43], pp8[42], S[41], Cout[41]);
	Full_Adder FA32 (pp9[41], pp10[40], pp11[39], S[42], Cout[42]);
	Full_Adder FA33 (pp12[38], pp13[37], pp14[36], S[43], Cout[43]);
	Full_Adder FA34 (pp15[35], pp16[34], pp17[33], S[44], Cout[44]);
	Full_Adder FA35 (pp18[32], pp19[31], pp20[30], S[45], Cout[45]);
	Full_Adder FA36 (pp21[29], pp22[28], pp23[27], S[46], Cout[46]);
	Half_Adder HA11 (pp24[26], pp25[25], S[47], Cout[47]);
	Full_Adder FA37 (pp0[51], pp1[50], pp2[49], S[48], Cout[48]);
	Full_Adder FA38 (pp3[48], pp4[47], pp5[46], S[49], Cout[49]);
	Full_Adder FA39 (pp6[45], pp7[44], pp8[43], S[50], Cout[50]);
	Full_Adder FA40 (pp9[42], pp10[41], pp11[40], S[51], Cout[51]);
	Full_Adder FA41 (pp12[39], pp13[38], pp14[37], S[52], Cout[52]);
	Full_Adder FA42 (pp15[36], pp16[35], pp17[34], S[53], Cout[53]);
	Full_Adder FA43 (pp18[33], pp19[32], pp20[31], S[54], Cout[54]);
	Full_Adder FA44 (pp21[30], pp22[29], pp23[28], S[55], Cout[55]);
	Full_Adder FA45 (pp24[27], pp25[26], pp26[25], S[56], Cout[56]);
	Half_Adder HA12 (pp27[24], pp28[23], S[57], Cout[57]);
	Full_Adder FA46 (pp0[52], pp1[51], pp2[50], S[58], Cout[58]);
	Full_Adder FA47 (pp3[49], pp4[48], pp5[47], S[59], Cout[59]);
	Full_Adder FA48 (pp6[46], pp7[45], pp8[44], S[60], Cout[60]);
	Full_Adder FA49 (pp9[43], pp10[42], pp11[41], S[61], Cout[61]);
	Full_Adder FA50 (pp12[40], pp13[39], pp14[38], S[62], Cout[62]);
	Full_Adder FA51 (pp15[37], pp16[36], pp17[35], S[63], Cout[63]);
	Full_Adder FA52 (pp18[34], pp19[33], pp20[32], S[64], Cout[64]);
	Full_Adder FA53 (pp21[31], pp22[30], pp23[29], S[65], Cout[65]);
	Full_Adder FA54 (pp24[28], pp25[27], pp26[26], S[66], Cout[66]);
	Full_Adder FA55 (pp27[25], pp28[24], pp29[23], S[67], Cout[67]);
	Half_Adder HA13 (pp30[22], pp31[21], S[68], Cout[68]);
	Full_Adder FA56 (pp0[53], pp1[52], pp2[51], S[69], Cout[69]);
	Full_Adder FA57 (pp3[50], pp4[49], pp5[48], S[70], Cout[70]);
	Full_Adder FA58 (pp6[47], pp7[46], pp8[45], S[71], Cout[71]);
	Full_Adder FA59 (pp9[44], pp10[43], pp11[42], S[72], Cout[72]);
	Full_Adder FA60 (pp12[41], pp13[40], pp14[39], S[73], Cout[73]);
	Full_Adder FA61 (pp15[38], pp16[37], pp17[36], S[74], Cout[74]);
	Full_Adder FA62 (pp18[35], pp19[34], pp20[33], S[75], Cout[75]);
	Full_Adder FA63 (pp21[32], pp22[31], pp23[30], S[76], Cout[76]);
	Full_Adder FA64 (pp24[29], pp25[28], pp26[27], S[77], Cout[77]);
	Full_Adder FA65 (pp27[26], pp28[25], pp29[24], S[78], Cout[78]);
	Full_Adder FA66 (pp30[23], pp31[22], pp32[21], S[79], Cout[79]);
	Half_Adder HA14 (pp33[20], pp34[19], S[80], Cout[80]);
	Full_Adder FA67 (pp0[54], pp1[53], pp2[52], S[81], Cout[81]);
	Full_Adder FA68 (pp3[51], pp4[50], pp5[49], S[82], Cout[82]);
	Full_Adder FA69 (pp6[48], pp7[47], pp8[46], S[83], Cout[83]);
	Full_Adder FA70 (pp9[45], pp10[44], pp11[43], S[84], Cout[84]);
	Full_Adder FA71 (pp12[42], pp13[41], pp14[40], S[85], Cout[85]);
	Full_Adder FA72 (pp15[39], pp16[38], pp17[37], S[86], Cout[86]);
	Full_Adder FA73 (pp18[36], pp19[35], pp20[34], S[87], Cout[87]);
	Full_Adder FA74 (pp21[33], pp22[32], pp23[31], S[88], Cout[88]);
	Full_Adder FA75 (pp24[30], pp25[29], pp26[28], S[89], Cout[89]);
	Full_Adder FA76 (pp27[27], pp28[26], pp29[25], S[90], Cout[90]);
	Full_Adder FA77 (pp30[24], pp31[23], pp32[22], S[91], Cout[91]);
	Full_Adder FA78 (pp33[21], pp34[20], pp35[19], S[92], Cout[92]);
	Half_Adder HA15 (pp36[18], pp37[17], S[93], Cout[93]);
	Full_Adder FA79 (pp0[55], pp1[54], pp2[53], S[94], Cout[94]);
	Full_Adder FA80 (pp3[52], pp4[51], pp5[50], S[95], Cout[95]);
	Full_Adder FA81 (pp6[49], pp7[48], pp8[47], S[96], Cout[96]);
	Full_Adder FA82 (pp9[46], pp10[45], pp11[44], S[97], Cout[97]);
	Full_Adder FA83 (pp12[43], pp13[42], pp14[41], S[98], Cout[98]);
	Full_Adder FA84 (pp15[40], pp16[39], pp17[38], S[99], Cout[99]);
	Full_Adder FA85 (pp18[37], pp19[36], pp20[35], S[100], Cout[100]);
	Full_Adder FA86 (pp21[34], pp22[33], pp23[32], S[101], Cout[101]);
	Full_Adder FA87 (pp24[31], pp25[30], pp26[29], S[102], Cout[102]);
	Full_Adder FA88 (pp27[28], pp28[27], pp29[26], S[103], Cout[103]);
	Full_Adder FA89 (pp30[25], pp31[24], pp32[23], S[104], Cout[104]);
	Full_Adder FA90 (pp33[22], pp34[21], pp35[20], S[105], Cout[105]);
	Full_Adder FA91 (pp36[19], pp37[18], pp38[17], S[106], Cout[106]);
	Half_Adder HA16 (pp39[16], pp40[15], S[107], Cout[107]);
	Full_Adder FA92 (pp0[56], pp1[55], pp2[54], S[108], Cout[108]);
	Full_Adder FA93 (pp3[53], pp4[52], pp5[51], S[109], Cout[109]);
	Full_Adder FA94 (pp6[50], pp7[49], pp8[48], S[110], Cout[110]);
	Full_Adder FA95 (pp9[47], pp10[46], pp11[45], S[111], Cout[111]);
	Full_Adder FA96 (pp12[44], pp13[43], pp14[42], S[112], Cout[112]);
	Full_Adder FA97 (pp15[41], pp16[40], pp17[39], S[113], Cout[113]);
	Full_Adder FA98 (pp18[38], pp19[37], pp20[36], S[114], Cout[114]);
	Full_Adder FA99 (pp21[35], pp22[34], pp23[33], S[115], Cout[115]);
	Full_Adder FA100 (pp24[32], pp25[31], pp26[30], S[116], Cout[116]);
	Full_Adder FA101 (pp27[29], pp28[28], pp29[27], S[117], Cout[117]);
	Full_Adder FA102 (pp30[26], pp31[25], pp32[24], S[118], Cout[118]);
	Full_Adder FA103 (pp33[23], pp34[22], pp35[21], S[119], Cout[119]);
	Full_Adder FA104 (pp36[20], pp37[19], pp38[18], S[120], Cout[120]);
	Full_Adder FA105 (pp39[17], pp40[16], pp41[15], S[121], Cout[121]);
	Half_Adder HA17 (pp42[14], pp43[13], S[122], Cout[122]);
	Full_Adder FA106 (pp0[57], pp1[56], pp2[55], S[123], Cout[123]);
	Full_Adder FA107 (pp3[54], pp4[53], pp5[52], S[124], Cout[124]);
	Full_Adder FA108 (pp6[51], pp7[50], pp8[49], S[125], Cout[125]);
	Full_Adder FA109 (pp9[48], pp10[47], pp11[46], S[126], Cout[126]);
	Full_Adder FA110 (pp12[45], pp13[44], pp14[43], S[127], Cout[127]);
	Full_Adder FA111 (pp15[42], pp16[41], pp17[40], S[128], Cout[128]);
	Full_Adder FA112 (pp18[39], pp19[38], pp20[37], S[129], Cout[129]);
	Full_Adder FA113 (pp21[36], pp22[35], pp23[34], S[130], Cout[130]);
	Full_Adder FA114 (pp24[33], pp25[32], pp26[31], S[131], Cout[131]);
	Full_Adder FA115 (pp27[30], pp28[29], pp29[28], S[132], Cout[132]);
	Full_Adder FA116 (pp30[27], pp31[26], pp32[25], S[133], Cout[133]);
	Full_Adder FA117 (pp33[24], pp34[23], pp35[22], S[134], Cout[134]);
	Full_Adder FA118 (pp36[21], pp37[20], pp38[19], S[135], Cout[135]);
	Full_Adder FA119 (pp39[18], pp40[17], pp41[16], S[136], Cout[136]);
	Full_Adder FA120 (pp42[15], pp43[14], pp44[13], S[137], Cout[137]);
	Half_Adder HA18 (pp45[12], pp46[11], S[138], Cout[138]);
	Full_Adder FA121 (pp0[58], pp1[57], pp2[56], S[139], Cout[139]);
	Full_Adder FA122 (pp3[55], pp4[54], pp5[53], S[140], Cout[140]);
	Full_Adder FA123 (pp6[52], pp7[51], pp8[50], S[141], Cout[141]);
	Full_Adder FA124 (pp9[49], pp10[48], pp11[47], S[142], Cout[142]);
	Full_Adder FA125 (pp12[46], pp13[45], pp14[44], S[143], Cout[143]);
	Full_Adder FA126 (pp15[43], pp16[42], pp17[41], S[144], Cout[144]);
	Full_Adder FA127 (pp18[40], pp19[39], pp20[38], S[145], Cout[145]);
	Full_Adder FA128 (pp21[37], pp22[36], pp23[35], S[146], Cout[146]);
	Full_Adder FA129 (pp24[34], pp25[33], pp26[32], S[147], Cout[147]);
	Full_Adder FA130 (pp27[31], pp28[30], pp29[29], S[148], Cout[148]);
	Full_Adder FA131 (pp30[28], pp31[27], pp32[26], S[149], Cout[149]);
	Full_Adder FA132 (pp33[25], pp34[24], pp35[23], S[150], Cout[150]);
	Full_Adder FA133 (pp36[22], pp37[21], pp38[20], S[151], Cout[151]);
	Full_Adder FA134 (pp39[19], pp40[18], pp41[17], S[152], Cout[152]);
	Full_Adder FA135 (pp42[16], pp43[15], pp44[14], S[153], Cout[153]);
	Full_Adder FA136 (pp45[13], pp46[12], pp47[11], S[154], Cout[154]);
	Half_Adder HA19 (pp48[10], pp49[9], S[155], Cout[155]);
	Full_Adder FA137 (pp0[59], pp1[58], pp2[57], S[156], Cout[156]);
	Full_Adder FA138 (pp3[56], pp4[55], pp5[54], S[157], Cout[157]);
	Full_Adder FA139 (pp6[53], pp7[52], pp8[51], S[158], Cout[158]);
	Full_Adder FA140 (pp9[50], pp10[49], pp11[48], S[159], Cout[159]);
	Full_Adder FA141 (pp12[47], pp13[46], pp14[45], S[160], Cout[160]);
	Full_Adder FA142 (pp15[44], pp16[43], pp17[42], S[161], Cout[161]);
	Full_Adder FA143 (pp18[41], pp19[40], pp20[39], S[162], Cout[162]);
	Full_Adder FA144 (pp21[38], pp22[37], pp23[36], S[163], Cout[163]);
	Full_Adder FA145 (pp24[35], pp25[34], pp26[33], S[164], Cout[164]);
	Full_Adder FA146 (pp27[32], pp28[31], pp29[30], S[165], Cout[165]);
	Full_Adder FA147 (pp30[29], pp31[28], pp32[27], S[166], Cout[166]);
	Full_Adder FA148 (pp33[26], pp34[25], pp35[24], S[167], Cout[167]);
	Full_Adder FA149 (pp36[23], pp37[22], pp38[21], S[168], Cout[168]);
	Full_Adder FA150 (pp39[20], pp40[19], pp41[18], S[169], Cout[169]);
	Full_Adder FA151 (pp42[17], pp43[16], pp44[15], S[170], Cout[170]);
	Full_Adder FA152 (pp45[14], pp46[13], pp47[12], S[171], Cout[171]);
	Full_Adder FA153 (pp48[11], pp49[10], pp50[9], S[172], Cout[172]);
	Half_Adder HA20 (pp51[8], pp52[7], S[173], Cout[173]);
	Full_Adder FA154 (pp0[60], pp1[59], pp2[58], S[174], Cout[174]);
	Full_Adder FA155 (pp3[57], pp4[56], pp5[55], S[175], Cout[175]);
	Full_Adder FA156 (pp6[54], pp7[53], pp8[52], S[176], Cout[176]);
	Full_Adder FA157 (pp9[51], pp10[50], pp11[49], S[177], Cout[177]);
	Full_Adder FA158 (pp12[48], pp13[47], pp14[46], S[178], Cout[178]);
	Full_Adder FA159 (pp15[45], pp16[44], pp17[43], S[179], Cout[179]);
	Full_Adder FA160 (pp18[42], pp19[41], pp20[40], S[180], Cout[180]);
	Full_Adder FA161 (pp21[39], pp22[38], pp23[37], S[181], Cout[181]);
	Full_Adder FA162 (pp24[36], pp25[35], pp26[34], S[182], Cout[182]);
	Full_Adder FA163 (pp27[33], pp28[32], pp29[31], S[183], Cout[183]);
	Full_Adder FA164 (pp30[30], pp31[29], pp32[28], S[184], Cout[184]);
	Full_Adder FA165 (pp33[27], pp34[26], pp35[25], S[185], Cout[185]);
	Full_Adder FA166 (pp36[24], pp37[23], pp38[22], S[186], Cout[186]);
	Full_Adder FA167 (pp39[21], pp40[20], pp41[19], S[187], Cout[187]);
	Full_Adder FA168 (pp42[18], pp43[17], pp44[16], S[188], Cout[188]);
	Full_Adder FA169 (pp45[15], pp46[14], pp47[13], S[189], Cout[189]);
	Full_Adder FA170 (pp48[12], pp49[11], pp50[10], S[190], Cout[190]);
	Full_Adder FA171 (pp51[9], pp52[8], pp53[7], S[191], Cout[191]);
	Half_Adder HA21 (pp54[6], pp55[5], S[192], Cout[192]);
	Full_Adder FA172 (pp0[61], pp1[60], pp2[59], S[193], Cout[193]);
	Full_Adder FA173 (pp3[58], pp4[57], pp5[56], S[194], Cout[194]);
	Full_Adder FA174 (pp6[55], pp7[54], pp8[53], S[195], Cout[195]);
	Full_Adder FA175 (pp9[52], pp10[51], pp11[50], S[196], Cout[196]);
	Full_Adder FA176 (pp12[49], pp13[48], pp14[47], S[197], Cout[197]);
	Full_Adder FA177 (pp15[46], pp16[45], pp17[44], S[198], Cout[198]);
	Full_Adder FA178 (pp18[43], pp19[42], pp20[41], S[199], Cout[199]);
	Full_Adder FA179 (pp21[40], pp22[39], pp23[38], S[200], Cout[200]);
	Full_Adder FA180 (pp24[37], pp25[36], pp26[35], S[201], Cout[201]);
	Full_Adder FA181 (pp27[34], pp28[33], pp29[32], S[202], Cout[202]);
	Full_Adder FA182 (pp30[31], pp31[30], pp32[29], S[203], Cout[203]);
	Full_Adder FA183 (pp33[28], pp34[27], pp35[26], S[204], Cout[204]);
	Full_Adder FA184 (pp36[25], pp37[24], pp38[23], S[205], Cout[205]);
	Full_Adder FA185 (pp39[22], pp40[21], pp41[20], S[206], Cout[206]);
	Full_Adder FA186 (pp42[19], pp43[18], pp44[17], S[207], Cout[207]);
	Full_Adder FA187 (pp45[16], pp46[15], pp47[14], S[208], Cout[208]);
	Full_Adder FA188 (pp48[13], pp49[12], pp50[11], S[209], Cout[209]);
	Full_Adder FA189 (pp51[10], pp52[9], pp53[8], S[210], Cout[210]);
	Full_Adder FA190 (pp54[7], pp55[6], pp56[5], S[211], Cout[211]);
	Half_Adder HA22 (pp57[4], pp58[3], S[212], Cout[212]);
	Full_Adder FA191 (pp0[62], pp1[61], pp2[60], S[213], Cout[213]);
	Full_Adder FA192 (pp3[59], pp4[58], pp5[57], S[214], Cout[214]);
	Full_Adder FA193 (pp6[56], pp7[55], pp8[54], S[215], Cout[215]);
	Full_Adder FA194 (pp9[53], pp10[52], pp11[51], S[216], Cout[216]);
	Full_Adder FA195 (pp12[50], pp13[49], pp14[48], S[217], Cout[217]);
	Full_Adder FA196 (pp15[47], pp16[46], pp17[45], S[218], Cout[218]);
	Full_Adder FA197 (pp18[44], pp19[43], pp20[42], S[219], Cout[219]);
	Full_Adder FA198 (pp21[41], pp22[40], pp23[39], S[220], Cout[220]);
	Full_Adder FA199 (pp24[38], pp25[37], pp26[36], S[221], Cout[221]);
	Full_Adder FA200 (pp27[35], pp28[34], pp29[33], S[222], Cout[222]);
	Full_Adder FA201 (pp30[32], pp31[31], pp32[30], S[223], Cout[223]);
	Full_Adder FA202 (pp33[29], pp34[28], pp35[27], S[224], Cout[224]);
	Full_Adder FA203 (pp36[26], pp37[25], pp38[24], S[225], Cout[225]);
	Full_Adder FA204 (pp39[23], pp40[22], pp41[21], S[226], Cout[226]);
	Full_Adder FA205 (pp42[20], pp43[19], pp44[18], S[227], Cout[227]);
	Full_Adder FA206 (pp45[17], pp46[16], pp47[15], S[228], Cout[228]);
	Full_Adder FA207 (pp48[14], pp49[13], pp50[12], S[229], Cout[229]);
	Full_Adder FA208 (pp51[11], pp52[10], pp53[9], S[230], Cout[230]);
	Full_Adder FA209 (pp54[8], pp55[7], pp56[6], S[231], Cout[231]);
	Full_Adder FA210 (pp57[5], pp58[4], pp59[3], S[232], Cout[232]);
	Half_Adder HA23 (pp60[2], pp61[1], S[233], Cout[233]);
	Full_Adder FA211 (pp2[61], pp3[60], pp4[59], S[234], Cout[234]);
	Full_Adder FA212 (pp5[58], pp6[57], pp7[56], S[235], Cout[235]);
	Full_Adder FA213 (pp8[55], pp9[54], pp10[53], S[236], Cout[236]);
	Full_Adder FA214 (pp11[52], pp12[51], pp13[50], S[237], Cout[237]);
	Full_Adder FA215 (pp14[49], pp15[48], pp16[47], S[238], Cout[238]);
	Full_Adder FA216 (pp17[46], pp18[45], pp19[44], S[239], Cout[239]);
	Full_Adder FA217 (pp20[43], pp21[42], pp22[41], S[240], Cout[240]);
	Full_Adder FA218 (pp23[40], pp24[39], pp25[38], S[241], Cout[241]);
	Full_Adder FA219 (pp26[37], pp27[36], pp28[35], S[242], Cout[242]);
	Full_Adder FA220 (pp29[34], pp30[33], pp31[32], S[243], Cout[243]);
	Full_Adder FA221 (pp32[31], pp33[30], pp34[29], S[244], Cout[244]);
	Full_Adder FA222 (pp35[28], pp36[27], pp37[26], S[245], Cout[245]);
	Full_Adder FA223 (pp38[25], pp39[24], pp40[23], S[246], Cout[246]);
	Full_Adder FA224 (pp41[22], pp42[21], pp43[20], S[247], Cout[247]);
	Full_Adder FA225 (pp44[19], pp45[18], pp46[17], S[248], Cout[248]);
	Full_Adder FA226 (pp47[16], pp48[15], pp49[14], S[249], Cout[249]);
	Full_Adder FA227 (pp50[13], pp51[12], pp52[11], S[250], Cout[250]);
	Full_Adder FA228 (pp53[10], pp54[9], pp55[8], S[251], Cout[251]);
	Full_Adder FA229 (pp56[7], pp57[6], pp58[5], S[252], Cout[252]);
	Full_Adder FA230 (pp59[4], pp60[3], pp61[2], S[253], Cout[253]);
	Full_Adder FA231 (pp62[1], pp63[0], S[1], S[254], Cout[254]);
	Full_Adder FA232 (pp3[61], pp4[60], pp5[59], S[255], Cout[255]);
	Full_Adder FA233 (pp6[58], pp7[57], pp8[56], S[256], Cout[256]);
	Full_Adder FA234 (pp9[55], pp10[54], pp11[53], S[257], Cout[257]);
	Full_Adder FA235 (pp12[52], pp13[51], pp14[50], S[258], Cout[258]);
	Full_Adder FA236 (pp15[49], pp16[48], pp17[47], S[259], Cout[259]);
	Full_Adder FA237 (pp18[46], pp19[45], pp20[44], S[260], Cout[260]);
	Full_Adder FA238 (pp21[43], pp22[42], pp23[41], S[261], Cout[261]);
	Full_Adder FA239 (pp24[40], pp25[39], pp26[38], S[262], Cout[262]);
	Full_Adder FA240 (pp27[37], pp28[36], pp29[35], S[263], Cout[263]);
	Full_Adder FA241 (pp30[34], pp31[33], pp32[32], S[264], Cout[264]);
	Full_Adder FA242 (pp33[31], pp34[30], pp35[29], S[265], Cout[265]);
	Full_Adder FA243 (pp36[28], pp37[27], pp38[26], S[266], Cout[266]);
	Full_Adder FA244 (pp39[25], pp40[24], pp41[23], S[267], Cout[267]);
	Full_Adder FA245 (pp42[22], pp43[21], pp44[20], S[268], Cout[268]);
	Full_Adder FA246 (pp45[19], pp46[18], pp47[17], S[269], Cout[269]);
	Full_Adder FA247 (pp48[16], pp49[15], pp50[14], S[270], Cout[270]);
	Full_Adder FA248 (pp51[13], pp52[12], pp53[11], S[271], Cout[271]);
	Full_Adder FA249 (pp54[10], pp55[9], pp56[8], S[272], Cout[272]);
	Full_Adder FA250 (pp57[7], pp58[6], pp59[5], S[273], Cout[273]);
	Full_Adder FA251 (pp60[4], pp61[3], pp62[2], S[274], Cout[274]);
	Full_Adder FA252 (pp63[1], Cout[1], S[2], S[275], Cout[275]);
	Full_Adder FA253 (pp2[63], pp3[62], pp4[61], S[276], Cout[276]);
	Full_Adder FA254 (pp5[60], pp6[59], pp7[58], S[277], Cout[277]);
	Full_Adder FA255 (pp8[57], pp9[56], pp10[55], S[278], Cout[278]);
	Full_Adder FA256 (pp11[54], pp12[53], pp13[52], S[279], Cout[279]);
	Full_Adder FA257 (pp14[51], pp15[50], pp16[49], S[280], Cout[280]);
	Full_Adder FA258 (pp17[48], pp18[47], pp19[46], S[281], Cout[281]);
	Full_Adder FA259 (pp20[45], pp21[44], pp22[43], S[282], Cout[282]);
	Full_Adder FA260 (pp23[42], pp24[41], pp25[40], S[283], Cout[283]);
	Full_Adder FA261 (pp26[39], pp27[38], pp28[37], S[284], Cout[284]);
	Full_Adder FA262 (pp29[36], pp30[35], pp31[34], S[285], Cout[285]);
	Full_Adder FA263 (pp32[33], pp33[32], pp34[31], S[286], Cout[286]);
	Full_Adder FA264 (pp35[30], pp36[29], pp37[28], S[287], Cout[287]);
	Full_Adder FA265 (pp38[27], pp39[26], pp40[25], S[288], Cout[288]);
	Full_Adder FA266 (pp41[24], pp42[23], pp43[22], S[289], Cout[289]);
	Full_Adder FA267 (pp44[21], pp45[20], pp46[19], S[290], Cout[290]);
	Full_Adder FA268 (pp47[18], pp48[17], pp49[16], S[291], Cout[291]);
	Full_Adder FA269 (pp50[15], pp51[14], pp52[13], S[292], Cout[292]);
	Full_Adder FA270 (pp53[12], pp54[11], pp55[10], S[293], Cout[293]);
	Full_Adder FA271 (pp56[9], pp57[8], pp58[7], S[294], Cout[294]);
	Full_Adder FA272 (pp59[6], pp60[5], pp61[4], S[295], Cout[295]);
	Full_Adder FA273 (pp62[3], pp63[2], Cout[2], S[296], Cout[296]);
	Full_Adder FA274 (pp3[63], pp4[62], pp5[61], S[297], Cout[297]);
	Full_Adder FA275 (pp6[60], pp7[59], pp8[58], S[298], Cout[298]);
	Full_Adder FA276 (pp9[57], pp10[56], pp11[55], S[299], Cout[299]);
	Full_Adder FA277 (pp12[54], pp13[53], pp14[52], S[300], Cout[300]);
	Full_Adder FA278 (pp15[51], pp16[50], pp17[49], S[301], Cout[301]);
	Full_Adder FA279 (pp18[48], pp19[47], pp20[46], S[302], Cout[302]);
	Full_Adder FA280 (pp21[45], pp22[44], pp23[43], S[303], Cout[303]);
	Full_Adder FA281 (pp24[42], pp25[41], pp26[40], S[304], Cout[304]);
	Full_Adder FA282 (pp27[39], pp28[38], pp29[37], S[305], Cout[305]);
	Full_Adder FA283 (pp30[36], pp31[35], pp32[34], S[306], Cout[306]);
	Full_Adder FA284 (pp33[33], pp34[32], pp35[31], S[307], Cout[307]);
	Full_Adder FA285 (pp36[30], pp37[29], pp38[28], S[308], Cout[308]);
	Full_Adder FA286 (pp39[27], pp40[26], pp41[25], S[309], Cout[309]);
	Full_Adder FA287 (pp42[24], pp43[23], pp44[22], S[310], Cout[310]);
	Full_Adder FA288 (pp45[21], pp46[20], pp47[19], S[311], Cout[311]);
	Full_Adder FA289 (pp48[18], pp49[17], pp50[16], S[312], Cout[312]);
	Full_Adder FA290 (pp51[15], pp52[14], pp53[13], S[313], Cout[313]);
	Full_Adder FA291 (pp54[12], pp55[11], pp56[10], S[314], Cout[314]);
	Full_Adder FA292 (pp57[9], pp58[8], pp59[7], S[315], Cout[315]);
	Full_Adder FA293 (pp60[6], pp61[5], pp62[4], S[316], Cout[316]);
	Full_Adder FA294 (pp4[63], pp5[62], pp6[61], S[317], Cout[317]);
	Full_Adder FA295 (pp7[60], pp8[59], pp9[58], S[318], Cout[318]);
	Full_Adder FA296 (pp10[57], pp11[56], pp12[55], S[319], Cout[319]);
	Full_Adder FA297 (pp13[54], pp14[53], pp15[52], S[320], Cout[320]);
	Full_Adder FA298 (pp16[51], pp17[50], pp18[49], S[321], Cout[321]);
	Full_Adder FA299 (pp19[48], pp20[47], pp21[46], S[322], Cout[322]);
	Full_Adder FA300 (pp22[45], pp23[44], pp24[43], S[323], Cout[323]);
	Full_Adder FA301 (pp25[42], pp26[41], pp27[40], S[324], Cout[324]);
	Full_Adder FA302 (pp28[39], pp29[38], pp30[37], S[325], Cout[325]);
	Full_Adder FA303 (pp31[36], pp32[35], pp33[34], S[326], Cout[326]);
	Full_Adder FA304 (pp34[33], pp35[32], pp36[31], S[327], Cout[327]);
	Full_Adder FA305 (pp37[30], pp38[29], pp39[28], S[328], Cout[328]);
	Full_Adder FA306 (pp40[27], pp41[26], pp42[25], S[329], Cout[329]);
	Full_Adder FA307 (pp43[24], pp44[23], pp45[22], S[330], Cout[330]);
	Full_Adder FA308 (pp46[21], pp47[20], pp48[19], S[331], Cout[331]);
	Full_Adder FA309 (pp49[18], pp50[17], pp51[16], S[332], Cout[332]);
	Full_Adder FA310 (pp52[15], pp53[14], pp54[13], S[333], Cout[333]);
	Full_Adder FA311 (pp55[12], pp56[11], pp57[10], S[334], Cout[334]);
	Full_Adder FA312 (pp58[9], pp59[8], pp60[7], S[335], Cout[335]);
	Full_Adder FA313 (pp5[63], pp6[62], pp7[61], S[336], Cout[336]);
	Full_Adder FA314 (pp8[60], pp9[59], pp10[58], S[337], Cout[337]);
	Full_Adder FA315 (pp11[57], pp12[56], pp13[55], S[338], Cout[338]);
	Full_Adder FA316 (pp14[54], pp15[53], pp16[52], S[339], Cout[339]);
	Full_Adder FA317 (pp17[51], pp18[50], pp19[49], S[340], Cout[340]);
	Full_Adder FA318 (pp20[48], pp21[47], pp22[46], S[341], Cout[341]);
	Full_Adder FA319 (pp23[45], pp24[44], pp25[43], S[342], Cout[342]);
	Full_Adder FA320 (pp26[42], pp27[41], pp28[40], S[343], Cout[343]);
	Full_Adder FA321 (pp29[39], pp30[38], pp31[37], S[344], Cout[344]);
	Full_Adder FA322 (pp32[36], pp33[35], pp34[34], S[345], Cout[345]);
	Full_Adder FA323 (pp35[33], pp36[32], pp37[31], S[346], Cout[346]);
	Full_Adder FA324 (pp38[30], pp39[29], pp40[28], S[347], Cout[347]);
	Full_Adder FA325 (pp41[27], pp42[26], pp43[25], S[348], Cout[348]);
	Full_Adder FA326 (pp44[24], pp45[23], pp46[22], S[349], Cout[349]);
	Full_Adder FA327 (pp47[21], pp48[20], pp49[19], S[350], Cout[350]);
	Full_Adder FA328 (pp50[18], pp51[17], pp52[16], S[351], Cout[351]);
	Full_Adder FA329 (pp53[15], pp54[14], pp55[13], S[352], Cout[352]);
	Full_Adder FA330 (pp56[12], pp57[11], pp58[10], S[353], Cout[353]);
	Full_Adder FA331 (pp6[63], pp7[62], pp8[61], S[354], Cout[354]);
	Full_Adder FA332 (pp9[60], pp10[59], pp11[58], S[355], Cout[355]);
	Full_Adder FA333 (pp12[57], pp13[56], pp14[55], S[356], Cout[356]);
	Full_Adder FA334 (pp15[54], pp16[53], pp17[52], S[357], Cout[357]);
	Full_Adder FA335 (pp18[51], pp19[50], pp20[49], S[358], Cout[358]);
	Full_Adder FA336 (pp21[48], pp22[47], pp23[46], S[359], Cout[359]);
	Full_Adder FA337 (pp24[45], pp25[44], pp26[43], S[360], Cout[360]);
	Full_Adder FA338 (pp27[42], pp28[41], pp29[40], S[361], Cout[361]);
	Full_Adder FA339 (pp30[39], pp31[38], pp32[37], S[362], Cout[362]);
	Full_Adder FA340 (pp33[36], pp34[35], pp35[34], S[363], Cout[363]);
	Full_Adder FA341 (pp36[33], pp37[32], pp38[31], S[364], Cout[364]);
	Full_Adder FA342 (pp39[30], pp40[29], pp41[28], S[365], Cout[365]);
	Full_Adder FA343 (pp42[27], pp43[26], pp44[25], S[366], Cout[366]);
	Full_Adder FA344 (pp45[24], pp46[23], pp47[22], S[367], Cout[367]);
	Full_Adder FA345 (pp48[21], pp49[20], pp50[19], S[368], Cout[368]);
	Full_Adder FA346 (pp51[18], pp52[17], pp53[16], S[369], Cout[369]);
	Full_Adder FA347 (pp54[15], pp55[14], pp56[13], S[370], Cout[370]);
	Full_Adder FA348 (pp7[63], pp8[62], pp9[61], S[371], Cout[371]);
	Full_Adder FA349 (pp10[60], pp11[59], pp12[58], S[372], Cout[372]);
	Full_Adder FA350 (pp13[57], pp14[56], pp15[55], S[373], Cout[373]);
	Full_Adder FA351 (pp16[54], pp17[53], pp18[52], S[374], Cout[374]);
	Full_Adder FA352 (pp19[51], pp20[50], pp21[49], S[375], Cout[375]);
	Full_Adder FA353 (pp22[48], pp23[47], pp24[46], S[376], Cout[376]);
	Full_Adder FA354 (pp25[45], pp26[44], pp27[43], S[377], Cout[377]);
	Full_Adder FA355 (pp28[42], pp29[41], pp30[40], S[378], Cout[378]);
	Full_Adder FA356 (pp31[39], pp32[38], pp33[37], S[379], Cout[379]);
	Full_Adder FA357 (pp34[36], pp35[35], pp36[34], S[380], Cout[380]);
	Full_Adder FA358 (pp37[33], pp38[32], pp39[31], S[381], Cout[381]);
	Full_Adder FA359 (pp40[30], pp41[29], pp42[28], S[382], Cout[382]);
	Full_Adder FA360 (pp43[27], pp44[26], pp45[25], S[383], Cout[383]);
	Full_Adder FA361 (pp46[24], pp47[23], pp48[22], S[384], Cout[384]);
	Full_Adder FA362 (pp49[21], pp50[20], pp51[19], S[385], Cout[385]);
	Full_Adder FA363 (pp52[18], pp53[17], pp54[16], S[386], Cout[386]);
	Full_Adder FA364 (pp8[63], pp9[62], pp10[61], S[387], Cout[387]);
	Full_Adder FA365 (pp11[60], pp12[59], pp13[58], S[388], Cout[388]);
	Full_Adder FA366 (pp14[57], pp15[56], pp16[55], S[389], Cout[389]);
	Full_Adder FA367 (pp17[54], pp18[53], pp19[52], S[390], Cout[390]);
	Full_Adder FA368 (pp20[51], pp21[50], pp22[49], S[391], Cout[391]);
	Full_Adder FA369 (pp23[48], pp24[47], pp25[46], S[392], Cout[392]);
	Full_Adder FA370 (pp26[45], pp27[44], pp28[43], S[393], Cout[393]);
	Full_Adder FA371 (pp29[42], pp30[41], pp31[40], S[394], Cout[394]);
	Full_Adder FA372 (pp32[39], pp33[38], pp34[37], S[395], Cout[395]);
	Full_Adder FA373 (pp35[36], pp36[35], pp37[34], S[396], Cout[396]);
	Full_Adder FA374 (pp38[33], pp39[32], pp40[31], S[397], Cout[397]);
	Full_Adder FA375 (pp41[30], pp42[29], pp43[28], S[398], Cout[398]);
	Full_Adder FA376 (pp44[27], pp45[26], pp46[25], S[399], Cout[399]);
	Full_Adder FA377 (pp47[24], pp48[23], pp49[22], S[400], Cout[400]);
	Full_Adder FA378 (pp50[21], pp51[20], pp52[19], S[401], Cout[401]);
	Full_Adder FA379 (pp9[63], pp10[62], pp11[61], S[402], Cout[402]);
	Full_Adder FA380 (pp12[60], pp13[59], pp14[58], S[403], Cout[403]);
	Full_Adder FA381 (pp15[57], pp16[56], pp17[55], S[404], Cout[404]);
	Full_Adder FA382 (pp18[54], pp19[53], pp20[52], S[405], Cout[405]);
	Full_Adder FA383 (pp21[51], pp22[50], pp23[49], S[406], Cout[406]);
	Full_Adder FA384 (pp24[48], pp25[47], pp26[46], S[407], Cout[407]);
	Full_Adder FA385 (pp27[45], pp28[44], pp29[43], S[408], Cout[408]);
	Full_Adder FA386 (pp30[42], pp31[41], pp32[40], S[409], Cout[409]);
	Full_Adder FA387 (pp33[39], pp34[38], pp35[37], S[410], Cout[410]);
	Full_Adder FA388 (pp36[36], pp37[35], pp38[34], S[411], Cout[411]);
	Full_Adder FA389 (pp39[33], pp40[32], pp41[31], S[412], Cout[412]);
	Full_Adder FA390 (pp42[30], pp43[29], pp44[28], S[413], Cout[413]);
	Full_Adder FA391 (pp45[27], pp46[26], pp47[25], S[414], Cout[414]);
	Full_Adder FA392 (pp48[24], pp49[23], pp50[22], S[415], Cout[415]);
	Full_Adder FA393 (pp10[63], pp11[62], pp12[61], S[416], Cout[416]);
	Full_Adder FA394 (pp13[60], pp14[59], pp15[58], S[417], Cout[417]);
	Full_Adder FA395 (pp16[57], pp17[56], pp18[55], S[418], Cout[418]);
	Full_Adder FA396 (pp19[54], pp20[53], pp21[52], S[419], Cout[419]);
	Full_Adder FA397 (pp22[51], pp23[50], pp24[49], S[420], Cout[420]);
	Full_Adder FA398 (pp25[48], pp26[47], pp27[46], S[421], Cout[421]);
	Full_Adder FA399 (pp28[45], pp29[44], pp30[43], S[422], Cout[422]);
	Full_Adder FA400 (pp31[42], pp32[41], pp33[40], S[423], Cout[423]);
	Full_Adder FA401 (pp34[39], pp35[38], pp36[37], S[424], Cout[424]);
	Full_Adder FA402 (pp37[36], pp38[35], pp39[34], S[425], Cout[425]);
	Full_Adder FA403 (pp40[33], pp41[32], pp42[31], S[426], Cout[426]);
	Full_Adder FA404 (pp43[30], pp44[29], pp45[28], S[427], Cout[427]);
	Full_Adder FA405 (pp46[27], pp47[26], pp48[25], S[428], Cout[428]);
	Full_Adder FA406 (pp11[63], pp12[62], pp13[61], S[429], Cout[429]);
	Full_Adder FA407 (pp14[60], pp15[59], pp16[58], S[430], Cout[430]);
	Full_Adder FA408 (pp17[57], pp18[56], pp19[55], S[431], Cout[431]);
	Full_Adder FA409 (pp20[54], pp21[53], pp22[52], S[432], Cout[432]);
	Full_Adder FA410 (pp23[51], pp24[50], pp25[49], S[433], Cout[433]);
	Full_Adder FA411 (pp26[48], pp27[47], pp28[46], S[434], Cout[434]);
	Full_Adder FA412 (pp29[45], pp30[44], pp31[43], S[435], Cout[435]);
	Full_Adder FA413 (pp32[42], pp33[41], pp34[40], S[436], Cout[436]);
	Full_Adder FA414 (pp35[39], pp36[38], pp37[37], S[437], Cout[437]);
	Full_Adder FA415 (pp38[36], pp39[35], pp40[34], S[438], Cout[438]);
	Full_Adder FA416 (pp41[33], pp42[32], pp43[31], S[439], Cout[439]);
	Full_Adder FA417 (pp44[30], pp45[29], pp46[28], S[440], Cout[440]);
	Full_Adder FA418 (pp12[63], pp13[62], pp14[61], S[441], Cout[441]);
	Full_Adder FA419 (pp15[60], pp16[59], pp17[58], S[442], Cout[442]);
	Full_Adder FA420 (pp18[57], pp19[56], pp20[55], S[443], Cout[443]);
	Full_Adder FA421 (pp21[54], pp22[53], pp23[52], S[444], Cout[444]);
	Full_Adder FA422 (pp24[51], pp25[50], pp26[49], S[445], Cout[445]);
	Full_Adder FA423 (pp27[48], pp28[47], pp29[46], S[446], Cout[446]);
	Full_Adder FA424 (pp30[45], pp31[44], pp32[43], S[447], Cout[447]);
	Full_Adder FA425 (pp33[42], pp34[41], pp35[40], S[448], Cout[448]);
	Full_Adder FA426 (pp36[39], pp37[38], pp38[37], S[449], Cout[449]);
	Full_Adder FA427 (pp39[36], pp40[35], pp41[34], S[450], Cout[450]);
	Full_Adder FA428 (pp42[33], pp43[32], pp44[31], S[451], Cout[451]);
	Full_Adder FA429 (pp13[63], pp14[62], pp15[61], S[452], Cout[452]);
	Full_Adder FA430 (pp16[60], pp17[59], pp18[58], S[453], Cout[453]);
	Full_Adder FA431 (pp19[57], pp20[56], pp21[55], S[454], Cout[454]);
	Full_Adder FA432 (pp22[54], pp23[53], pp24[52], S[455], Cout[455]);
	Full_Adder FA433 (pp25[51], pp26[50], pp27[49], S[456], Cout[456]);
	Full_Adder FA434 (pp28[48], pp29[47], pp30[46], S[457], Cout[457]);
	Full_Adder FA435 (pp31[45], pp32[44], pp33[43], S[458], Cout[458]);
	Full_Adder FA436 (pp34[42], pp35[41], pp36[40], S[459], Cout[459]);
	Full_Adder FA437 (pp37[39], pp38[38], pp39[37], S[460], Cout[460]);
	Full_Adder FA438 (pp40[36], pp41[35], pp42[34], S[461], Cout[461]);
	Full_Adder FA439 (pp14[63], pp15[62], pp16[61], S[462], Cout[462]);
	Full_Adder FA440 (pp17[60], pp18[59], pp19[58], S[463], Cout[463]);
	Full_Adder FA441 (pp20[57], pp21[56], pp22[55], S[464], Cout[464]);
	Full_Adder FA442 (pp23[54], pp24[53], pp25[52], S[465], Cout[465]);
	Full_Adder FA443 (pp26[51], pp27[50], pp28[49], S[466], Cout[466]);
	Full_Adder FA444 (pp29[48], pp30[47], pp31[46], S[467], Cout[467]);
	Full_Adder FA445 (pp32[45], pp33[44], pp34[43], S[468], Cout[468]);
	Full_Adder FA446 (pp35[42], pp36[41], pp37[40], S[469], Cout[469]);
	Full_Adder FA447 (pp38[39], pp39[38], pp40[37], S[470], Cout[470]);
	Full_Adder FA448 (pp15[63], pp16[62], pp17[61], S[471], Cout[471]);
	Full_Adder FA449 (pp18[60], pp19[59], pp20[58], S[472], Cout[472]);
	Full_Adder FA450 (pp21[57], pp22[56], pp23[55], S[473], Cout[473]);
	Full_Adder FA451 (pp24[54], pp25[53], pp26[52], S[474], Cout[474]);
	Full_Adder FA452 (pp27[51], pp28[50], pp29[49], S[475], Cout[475]);
	Full_Adder FA453 (pp30[48], pp31[47], pp32[46], S[476], Cout[476]);
	Full_Adder FA454 (pp33[45], pp34[44], pp35[43], S[477], Cout[477]);
	Full_Adder FA455 (pp36[42], pp37[41], pp38[40], S[478], Cout[478]);
	Full_Adder FA456 (pp16[63], pp17[62], pp18[61], S[479], Cout[479]);
	Full_Adder FA457 (pp19[60], pp20[59], pp21[58], S[480], Cout[480]);
	Full_Adder FA458 (pp22[57], pp23[56], pp24[55], S[481], Cout[481]);
	Full_Adder FA459 (pp25[54], pp26[53], pp27[52], S[482], Cout[482]);
	Full_Adder FA460 (pp28[51], pp29[50], pp30[49], S[483], Cout[483]);
	Full_Adder FA461 (pp31[48], pp32[47], pp33[46], S[484], Cout[484]);
	Full_Adder FA462 (pp34[45], pp35[44], pp36[43], S[485], Cout[485]);
	Full_Adder FA463 (pp17[63], pp18[62], pp19[61], S[486], Cout[486]);
	Full_Adder FA464 (pp20[60], pp21[59], pp22[58], S[487], Cout[487]);
	Full_Adder FA465 (pp23[57], pp24[56], pp25[55], S[488], Cout[488]);
	Full_Adder FA466 (pp26[54], pp27[53], pp28[52], S[489], Cout[489]);
	Full_Adder FA467 (pp29[51], pp30[50], pp31[49], S[490], Cout[490]);
	Full_Adder FA468 (pp32[48], pp33[47], pp34[46], S[491], Cout[491]);
	Full_Adder FA469 (pp18[63], pp19[62], pp20[61], S[492], Cout[492]);
	Full_Adder FA470 (pp21[60], pp22[59], pp23[58], S[493], Cout[493]);
	Full_Adder FA471 (pp24[57], pp25[56], pp26[55], S[494], Cout[494]);
	Full_Adder FA472 (pp27[54], pp28[53], pp29[52], S[495], Cout[495]);
	Full_Adder FA473 (pp30[51], pp31[50], pp32[49], S[496], Cout[496]);
	Full_Adder FA474 (pp19[63], pp20[62], pp21[61], S[497], Cout[497]);
	Full_Adder FA475 (pp22[60], pp23[59], pp24[58], S[498], Cout[498]);
	Full_Adder FA476 (pp25[57], pp26[56], pp27[55], S[499], Cout[499]);
	Full_Adder FA477 (pp28[54], pp29[53], pp30[52], S[500], Cout[500]);
	Full_Adder FA478 (pp20[63], pp21[62], pp22[61], S[501], Cout[501]);
	Full_Adder FA479 (pp23[60], pp24[59], pp25[58], S[502], Cout[502]);
	Full_Adder FA480 (pp26[57], pp27[56], pp28[55], S[503], Cout[503]);
	Full_Adder FA481 (pp21[63], pp22[62], pp23[61], S[504], Cout[504]);
	Full_Adder FA482 (pp24[60], pp25[59], pp26[58], S[505], Cout[505]);
	Full_Adder FA483 (pp22[63], pp23[62], pp24[61], S[506], Cout[506]);
	Half_Adder HA24 (pp0[28], pp1[27], S[507], Cout[507]);
	Full_Adder FA484 (pp0[29], pp1[28], pp2[27], S[508], Cout[508]);
	Half_Adder HA25 (pp3[26], pp4[25], S[509], Cout[509]);
	Full_Adder FA485 (pp0[30], pp1[29], pp2[28], S[510], Cout[510]);
	Full_Adder FA486 (pp3[27], pp4[26], pp5[25], S[511], Cout[511]);
	Half_Adder HA26 (pp6[24], pp7[23], S[512], Cout[512]);
	Full_Adder FA487 (pp0[31], pp1[30], pp2[29], S[513], Cout[513]);
	Full_Adder FA488 (pp3[28], pp4[27], pp5[26], S[514], Cout[514]);
	Full_Adder FA489 (pp6[25], pp7[24], pp8[23], S[515], Cout[515]);
	Half_Adder HA27 (pp9[22], pp10[21], S[516], Cout[516]);
	Full_Adder FA490 (pp0[32], pp1[31], pp2[30], S[517], Cout[517]);
	Full_Adder FA491 (pp3[29], pp4[28], pp5[27], S[518], Cout[518]);
	Full_Adder FA492 (pp6[26], pp7[25], pp8[24], S[519], Cout[519]);
	Full_Adder FA493 (pp9[23], pp10[22], pp11[21], S[520], Cout[520]);
	Half_Adder HA28 (pp12[20], pp13[19], S[521], Cout[521]);
	Full_Adder FA494 (pp0[33], pp1[32], pp2[31], S[522], Cout[522]);
	Full_Adder FA495 (pp3[30], pp4[29], pp5[28], S[523], Cout[523]);
	Full_Adder FA496 (pp6[27], pp7[26], pp8[25], S[524], Cout[524]);
	Full_Adder FA497 (pp9[24], pp10[23], pp11[22], S[525], Cout[525]);
	Full_Adder FA498 (pp12[21], pp13[20], pp14[19], S[526], Cout[526]);
	Half_Adder HA29 (pp15[18], pp16[17], S[527], Cout[527]);
	Full_Adder FA499 (pp0[34], pp1[33], pp2[32], S[528], Cout[528]);
	Full_Adder FA500 (pp3[31], pp4[30], pp5[29], S[529], Cout[529]);
	Full_Adder FA501 (pp6[28], pp7[27], pp8[26], S[530], Cout[530]);
	Full_Adder FA502 (pp9[25], pp10[24], pp11[23], S[531], Cout[531]);
	Full_Adder FA503 (pp12[22], pp13[21], pp14[20], S[532], Cout[532]);
	Full_Adder FA504 (pp15[19], pp16[18], pp17[17], S[533], Cout[533]);
	Half_Adder HA30 (pp18[16], pp19[15], S[534], Cout[534]);
	Full_Adder FA505 (pp0[35], pp1[34], pp2[33], S[535], Cout[535]);
	Full_Adder FA506 (pp3[32], pp4[31], pp5[30], S[536], Cout[536]);
	Full_Adder FA507 (pp6[29], pp7[28], pp8[27], S[537], Cout[537]);
	Full_Adder FA508 (pp9[26], pp10[25], pp11[24], S[538], Cout[538]);
	Full_Adder FA509 (pp12[23], pp13[22], pp14[21], S[539], Cout[539]);
	Full_Adder FA510 (pp15[20], pp16[19], pp17[18], S[540], Cout[540]);
	Full_Adder FA511 (pp18[17], pp19[16], pp20[15], S[541], Cout[541]);
	Half_Adder HA31 (pp21[14], pp22[13], S[542], Cout[542]);
	Full_Adder FA512 (pp0[36], pp1[35], pp2[34], S[543], Cout[543]);
	Full_Adder FA513 (pp3[33], pp4[32], pp5[31], S[544], Cout[544]);
	Full_Adder FA514 (pp6[30], pp7[29], pp8[28], S[545], Cout[545]);
	Full_Adder FA515 (pp9[27], pp10[26], pp11[25], S[546], Cout[546]);
	Full_Adder FA516 (pp12[24], pp13[23], pp14[22], S[547], Cout[547]);
	Full_Adder FA517 (pp15[21], pp16[20], pp17[19], S[548], Cout[548]);
	Full_Adder FA518 (pp18[18], pp19[17], pp20[16], S[549], Cout[549]);
	Full_Adder FA519 (pp21[15], pp22[14], pp23[13], S[550], Cout[550]);
	Half_Adder HA32 (pp24[12], pp25[11], S[551], Cout[551]);
	Full_Adder FA520 (pp0[37], pp1[36], pp2[35], S[552], Cout[552]);
	Full_Adder FA521 (pp3[34], pp4[33], pp5[32], S[553], Cout[553]);
	Full_Adder FA522 (pp6[31], pp7[30], pp8[29], S[554], Cout[554]);
	Full_Adder FA523 (pp9[28], pp10[27], pp11[26], S[555], Cout[555]);
	Full_Adder FA524 (pp12[25], pp13[24], pp14[23], S[556], Cout[556]);
	Full_Adder FA525 (pp15[22], pp16[21], pp17[20], S[557], Cout[557]);
	Full_Adder FA526 (pp18[19], pp19[18], pp20[17], S[558], Cout[558]);
	Full_Adder FA527 (pp21[16], pp22[15], pp23[14], S[559], Cout[559]);
	Full_Adder FA528 (pp24[13], pp25[12], pp26[11], S[560], Cout[560]);
	Half_Adder HA33 (pp27[10], pp28[9], S[561], Cout[561]);
	Full_Adder FA529 (pp0[38], pp1[37], pp2[36], S[562], Cout[562]);
	Full_Adder FA530 (pp3[35], pp4[34], pp5[33], S[563], Cout[563]);
	Full_Adder FA531 (pp6[32], pp7[31], pp8[30], S[564], Cout[564]);
	Full_Adder FA532 (pp9[29], pp10[28], pp11[27], S[565], Cout[565]);
	Full_Adder FA533 (pp12[26], pp13[25], pp14[24], S[566], Cout[566]);
	Full_Adder FA534 (pp15[23], pp16[22], pp17[21], S[567], Cout[567]);
	Full_Adder FA535 (pp18[20], pp19[19], pp20[18], S[568], Cout[568]);
	Full_Adder FA536 (pp21[17], pp22[16], pp23[15], S[569], Cout[569]);
	Full_Adder FA537 (pp24[14], pp25[13], pp26[12], S[570], Cout[570]);
	Full_Adder FA538 (pp27[11], pp28[10], pp29[9], S[571], Cout[571]);
	Half_Adder HA34 (pp30[8], pp31[7], S[572], Cout[572]);
	Full_Adder FA539 (pp0[39], pp1[38], pp2[37], S[573], Cout[573]);
	Full_Adder FA540 (pp3[36], pp4[35], pp5[34], S[574], Cout[574]);
	Full_Adder FA541 (pp6[33], pp7[32], pp8[31], S[575], Cout[575]);
	Full_Adder FA542 (pp9[30], pp10[29], pp11[28], S[576], Cout[576]);
	Full_Adder FA543 (pp12[27], pp13[26], pp14[25], S[577], Cout[577]);
	Full_Adder FA544 (pp15[24], pp16[23], pp17[22], S[578], Cout[578]);
	Full_Adder FA545 (pp18[21], pp19[20], pp20[19], S[579], Cout[579]);
	Full_Adder FA546 (pp21[18], pp22[17], pp23[16], S[580], Cout[580]);
	Full_Adder FA547 (pp24[15], pp25[14], pp26[13], S[581], Cout[581]);
	Full_Adder FA548 (pp27[12], pp28[11], pp29[10], S[582], Cout[582]);
	Full_Adder FA549 (pp30[9], pp31[8], pp32[7], S[583], Cout[583]);
	Half_Adder HA35 (pp33[6], pp34[5], S[584], Cout[584]);
	Full_Adder FA550 (pp0[40], pp1[39], pp2[38], S[585], Cout[585]);
	Full_Adder FA551 (pp3[37], pp4[36], pp5[35], S[586], Cout[586]);
	Full_Adder FA552 (pp6[34], pp7[33], pp8[32], S[587], Cout[587]);
	Full_Adder FA553 (pp9[31], pp10[30], pp11[29], S[588], Cout[588]);
	Full_Adder FA554 (pp12[28], pp13[27], pp14[26], S[589], Cout[589]);
	Full_Adder FA555 (pp15[25], pp16[24], pp17[23], S[590], Cout[590]);
	Full_Adder FA556 (pp18[22], pp19[21], pp20[20], S[591], Cout[591]);
	Full_Adder FA557 (pp21[19], pp22[18], pp23[17], S[592], Cout[592]);
	Full_Adder FA558 (pp24[16], pp25[15], pp26[14], S[593], Cout[593]);
	Full_Adder FA559 (pp27[13], pp28[12], pp29[11], S[594], Cout[594]);
	Full_Adder FA560 (pp30[10], pp31[9], pp32[8], S[595], Cout[595]);
	Full_Adder FA561 (pp33[7], pp34[6], pp35[5], S[596], Cout[596]);
	Half_Adder HA36 (pp36[4], pp37[3], S[597], Cout[597]);
	Full_Adder FA562 (pp0[41], pp1[40], pp2[39], S[598], Cout[598]);
	Full_Adder FA563 (pp3[38], pp4[37], pp5[36], S[599], Cout[599]);
	Full_Adder FA564 (pp6[35], pp7[34], pp8[33], S[600], Cout[600]);
	Full_Adder FA565 (pp9[32], pp10[31], pp11[30], S[601], Cout[601]);
	Full_Adder FA566 (pp12[29], pp13[28], pp14[27], S[602], Cout[602]);
	Full_Adder FA567 (pp15[26], pp16[25], pp17[24], S[603], Cout[603]);
	Full_Adder FA568 (pp18[23], pp19[22], pp20[21], S[604], Cout[604]);
	Full_Adder FA569 (pp21[20], pp22[19], pp23[18], S[605], Cout[605]);
	Full_Adder FA570 (pp24[17], pp25[16], pp26[15], S[606], Cout[606]);
	Full_Adder FA571 (pp27[14], pp28[13], pp29[12], S[607], Cout[607]);
	Full_Adder FA572 (pp30[11], pp31[10], pp32[9], S[608], Cout[608]);
	Full_Adder FA573 (pp33[8], pp34[7], pp35[6], S[609], Cout[609]);
	Full_Adder FA574 (pp36[5], pp37[4], pp38[3], S[610], Cout[610]);
	Half_Adder HA37 (pp39[2], pp40[1], S[611], Cout[611]);
	Full_Adder FA575 (pp2[40], pp3[39], pp4[38], S[612], Cout[612]);
	Full_Adder FA576 (pp5[37], pp6[36], pp7[35], S[613], Cout[613]);
	Full_Adder FA577 (pp8[34], pp9[33], pp10[32], S[614], Cout[614]);
	Full_Adder FA578 (pp11[31], pp12[30], pp13[29], S[615], Cout[615]);
	Full_Adder FA579 (pp14[28], pp15[27], pp16[26], S[616], Cout[616]);
	Full_Adder FA580 (pp17[25], pp18[24], pp19[23], S[617], Cout[617]);
	Full_Adder FA581 (pp20[22], pp21[21], pp22[20], S[618], Cout[618]);
	Full_Adder FA582 (pp23[19], pp24[18], pp25[17], S[619], Cout[619]);
	Full_Adder FA583 (pp26[16], pp27[15], pp28[14], S[620], Cout[620]);
	Full_Adder FA584 (pp29[13], pp30[12], pp31[11], S[621], Cout[621]);
	Full_Adder FA585 (pp32[10], pp33[9], pp34[8], S[622], Cout[622]);
	Full_Adder FA586 (pp35[7], pp36[6], pp37[5], S[623], Cout[623]);
	Full_Adder FA587 (pp38[4], pp39[3], pp40[2], S[624], Cout[624]);
	Full_Adder FA588 (pp41[1], pp42[0], S[3], S[625], Cout[625]);
	Full_Adder FA589 (pp5[38], pp6[37], pp7[36], S[626], Cout[626]);
	Full_Adder FA590 (pp8[35], pp9[34], pp10[33], S[627], Cout[627]);
	Full_Adder FA591 (pp11[32], pp12[31], pp13[30], S[628], Cout[628]);
	Full_Adder FA592 (pp14[29], pp15[28], pp16[27], S[629], Cout[629]);
	Full_Adder FA593 (pp17[26], pp18[25], pp19[24], S[630], Cout[630]);
	Full_Adder FA594 (pp20[23], pp21[22], pp22[21], S[631], Cout[631]);
	Full_Adder FA595 (pp23[20], pp24[19], pp25[18], S[632], Cout[632]);
	Full_Adder FA596 (pp26[17], pp27[16], pp28[15], S[633], Cout[633]);
	Full_Adder FA597 (pp29[14], pp30[13], pp31[12], S[634], Cout[634]);
	Full_Adder FA598 (pp32[11], pp33[10], pp34[9], S[635], Cout[635]);
	Full_Adder FA599 (pp35[8], pp36[7], pp37[6], S[636], Cout[636]);
	Full_Adder FA600 (pp38[5], pp39[4], pp40[3], S[637], Cout[637]);
	Full_Adder FA601 (pp41[2], pp42[1], pp43[0], S[638], Cout[638]);
	Full_Adder FA602 (Cout[3], S[4], S[5], S[639], Cout[639]);
	Full_Adder FA603 (pp8[36], pp9[35], pp10[34], S[640], Cout[640]);
	Full_Adder FA604 (pp11[33], pp12[32], pp13[31], S[641], Cout[641]);
	Full_Adder FA605 (pp14[30], pp15[29], pp16[28], S[642], Cout[642]);
	Full_Adder FA606 (pp17[27], pp18[26], pp19[25], S[643], Cout[643]);
	Full_Adder FA607 (pp20[24], pp21[23], pp22[22], S[644], Cout[644]);
	Full_Adder FA608 (pp23[21], pp24[20], pp25[19], S[645], Cout[645]);
	Full_Adder FA609 (pp26[18], pp27[17], pp28[16], S[646], Cout[646]);
	Full_Adder FA610 (pp29[15], pp30[14], pp31[13], S[647], Cout[647]);
	Full_Adder FA611 (pp32[12], pp33[11], pp34[10], S[648], Cout[648]);
	Full_Adder FA612 (pp35[9], pp36[8], pp37[7], S[649], Cout[649]);
	Full_Adder FA613 (pp38[6], pp39[5], pp40[4], S[650], Cout[650]);
	Full_Adder FA614 (pp41[3], pp42[2], pp43[1], S[651], Cout[651]);
	Full_Adder FA615 (pp44[0], Cout[4], Cout[5], S[652], Cout[652]);
	Full_Adder FA616 (S[6], S[7], S[8], S[653], Cout[653]);
	Full_Adder FA617 (pp11[34], pp12[33], pp13[32], S[654], Cout[654]);
	Full_Adder FA618 (pp14[31], pp15[30], pp16[29], S[655], Cout[655]);
	Full_Adder FA619 (pp17[28], pp18[27], pp19[26], S[656], Cout[656]);
	Full_Adder FA620 (pp20[25], pp21[24], pp22[23], S[657], Cout[657]);
	Full_Adder FA621 (pp23[22], pp24[21], pp25[20], S[658], Cout[658]);
	Full_Adder FA622 (pp26[19], pp27[18], pp28[17], S[659], Cout[659]);
	Full_Adder FA623 (pp29[16], pp30[15], pp31[14], S[660], Cout[660]);
	Full_Adder FA624 (pp32[13], pp33[12], pp34[11], S[661], Cout[661]);
	Full_Adder FA625 (pp35[10], pp36[9], pp37[8], S[662], Cout[662]);
	Full_Adder FA626 (pp38[7], pp39[6], pp40[5], S[663], Cout[663]);
	Full_Adder FA627 (pp41[4], pp42[3], pp43[2], S[664], Cout[664]);
	Full_Adder FA628 (pp44[1], pp45[0], Cout[6], S[665], Cout[665]);
	Full_Adder FA629 (Cout[7], Cout[8], S[9], S[666], Cout[666]);
	Full_Adder FA630 (S[10], S[11], S[12], S[667], Cout[667]);
	Full_Adder FA631 (pp14[32], pp15[31], pp16[30], S[668], Cout[668]);
	Full_Adder FA632 (pp17[29], pp18[28], pp19[27], S[669], Cout[669]);
	Full_Adder FA633 (pp20[26], pp21[25], pp22[24], S[670], Cout[670]);
	Full_Adder FA634 (pp23[23], pp24[22], pp25[21], S[671], Cout[671]);
	Full_Adder FA635 (pp26[20], pp27[19], pp28[18], S[672], Cout[672]);
	Full_Adder FA636 (pp29[17], pp30[16], pp31[15], S[673], Cout[673]);
	Full_Adder FA637 (pp32[14], pp33[13], pp34[12], S[674], Cout[674]);
	Full_Adder FA638 (pp35[11], pp36[10], pp37[9], S[675], Cout[675]);
	Full_Adder FA639 (pp38[8], pp39[7], pp40[6], S[676], Cout[676]);
	Full_Adder FA640 (pp41[5], pp42[4], pp43[3], S[677], Cout[677]);
	Full_Adder FA641 (pp44[2], pp45[1], pp46[0], S[678], Cout[678]);
	Full_Adder FA642 (Cout[9], Cout[10], Cout[11], S[679], Cout[679]);
	Full_Adder FA643 (Cout[12], S[13], S[14], S[680], Cout[680]);
	Full_Adder FA644 (S[15], S[16], S[17], S[681], Cout[681]);
	Full_Adder FA645 (pp17[30], pp18[29], pp19[28], S[682], Cout[682]);
	Full_Adder FA646 (pp20[27], pp21[26], pp22[25], S[683], Cout[683]);
	Full_Adder FA647 (pp23[24], pp24[23], pp25[22], S[684], Cout[684]);
	Full_Adder FA648 (pp26[21], pp27[20], pp28[19], S[685], Cout[685]);
	Full_Adder FA649 (pp29[18], pp30[17], pp31[16], S[686], Cout[686]);
	Full_Adder FA650 (pp32[15], pp33[14], pp34[13], S[687], Cout[687]);
	Full_Adder FA651 (pp35[12], pp36[11], pp37[10], S[688], Cout[688]);
	Full_Adder FA652 (pp38[9], pp39[8], pp40[7], S[689], Cout[689]);
	Full_Adder FA653 (pp41[6], pp42[5], pp43[4], S[690], Cout[690]);
	Full_Adder FA654 (pp44[3], pp45[2], pp46[1], S[691], Cout[691]);
	Full_Adder FA655 (pp47[0], Cout[13], Cout[14], S[692], Cout[692]);
	Full_Adder FA656 (Cout[15], Cout[16], Cout[17], S[693], Cout[693]);
	Full_Adder FA657 (S[18], S[19], S[20], S[694], Cout[694]);
	Full_Adder FA658 (S[21], S[22], S[23], S[695], Cout[695]);
	Full_Adder FA659 (pp20[28], pp21[27], pp22[26], S[696], Cout[696]);
	Full_Adder FA660 (pp23[25], pp24[24], pp25[23], S[697], Cout[697]);
	Full_Adder FA661 (pp26[22], pp27[21], pp28[20], S[698], Cout[698]);
	Full_Adder FA662 (pp29[19], pp30[18], pp31[17], S[699], Cout[699]);
	Full_Adder FA663 (pp32[16], pp33[15], pp34[14], S[700], Cout[700]);
	Full_Adder FA664 (pp35[13], pp36[12], pp37[11], S[701], Cout[701]);
	Full_Adder FA665 (pp38[10], pp39[9], pp40[8], S[702], Cout[702]);
	Full_Adder FA666 (pp41[7], pp42[6], pp43[5], S[703], Cout[703]);
	Full_Adder FA667 (pp44[4], pp45[3], pp46[2], S[704], Cout[704]);
	Full_Adder FA668 (pp47[1], pp48[0], Cout[18], S[705], Cout[705]);
	Full_Adder FA669 (Cout[19], Cout[20], Cout[21], S[706], Cout[706]);
	Full_Adder FA670 (Cout[22], Cout[23], S[24], S[707], Cout[707]);
	Full_Adder FA671 (S[25], S[26], S[27], S[708], Cout[708]);
	Full_Adder FA672 (S[28], S[29], S[30], S[709], Cout[709]);
	Full_Adder FA673 (pp23[26], pp24[25], pp25[24], S[710], Cout[710]);
	Full_Adder FA674 (pp26[23], pp27[22], pp28[21], S[711], Cout[711]);
	Full_Adder FA675 (pp29[20], pp30[19], pp31[18], S[712], Cout[712]);
	Full_Adder FA676 (pp32[17], pp33[16], pp34[15], S[713], Cout[713]);
	Full_Adder FA677 (pp35[14], pp36[13], pp37[12], S[714], Cout[714]);
	Full_Adder FA678 (pp38[11], pp39[10], pp40[9], S[715], Cout[715]);
	Full_Adder FA679 (pp41[8], pp42[7], pp43[6], S[716], Cout[716]);
	Full_Adder FA680 (pp44[5], pp45[4], pp46[3], S[717], Cout[717]);
	Full_Adder FA681 (pp47[2], pp48[1], pp49[0], S[718], Cout[718]);
	Full_Adder FA682 (Cout[24], Cout[25], Cout[26], S[719], Cout[719]);
	Full_Adder FA683 (Cout[27], Cout[28], Cout[29], S[720], Cout[720]);
	Full_Adder FA684 (Cout[30], S[31], S[32], S[721], Cout[721]);
	Full_Adder FA685 (S[33], S[34], S[35], S[722], Cout[722]);
	Full_Adder FA686 (S[36], S[37], S[38], S[723], Cout[723]);
	Full_Adder FA687 (pp26[24], pp27[23], pp28[22], S[724], Cout[724]);
	Full_Adder FA688 (pp29[21], pp30[20], pp31[19], S[725], Cout[725]);
	Full_Adder FA689 (pp32[18], pp33[17], pp34[16], S[726], Cout[726]);
	Full_Adder FA690 (pp35[15], pp36[14], pp37[13], S[727], Cout[727]);
	Full_Adder FA691 (pp38[12], pp39[11], pp40[10], S[728], Cout[728]);
	Full_Adder FA692 (pp41[9], pp42[8], pp43[7], S[729], Cout[729]);
	Full_Adder FA693 (pp44[6], pp45[5], pp46[4], S[730], Cout[730]);
	Full_Adder FA694 (pp47[3], pp48[2], pp49[1], S[731], Cout[731]);
	Full_Adder FA695 (pp50[0], Cout[31], Cout[32], S[732], Cout[732]);
	Full_Adder FA696 (Cout[33], Cout[34], Cout[35], S[733], Cout[733]);
	Full_Adder FA697 (Cout[36], Cout[37], Cout[38], S[734], Cout[734]);
	Full_Adder FA698 (S[39], S[40], S[41], S[735], Cout[735]);
	Full_Adder FA699 (S[42], S[43], S[44], S[736], Cout[736]);
	Full_Adder FA700 (S[45], S[46], S[47], S[737], Cout[737]);
	Full_Adder FA701 (pp29[22], pp30[21], pp31[20], S[738], Cout[738]);
	Full_Adder FA702 (pp32[19], pp33[18], pp34[17], S[739], Cout[739]);
	Full_Adder FA703 (pp35[16], pp36[15], pp37[14], S[740], Cout[740]);
	Full_Adder FA704 (pp38[13], pp39[12], pp40[11], S[741], Cout[741]);
	Full_Adder FA705 (pp41[10], pp42[9], pp43[8], S[742], Cout[742]);
	Full_Adder FA706 (pp44[7], pp45[6], pp46[5], S[743], Cout[743]);
	Full_Adder FA707 (pp47[4], pp48[3], pp49[2], S[744], Cout[744]);
	Full_Adder FA708 (pp50[1], pp51[0], Cout[39], S[745], Cout[745]);
	Full_Adder FA709 (Cout[40], Cout[41], Cout[42], S[746], Cout[746]);
	Full_Adder FA710 (Cout[43], Cout[44], Cout[45], S[747], Cout[747]);
	Full_Adder FA711 (Cout[46], Cout[47], S[48], S[748], Cout[748]);
	Full_Adder FA712 (S[49], S[50], S[51], S[749], Cout[749]);
	Full_Adder FA713 (S[52], S[53], S[54], S[750], Cout[750]);
	Full_Adder FA714 (S[55], S[56], S[57], S[751], Cout[751]);
	Full_Adder FA715 (pp32[20], pp33[19], pp34[18], S[752], Cout[752]);
	Full_Adder FA716 (pp35[17], pp36[16], pp37[15], S[753], Cout[753]);
	Full_Adder FA717 (pp38[14], pp39[13], pp40[12], S[754], Cout[754]);
	Full_Adder FA718 (pp41[11], pp42[10], pp43[9], S[755], Cout[755]);
	Full_Adder FA719 (pp44[8], pp45[7], pp46[6], S[756], Cout[756]);
	Full_Adder FA720 (pp47[5], pp48[4], pp49[3], S[757], Cout[757]);
	Full_Adder FA721 (pp50[2], pp51[1], pp52[0], S[758], Cout[758]);
	Full_Adder FA722 (Cout[48], Cout[49], Cout[50], S[759], Cout[759]);
	Full_Adder FA723 (Cout[51], Cout[52], Cout[53], S[760], Cout[760]);
	Full_Adder FA724 (Cout[54], Cout[55], Cout[56], S[761], Cout[761]);
	Full_Adder FA725 (Cout[57], S[58], S[59], S[762], Cout[762]);
	Full_Adder FA726 (S[60], S[61], S[62], S[763], Cout[763]);
	Full_Adder FA727 (S[63], S[64], S[65], S[764], Cout[764]);
	Full_Adder FA728 (S[66], S[67], S[68], S[765], Cout[765]);
	Full_Adder FA729 (pp35[18], pp36[17], pp37[16], S[766], Cout[766]);
	Full_Adder FA730 (pp38[15], pp39[14], pp40[13], S[767], Cout[767]);
	Full_Adder FA731 (pp41[12], pp42[11], pp43[10], S[768], Cout[768]);
	Full_Adder FA732 (pp44[9], pp45[8], pp46[7], S[769], Cout[769]);
	Full_Adder FA733 (pp47[6], pp48[5], pp49[4], S[770], Cout[770]);
	Full_Adder FA734 (pp50[3], pp51[2], pp52[1], S[771], Cout[771]);
	Full_Adder FA735 (pp53[0], Cout[58], Cout[59], S[772], Cout[772]);
	Full_Adder FA736 (Cout[60], Cout[61], Cout[62], S[773], Cout[773]);
	Full_Adder FA737 (Cout[63], Cout[64], Cout[65], S[774], Cout[774]);
	Full_Adder FA738 (Cout[66], Cout[67], Cout[68], S[775], Cout[775]);
	Full_Adder FA739 (S[69], S[70], S[71], S[776], Cout[776]);
	Full_Adder FA740 (S[72], S[73], S[74], S[777], Cout[777]);
	Full_Adder FA741 (S[75], S[76], S[77], S[778], Cout[778]);
	Full_Adder FA742 (S[78], S[79], S[80], S[779], Cout[779]);
	Full_Adder FA743 (pp38[16], pp39[15], pp40[14], S[780], Cout[780]);
	Full_Adder FA744 (pp41[13], pp42[12], pp43[11], S[781], Cout[781]);
	Full_Adder FA745 (pp44[10], pp45[9], pp46[8], S[782], Cout[782]);
	Full_Adder FA746 (pp47[7], pp48[6], pp49[5], S[783], Cout[783]);
	Full_Adder FA747 (pp50[4], pp51[3], pp52[2], S[784], Cout[784]);
	Full_Adder FA748 (pp53[1], pp54[0], Cout[69], S[785], Cout[785]);
	Full_Adder FA749 (Cout[70], Cout[71], Cout[72], S[786], Cout[786]);
	Full_Adder FA750 (Cout[73], Cout[74], Cout[75], S[787], Cout[787]);
	Full_Adder FA751 (Cout[76], Cout[77], Cout[78], S[788], Cout[788]);
	Full_Adder FA752 (Cout[79], Cout[80], S[81], S[789], Cout[789]);
	Full_Adder FA753 (S[82], S[83], S[84], S[790], Cout[790]);
	Full_Adder FA754 (S[85], S[86], S[87], S[791], Cout[791]);
	Full_Adder FA755 (S[88], S[89], S[90], S[792], Cout[792]);
	Full_Adder FA756 (S[91], S[92], S[93], S[793], Cout[793]);
	Full_Adder FA757 (pp41[14], pp42[13], pp43[12], S[794], Cout[794]);
	Full_Adder FA758 (pp44[11], pp45[10], pp46[9], S[795], Cout[795]);
	Full_Adder FA759 (pp47[8], pp48[7], pp49[6], S[796], Cout[796]);
	Full_Adder FA760 (pp50[5], pp51[4], pp52[3], S[797], Cout[797]);
	Full_Adder FA761 (pp53[2], pp54[1], pp55[0], S[798], Cout[798]);
	Full_Adder FA762 (Cout[81], Cout[82], Cout[83], S[799], Cout[799]);
	Full_Adder FA763 (Cout[84], Cout[85], Cout[86], S[800], Cout[800]);
	Full_Adder FA764 (Cout[87], Cout[88], Cout[89], S[801], Cout[801]);
	Full_Adder FA765 (Cout[90], Cout[91], Cout[92], S[802], Cout[802]);
	Full_Adder FA766 (Cout[93], S[94], S[95], S[803], Cout[803]);
	Full_Adder FA767 (S[96], S[97], S[98], S[804], Cout[804]);
	Full_Adder FA768 (S[99], S[100], S[101], S[805], Cout[805]);
	Full_Adder FA769 (S[102], S[103], S[104], S[806], Cout[806]);
	Full_Adder FA770 (S[105], S[106], S[107], S[807], Cout[807]);
	Full_Adder FA771 (pp44[12], pp45[11], pp46[10], S[808], Cout[808]);
	Full_Adder FA772 (pp47[9], pp48[8], pp49[7], S[809], Cout[809]);
	Full_Adder FA773 (pp50[6], pp51[5], pp52[4], S[810], Cout[810]);
	Full_Adder FA774 (pp53[3], pp54[2], pp55[1], S[811], Cout[811]);
	Full_Adder FA775 (pp56[0], Cout[94], Cout[95], S[812], Cout[812]);
	Full_Adder FA776 (Cout[96], Cout[97], Cout[98], S[813], Cout[813]);
	Full_Adder FA777 (Cout[99], Cout[100], Cout[101], S[814], Cout[814]);
	Full_Adder FA778 (Cout[102], Cout[103], Cout[104], S[815], Cout[815]);
	Full_Adder FA779 (Cout[105], Cout[106], Cout[107], S[816], Cout[816]);
	Full_Adder FA780 (S[108], S[109], S[110], S[817], Cout[817]);
	Full_Adder FA781 (S[111], S[112], S[113], S[818], Cout[818]);
	Full_Adder FA782 (S[114], S[115], S[116], S[819], Cout[819]);
	Full_Adder FA783 (S[117], S[118], S[119], S[820], Cout[820]);
	Full_Adder FA784 (S[120], S[121], S[122], S[821], Cout[821]);
	Full_Adder FA785 (pp47[10], pp48[9], pp49[8], S[822], Cout[822]);
	Full_Adder FA786 (pp50[7], pp51[6], pp52[5], S[823], Cout[823]);
	Full_Adder FA787 (pp53[4], pp54[3], pp55[2], S[824], Cout[824]);
	Full_Adder FA788 (pp56[1], pp57[0], Cout[108], S[825], Cout[825]);
	Full_Adder FA789 (Cout[109], Cout[110], Cout[111], S[826], Cout[826]);
	Full_Adder FA790 (Cout[112], Cout[113], Cout[114], S[827], Cout[827]);
	Full_Adder FA791 (Cout[115], Cout[116], Cout[117], S[828], Cout[828]);
	Full_Adder FA792 (Cout[118], Cout[119], Cout[120], S[829], Cout[829]);
	Full_Adder FA793 (Cout[121], Cout[122], S[123], S[830], Cout[830]);
	Full_Adder FA794 (S[124], S[125], S[126], S[831], Cout[831]);
	Full_Adder FA795 (S[127], S[128], S[129], S[832], Cout[832]);
	Full_Adder FA796 (S[130], S[131], S[132], S[833], Cout[833]);
	Full_Adder FA797 (S[133], S[134], S[135], S[834], Cout[834]);
	Full_Adder FA798 (S[136], S[137], S[138], S[835], Cout[835]);
	Full_Adder FA799 (pp50[8], pp51[7], pp52[6], S[836], Cout[836]);
	Full_Adder FA800 (pp53[5], pp54[4], pp55[3], S[837], Cout[837]);
	Full_Adder FA801 (pp56[2], pp57[1], pp58[0], S[838], Cout[838]);
	Full_Adder FA802 (Cout[123], Cout[124], Cout[125], S[839], Cout[839]);
	Full_Adder FA803 (Cout[126], Cout[127], Cout[128], S[840], Cout[840]);
	Full_Adder FA804 (Cout[129], Cout[130], Cout[131], S[841], Cout[841]);
	Full_Adder FA805 (Cout[132], Cout[133], Cout[134], S[842], Cout[842]);
	Full_Adder FA806 (Cout[135], Cout[136], Cout[137], S[843], Cout[843]);
	Full_Adder FA807 (Cout[138], S[139], S[140], S[844], Cout[844]);
	Full_Adder FA808 (S[141], S[142], S[143], S[845], Cout[845]);
	Full_Adder FA809 (S[144], S[145], S[146], S[846], Cout[846]);
	Full_Adder FA810 (S[147], S[148], S[149], S[847], Cout[847]);
	Full_Adder FA811 (S[150], S[151], S[152], S[848], Cout[848]);
	Full_Adder FA812 (S[153], S[154], S[155], S[849], Cout[849]);
	Full_Adder FA813 (pp53[6], pp54[5], pp55[4], S[850], Cout[850]);
	Full_Adder FA814 (pp56[3], pp57[2], pp58[1], S[851], Cout[851]);
	Full_Adder FA815 (pp59[0], Cout[139], Cout[140], S[852], Cout[852]);
	Full_Adder FA816 (Cout[141], Cout[142], Cout[143], S[853], Cout[853]);
	Full_Adder FA817 (Cout[144], Cout[145], Cout[146], S[854], Cout[854]);
	Full_Adder FA818 (Cout[147], Cout[148], Cout[149], S[855], Cout[855]);
	Full_Adder FA819 (Cout[150], Cout[151], Cout[152], S[856], Cout[856]);
	Full_Adder FA820 (Cout[153], Cout[154], Cout[155], S[857], Cout[857]);
	Full_Adder FA821 (S[156], S[157], S[158], S[858], Cout[858]);
	Full_Adder FA822 (S[159], S[160], S[161], S[859], Cout[859]);
	Full_Adder FA823 (S[162], S[163], S[164], S[860], Cout[860]);
	Full_Adder FA824 (S[165], S[166], S[167], S[861], Cout[861]);
	Full_Adder FA825 (S[168], S[169], S[170], S[862], Cout[862]);
	Full_Adder FA826 (S[171], S[172], S[173], S[863], Cout[863]);
	Full_Adder FA827 (pp56[4], pp57[3], pp58[2], S[864], Cout[864]);
	Full_Adder FA828 (pp59[1], pp60[0], Cout[156], S[865], Cout[865]);
	Full_Adder FA829 (Cout[157], Cout[158], Cout[159], S[866], Cout[866]);
	Full_Adder FA830 (Cout[160], Cout[161], Cout[162], S[867], Cout[867]);
	Full_Adder FA831 (Cout[163], Cout[164], Cout[165], S[868], Cout[868]);
	Full_Adder FA832 (Cout[166], Cout[167], Cout[168], S[869], Cout[869]);
	Full_Adder FA833 (Cout[169], Cout[170], Cout[171], S[870], Cout[870]);
	Full_Adder FA834 (Cout[172], Cout[173], S[174], S[871], Cout[871]);
	Full_Adder FA835 (S[175], S[176], S[177], S[872], Cout[872]);
	Full_Adder FA836 (S[178], S[179], S[180], S[873], Cout[873]);
	Full_Adder FA837 (S[181], S[182], S[183], S[874], Cout[874]);
	Full_Adder FA838 (S[184], S[185], S[186], S[875], Cout[875]);
	Full_Adder FA839 (S[187], S[188], S[189], S[876], Cout[876]);
	Full_Adder FA840 (S[190], S[191], S[192], S[877], Cout[877]);
	Full_Adder FA841 (pp59[2], pp60[1], pp61[0], S[878], Cout[878]);
	Full_Adder FA842 (Cout[174], Cout[175], Cout[176], S[879], Cout[879]);
	Full_Adder FA843 (Cout[177], Cout[178], Cout[179], S[880], Cout[880]);
	Full_Adder FA844 (Cout[180], Cout[181], Cout[182], S[881], Cout[881]);
	Full_Adder FA845 (Cout[183], Cout[184], Cout[185], S[882], Cout[882]);
	Full_Adder FA846 (Cout[186], Cout[187], Cout[188], S[883], Cout[883]);
	Full_Adder FA847 (Cout[189], Cout[190], Cout[191], S[884], Cout[884]);
	Full_Adder FA848 (Cout[192], S[193], S[194], S[885], Cout[885]);
	Full_Adder FA849 (S[195], S[196], S[197], S[886], Cout[886]);
	Full_Adder FA850 (S[198], S[199], S[200], S[887], Cout[887]);
	Full_Adder FA851 (S[201], S[202], S[203], S[888], Cout[888]);
	Full_Adder FA852 (S[204], S[205], S[206], S[889], Cout[889]);
	Full_Adder FA853 (S[207], S[208], S[209], S[890], Cout[890]);
	Full_Adder FA854 (S[210], S[211], S[212], S[891], Cout[891]);
	Full_Adder FA855 (pp62[0], Cout[193], Cout[194], S[892], Cout[892]);
	Full_Adder FA856 (Cout[195], Cout[196], Cout[197], S[893], Cout[893]);
	Full_Adder FA857 (Cout[198], Cout[199], Cout[200], S[894], Cout[894]);
	Full_Adder FA858 (Cout[201], Cout[202], Cout[203], S[895], Cout[895]);
	Full_Adder FA859 (Cout[204], Cout[205], Cout[206], S[896], Cout[896]);
	Full_Adder FA860 (Cout[207], Cout[208], Cout[209], S[897], Cout[897]);
	Full_Adder FA861 (Cout[210], Cout[211], Cout[212], S[898], Cout[898]);
	Full_Adder FA862 (S[213], S[214], S[215], S[899], Cout[899]);
	Full_Adder FA863 (S[216], S[217], S[218], S[900], Cout[900]);
	Full_Adder FA864 (S[219], S[220], S[221], S[901], Cout[901]);
	Full_Adder FA865 (S[222], S[223], S[224], S[902], Cout[902]);
	Full_Adder FA866 (S[225], S[226], S[227], S[903], Cout[903]);
	Full_Adder FA867 (S[228], S[229], S[230], S[904], Cout[904]);
	Full_Adder FA868 (S[231], S[232], S[233], S[905], Cout[905]);
	Full_Adder FA869 (Cout[213], Cout[214], Cout[215], S[906], Cout[906]);
	Full_Adder FA870 (Cout[216], Cout[217], Cout[218], S[907], Cout[907]);
	Full_Adder FA871 (Cout[219], Cout[220], Cout[221], S[908], Cout[908]);
	Full_Adder FA872 (Cout[222], Cout[223], Cout[224], S[909], Cout[909]);
	Full_Adder FA873 (Cout[225], Cout[226], Cout[227], S[910], Cout[910]);
	Full_Adder FA874 (Cout[228], Cout[229], Cout[230], S[911], Cout[911]);
	Full_Adder FA875 (Cout[231], Cout[232], Cout[233], S[912], Cout[912]);
	Full_Adder FA876 (S[234], S[235], S[236], S[913], Cout[913]);
	Full_Adder FA877 (S[237], S[238], S[239], S[914], Cout[914]);
	Full_Adder FA878 (S[240], S[241], S[242], S[915], Cout[915]);
	Full_Adder FA879 (S[243], S[244], S[245], S[916], Cout[916]);
	Full_Adder FA880 (S[246], S[247], S[248], S[917], Cout[917]);
	Full_Adder FA881 (S[249], S[250], S[251], S[918], Cout[918]);
	Full_Adder FA882 (S[252], S[253], S[254], S[919], Cout[919]);
	Full_Adder FA883 (Cout[234], Cout[235], Cout[236], S[920], Cout[920]);
	Full_Adder FA884 (Cout[237], Cout[238], Cout[239], S[921], Cout[921]);
	Full_Adder FA885 (Cout[240], Cout[241], Cout[242], S[922], Cout[922]);
	Full_Adder FA886 (Cout[243], Cout[244], Cout[245], S[923], Cout[923]);
	Full_Adder FA887 (Cout[246], Cout[247], Cout[248], S[924], Cout[924]);
	Full_Adder FA888 (Cout[249], Cout[250], Cout[251], S[925], Cout[925]);
	Full_Adder FA889 (Cout[252], Cout[253], Cout[254], S[926], Cout[926]);
	Full_Adder FA890 (S[255], S[256], S[257], S[927], Cout[927]);
	Full_Adder FA891 (S[258], S[259], S[260], S[928], Cout[928]);
	Full_Adder FA892 (S[261], S[262], S[263], S[929], Cout[929]);
	Full_Adder FA893 (S[264], S[265], S[266], S[930], Cout[930]);
	Full_Adder FA894 (S[267], S[268], S[269], S[931], Cout[931]);
	Full_Adder FA895 (S[270], S[271], S[272], S[932], Cout[932]);
	Full_Adder FA896 (S[273], S[274], S[275], S[933], Cout[933]);
	Full_Adder FA897 (Cout[255], Cout[256], Cout[257], S[934], Cout[934]);
	Full_Adder FA898 (Cout[258], Cout[259], Cout[260], S[935], Cout[935]);
	Full_Adder FA899 (Cout[261], Cout[262], Cout[263], S[936], Cout[936]);
	Full_Adder FA900 (Cout[264], Cout[265], Cout[266], S[937], Cout[937]);
	Full_Adder FA901 (Cout[267], Cout[268], Cout[269], S[938], Cout[938]);
	Full_Adder FA902 (Cout[270], Cout[271], Cout[272], S[939], Cout[939]);
	Full_Adder FA903 (Cout[273], Cout[274], Cout[275], S[940], Cout[940]);
	Full_Adder FA904 (S[276], S[277], S[278], S[941], Cout[941]);
	Full_Adder FA905 (S[279], S[280], S[281], S[942], Cout[942]);
	Full_Adder FA906 (S[282], S[283], S[284], S[943], Cout[943]);
	Full_Adder FA907 (S[285], S[286], S[287], S[944], Cout[944]);
	Full_Adder FA908 (S[288], S[289], S[290], S[945], Cout[945]);
	Full_Adder FA909 (S[291], S[292], S[293], S[946], Cout[946]);
	Full_Adder FA910 (S[294], S[295], S[296], S[947], Cout[947]);
	Full_Adder FA911 (pp63[3], Cout[276], Cout[277], S[948], Cout[948]);
	Full_Adder FA912 (Cout[278], Cout[279], Cout[280], S[949], Cout[949]);
	Full_Adder FA913 (Cout[281], Cout[282], Cout[283], S[950], Cout[950]);
	Full_Adder FA914 (Cout[284], Cout[285], Cout[286], S[951], Cout[951]);
	Full_Adder FA915 (Cout[287], Cout[288], Cout[289], S[952], Cout[952]);
	Full_Adder FA916 (Cout[290], Cout[291], Cout[292], S[953], Cout[953]);
	Full_Adder FA917 (Cout[293], Cout[294], Cout[295], S[954], Cout[954]);
	Full_Adder FA918 (Cout[296], S[297], S[298], S[955], Cout[955]);
	Full_Adder FA919 (S[299], S[300], S[301], S[956], Cout[956]);
	Full_Adder FA920 (S[302], S[303], S[304], S[957], Cout[957]);
	Full_Adder FA921 (S[305], S[306], S[307], S[958], Cout[958]);
	Full_Adder FA922 (S[308], S[309], S[310], S[959], Cout[959]);
	Full_Adder FA923 (S[311], S[312], S[313], S[960], Cout[960]);
	Full_Adder FA924 (S[314], S[315], S[316], S[961], Cout[961]);
	Full_Adder FA925 (pp61[6], pp62[5], pp63[4], S[962], Cout[962]);
	Full_Adder FA926 (Cout[297], Cout[298], Cout[299], S[963], Cout[963]);
	Full_Adder FA927 (Cout[300], Cout[301], Cout[302], S[964], Cout[964]);
	Full_Adder FA928 (Cout[303], Cout[304], Cout[305], S[965], Cout[965]);
	Full_Adder FA929 (Cout[306], Cout[307], Cout[308], S[966], Cout[966]);
	Full_Adder FA930 (Cout[309], Cout[310], Cout[311], S[967], Cout[967]);
	Full_Adder FA931 (Cout[312], Cout[313], Cout[314], S[968], Cout[968]);
	Full_Adder FA932 (Cout[315], Cout[316], S[317], S[969], Cout[969]);
	Full_Adder FA933 (S[318], S[319], S[320], S[970], Cout[970]);
	Full_Adder FA934 (S[321], S[322], S[323], S[971], Cout[971]);
	Full_Adder FA935 (S[324], S[325], S[326], S[972], Cout[972]);
	Full_Adder FA936 (S[327], S[328], S[329], S[973], Cout[973]);
	Full_Adder FA937 (S[330], S[331], S[332], S[974], Cout[974]);
	Full_Adder FA938 (S[333], S[334], S[335], S[975], Cout[975]);
	Full_Adder FA939 (pp59[9], pp60[8], pp61[7], S[976], Cout[976]);
	Full_Adder FA940 (pp62[6], pp63[5], Cout[317], S[977], Cout[977]);
	Full_Adder FA941 (Cout[318], Cout[319], Cout[320], S[978], Cout[978]);
	Full_Adder FA942 (Cout[321], Cout[322], Cout[323], S[979], Cout[979]);
	Full_Adder FA943 (Cout[324], Cout[325], Cout[326], S[980], Cout[980]);
	Full_Adder FA944 (Cout[327], Cout[328], Cout[329], S[981], Cout[981]);
	Full_Adder FA945 (Cout[330], Cout[331], Cout[332], S[982], Cout[982]);
	Full_Adder FA946 (Cout[333], Cout[334], Cout[335], S[983], Cout[983]);
	Full_Adder FA947 (S[336], S[337], S[338], S[984], Cout[984]);
	Full_Adder FA948 (S[339], S[340], S[341], S[985], Cout[985]);
	Full_Adder FA949 (S[342], S[343], S[344], S[986], Cout[986]);
	Full_Adder FA950 (S[345], S[346], S[347], S[987], Cout[987]);
	Full_Adder FA951 (S[348], S[349], S[350], S[988], Cout[988]);
	Full_Adder FA952 (S[351], S[352], S[353], S[989], Cout[989]);
	Full_Adder FA953 (pp57[12], pp58[11], pp59[10], S[990], Cout[990]);
	Full_Adder FA954 (pp60[9], pp61[8], pp62[7], S[991], Cout[991]);
	Full_Adder FA955 (pp63[6], Cout[336], Cout[337], S[992], Cout[992]);
	Full_Adder FA956 (Cout[338], Cout[339], Cout[340], S[993], Cout[993]);
	Full_Adder FA957 (Cout[341], Cout[342], Cout[343], S[994], Cout[994]);
	Full_Adder FA958 (Cout[344], Cout[345], Cout[346], S[995], Cout[995]);
	Full_Adder FA959 (Cout[347], Cout[348], Cout[349], S[996], Cout[996]);
	Full_Adder FA960 (Cout[350], Cout[351], Cout[352], S[997], Cout[997]);
	Full_Adder FA961 (Cout[353], S[354], S[355], S[998], Cout[998]);
	Full_Adder FA962 (S[356], S[357], S[358], S[999], Cout[999]);
	Full_Adder FA963 (S[359], S[360], S[361], S[1000], Cout[1000]);
	Full_Adder FA964 (S[362], S[363], S[364], S[1001], Cout[1001]);
	Full_Adder FA965 (S[365], S[366], S[367], S[1002], Cout[1002]);
	Full_Adder FA966 (S[368], S[369], S[370], S[1003], Cout[1003]);
	Full_Adder FA967 (pp55[15], pp56[14], pp57[13], S[1004], Cout[1004]);
	Full_Adder FA968 (pp58[12], pp59[11], pp60[10], S[1005], Cout[1005]);
	Full_Adder FA969 (pp61[9], pp62[8], pp63[7], S[1006], Cout[1006]);
	Full_Adder FA970 (Cout[354], Cout[355], Cout[356], S[1007], Cout[1007]);
	Full_Adder FA971 (Cout[357], Cout[358], Cout[359], S[1008], Cout[1008]);
	Full_Adder FA972 (Cout[360], Cout[361], Cout[362], S[1009], Cout[1009]);
	Full_Adder FA973 (Cout[363], Cout[364], Cout[365], S[1010], Cout[1010]);
	Full_Adder FA974 (Cout[366], Cout[367], Cout[368], S[1011], Cout[1011]);
	Full_Adder FA975 (Cout[369], Cout[370], S[371], S[1012], Cout[1012]);
	Full_Adder FA976 (S[372], S[373], S[374], S[1013], Cout[1013]);
	Full_Adder FA977 (S[375], S[376], S[377], S[1014], Cout[1014]);
	Full_Adder FA978 (S[378], S[379], S[380], S[1015], Cout[1015]);
	Full_Adder FA979 (S[381], S[382], S[383], S[1016], Cout[1016]);
	Full_Adder FA980 (S[384], S[385], S[386], S[1017], Cout[1017]);
	Full_Adder FA981 (pp53[18], pp54[17], pp55[16], S[1018], Cout[1018]);
	Full_Adder FA982 (pp56[15], pp57[14], pp58[13], S[1019], Cout[1019]);
	Full_Adder FA983 (pp59[12], pp60[11], pp61[10], S[1020], Cout[1020]);
	Full_Adder FA984 (pp62[9], pp63[8], Cout[371], S[1021], Cout[1021]);
	Full_Adder FA985 (Cout[372], Cout[373], Cout[374], S[1022], Cout[1022]);
	Full_Adder FA986 (Cout[375], Cout[376], Cout[377], S[1023], Cout[1023]);
	Full_Adder FA987 (Cout[378], Cout[379], Cout[380], S[1024], Cout[1024]);
	Full_Adder FA988 (Cout[381], Cout[382], Cout[383], S[1025], Cout[1025]);
	Full_Adder FA989 (Cout[384], Cout[385], Cout[386], S[1026], Cout[1026]);
	Full_Adder FA990 (S[387], S[388], S[389], S[1027], Cout[1027]);
	Full_Adder FA991 (S[390], S[391], S[392], S[1028], Cout[1028]);
	Full_Adder FA992 (S[393], S[394], S[395], S[1029], Cout[1029]);
	Full_Adder FA993 (S[396], S[397], S[398], S[1030], Cout[1030]);
	Full_Adder FA994 (S[399], S[400], S[401], S[1031], Cout[1031]);
	Full_Adder FA995 (pp51[21], pp52[20], pp53[19], S[1032], Cout[1032]);
	Full_Adder FA996 (pp54[18], pp55[17], pp56[16], S[1033], Cout[1033]);
	Full_Adder FA997 (pp57[15], pp58[14], pp59[13], S[1034], Cout[1034]);
	Full_Adder FA998 (pp60[12], pp61[11], pp62[10], S[1035], Cout[1035]);
	Full_Adder FA999 (pp63[9], Cout[387], Cout[388], S[1036], Cout[1036]);
	Full_Adder FA1000 (Cout[389], Cout[390], Cout[391], S[1037], Cout[1037]);
	Full_Adder FA1001 (Cout[392], Cout[393], Cout[394], S[1038], Cout[1038]);
	Full_Adder FA1002 (Cout[395], Cout[396], Cout[397], S[1039], Cout[1039]);
	Full_Adder FA1003 (Cout[398], Cout[399], Cout[400], S[1040], Cout[1040]);
	Full_Adder FA1004 (Cout[401], S[402], S[403], S[1041], Cout[1041]);
	Full_Adder FA1005 (S[404], S[405], S[406], S[1042], Cout[1042]);
	Full_Adder FA1006 (S[407], S[408], S[409], S[1043], Cout[1043]);
	Full_Adder FA1007 (S[410], S[411], S[412], S[1044], Cout[1044]);
	Full_Adder FA1008 (S[413], S[414], S[415], S[1045], Cout[1045]);
	Full_Adder FA1009 (pp49[24], pp50[23], pp51[22], S[1046], Cout[1046]);
	Full_Adder FA1010 (pp52[21], pp53[20], pp54[19], S[1047], Cout[1047]);
	Full_Adder FA1011 (pp55[18], pp56[17], pp57[16], S[1048], Cout[1048]);
	Full_Adder FA1012 (pp58[15], pp59[14], pp60[13], S[1049], Cout[1049]);
	Full_Adder FA1013 (pp61[12], pp62[11], pp63[10], S[1050], Cout[1050]);
	Full_Adder FA1014 (Cout[402], Cout[403], Cout[404], S[1051], Cout[1051]);
	Full_Adder FA1015 (Cout[405], Cout[406], Cout[407], S[1052], Cout[1052]);
	Full_Adder FA1016 (Cout[408], Cout[409], Cout[410], S[1053], Cout[1053]);
	Full_Adder FA1017 (Cout[411], Cout[412], Cout[413], S[1054], Cout[1054]);
	Full_Adder FA1018 (Cout[414], Cout[415], S[416], S[1055], Cout[1055]);
	Full_Adder FA1019 (S[417], S[418], S[419], S[1056], Cout[1056]);
	Full_Adder FA1020 (S[420], S[421], S[422], S[1057], Cout[1057]);
	Full_Adder FA1021 (S[423], S[424], S[425], S[1058], Cout[1058]);
	Full_Adder FA1022 (S[426], S[427], S[428], S[1059], Cout[1059]);
	Full_Adder FA1023 (pp47[27], pp48[26], pp49[25], S[1060], Cout[1060]);
	Full_Adder FA1024 (pp50[24], pp51[23], pp52[22], S[1061], Cout[1061]);
	Full_Adder FA1025 (pp53[21], pp54[20], pp55[19], S[1062], Cout[1062]);
	Full_Adder FA1026 (pp56[18], pp57[17], pp58[16], S[1063], Cout[1063]);
	Full_Adder FA1027 (pp59[15], pp60[14], pp61[13], S[1064], Cout[1064]);
	Full_Adder FA1028 (pp62[12], pp63[11], Cout[416], S[1065], Cout[1065]);
	Full_Adder FA1029 (Cout[417], Cout[418], Cout[419], S[1066], Cout[1066]);
	Full_Adder FA1030 (Cout[420], Cout[421], Cout[422], S[1067], Cout[1067]);
	Full_Adder FA1031 (Cout[423], Cout[424], Cout[425], S[1068], Cout[1068]);
	Full_Adder FA1032 (Cout[426], Cout[427], Cout[428], S[1069], Cout[1069]);
	Full_Adder FA1033 (S[429], S[430], S[431], S[1070], Cout[1070]);
	Full_Adder FA1034 (S[432], S[433], S[434], S[1071], Cout[1071]);
	Full_Adder FA1035 (S[435], S[436], S[437], S[1072], Cout[1072]);
	Full_Adder FA1036 (S[438], S[439], S[440], S[1073], Cout[1073]);
	Full_Adder FA1037 (pp45[30], pp46[29], pp47[28], S[1074], Cout[1074]);
	Full_Adder FA1038 (pp48[27], pp49[26], pp50[25], S[1075], Cout[1075]);
	Full_Adder FA1039 (pp51[24], pp52[23], pp53[22], S[1076], Cout[1076]);
	Full_Adder FA1040 (pp54[21], pp55[20], pp56[19], S[1077], Cout[1077]);
	Full_Adder FA1041 (pp57[18], pp58[17], pp59[16], S[1078], Cout[1078]);
	Full_Adder FA1042 (pp60[15], pp61[14], pp62[13], S[1079], Cout[1079]);
	Full_Adder FA1043 (pp63[12], Cout[429], Cout[430], S[1080], Cout[1080]);
	Full_Adder FA1044 (Cout[431], Cout[432], Cout[433], S[1081], Cout[1081]);
	Full_Adder FA1045 (Cout[434], Cout[435], Cout[436], S[1082], Cout[1082]);
	Full_Adder FA1046 (Cout[437], Cout[438], Cout[439], S[1083], Cout[1083]);
	Full_Adder FA1047 (Cout[440], S[441], S[442], S[1084], Cout[1084]);
	Full_Adder FA1048 (S[443], S[444], S[445], S[1085], Cout[1085]);
	Full_Adder FA1049 (S[446], S[447], S[448], S[1086], Cout[1086]);
	Full_Adder FA1050 (S[449], S[450], S[451], S[1087], Cout[1087]);
	Full_Adder FA1051 (pp43[33], pp44[32], pp45[31], S[1088], Cout[1088]);
	Full_Adder FA1052 (pp46[30], pp47[29], pp48[28], S[1089], Cout[1089]);
	Full_Adder FA1053 (pp49[27], pp50[26], pp51[25], S[1090], Cout[1090]);
	Full_Adder FA1054 (pp52[24], pp53[23], pp54[22], S[1091], Cout[1091]);
	Full_Adder FA1055 (pp55[21], pp56[20], pp57[19], S[1092], Cout[1092]);
	Full_Adder FA1056 (pp58[18], pp59[17], pp60[16], S[1093], Cout[1093]);
	Full_Adder FA1057 (pp61[15], pp62[14], pp63[13], S[1094], Cout[1094]);
	Full_Adder FA1058 (Cout[441], Cout[442], Cout[443], S[1095], Cout[1095]);
	Full_Adder FA1059 (Cout[444], Cout[445], Cout[446], S[1096], Cout[1096]);
	Full_Adder FA1060 (Cout[447], Cout[448], Cout[449], S[1097], Cout[1097]);
	Full_Adder FA1061 (Cout[450], Cout[451], S[452], S[1098], Cout[1098]);
	Full_Adder FA1062 (S[453], S[454], S[455], S[1099], Cout[1099]);
	Full_Adder FA1063 (S[456], S[457], S[458], S[1100], Cout[1100]);
	Full_Adder FA1064 (S[459], S[460], S[461], S[1101], Cout[1101]);
	Full_Adder FA1065 (pp41[36], pp42[35], pp43[34], S[1102], Cout[1102]);
	Full_Adder FA1066 (pp44[33], pp45[32], pp46[31], S[1103], Cout[1103]);
	Full_Adder FA1067 (pp47[30], pp48[29], pp49[28], S[1104], Cout[1104]);
	Full_Adder FA1068 (pp50[27], pp51[26], pp52[25], S[1105], Cout[1105]);
	Full_Adder FA1069 (pp53[24], pp54[23], pp55[22], S[1106], Cout[1106]);
	Full_Adder FA1070 (pp56[21], pp57[20], pp58[19], S[1107], Cout[1107]);
	Full_Adder FA1071 (pp59[18], pp60[17], pp61[16], S[1108], Cout[1108]);
	Full_Adder FA1072 (pp62[15], pp63[14], Cout[452], S[1109], Cout[1109]);
	Full_Adder FA1073 (Cout[453], Cout[454], Cout[455], S[1110], Cout[1110]);
	Full_Adder FA1074 (Cout[456], Cout[457], Cout[458], S[1111], Cout[1111]);
	Full_Adder FA1075 (Cout[459], Cout[460], Cout[461], S[1112], Cout[1112]);
	Full_Adder FA1076 (S[462], S[463], S[464], S[1113], Cout[1113]);
	Full_Adder FA1077 (S[465], S[466], S[467], S[1114], Cout[1114]);
	Full_Adder FA1078 (S[468], S[469], S[470], S[1115], Cout[1115]);
	Full_Adder FA1079 (pp39[39], pp40[38], pp41[37], S[1116], Cout[1116]);
	Full_Adder FA1080 (pp42[36], pp43[35], pp44[34], S[1117], Cout[1117]);
	Full_Adder FA1081 (pp45[33], pp46[32], pp47[31], S[1118], Cout[1118]);
	Full_Adder FA1082 (pp48[30], pp49[29], pp50[28], S[1119], Cout[1119]);
	Full_Adder FA1083 (pp51[27], pp52[26], pp53[25], S[1120], Cout[1120]);
	Full_Adder FA1084 (pp54[24], pp55[23], pp56[22], S[1121], Cout[1121]);
	Full_Adder FA1085 (pp57[21], pp58[20], pp59[19], S[1122], Cout[1122]);
	Full_Adder FA1086 (pp60[18], pp61[17], pp62[16], S[1123], Cout[1123]);
	Full_Adder FA1087 (pp63[15], Cout[462], Cout[463], S[1124], Cout[1124]);
	Full_Adder FA1088 (Cout[464], Cout[465], Cout[466], S[1125], Cout[1125]);
	Full_Adder FA1089 (Cout[467], Cout[468], Cout[469], S[1126], Cout[1126]);
	Full_Adder FA1090 (Cout[470], S[471], S[472], S[1127], Cout[1127]);
	Full_Adder FA1091 (S[473], S[474], S[475], S[1128], Cout[1128]);
	Full_Adder FA1092 (S[476], S[477], S[478], S[1129], Cout[1129]);
	Full_Adder FA1093 (pp37[42], pp38[41], pp39[40], S[1130], Cout[1130]);
	Full_Adder FA1094 (pp40[39], pp41[38], pp42[37], S[1131], Cout[1131]);
	Full_Adder FA1095 (pp43[36], pp44[35], pp45[34], S[1132], Cout[1132]);
	Full_Adder FA1096 (pp46[33], pp47[32], pp48[31], S[1133], Cout[1133]);
	Full_Adder FA1097 (pp49[30], pp50[29], pp51[28], S[1134], Cout[1134]);
	Full_Adder FA1098 (pp52[27], pp53[26], pp54[25], S[1135], Cout[1135]);
	Full_Adder FA1099 (pp55[24], pp56[23], pp57[22], S[1136], Cout[1136]);
	Full_Adder FA1100 (pp58[21], pp59[20], pp60[19], S[1137], Cout[1137]);
	Full_Adder FA1101 (pp61[18], pp62[17], pp63[16], S[1138], Cout[1138]);
	Full_Adder FA1102 (Cout[471], Cout[472], Cout[473], S[1139], Cout[1139]);
	Full_Adder FA1103 (Cout[474], Cout[475], Cout[476], S[1140], Cout[1140]);
	Full_Adder FA1104 (Cout[477], Cout[478], S[479], S[1141], Cout[1141]);
	Full_Adder FA1105 (S[480], S[481], S[482], S[1142], Cout[1142]);
	Full_Adder FA1106 (S[483], S[484], S[485], S[1143], Cout[1143]);
	Full_Adder FA1107 (pp35[45], pp36[44], pp37[43], S[1144], Cout[1144]);
	Full_Adder FA1108 (pp38[42], pp39[41], pp40[40], S[1145], Cout[1145]);
	Full_Adder FA1109 (pp41[39], pp42[38], pp43[37], S[1146], Cout[1146]);
	Full_Adder FA1110 (pp44[36], pp45[35], pp46[34], S[1147], Cout[1147]);
	Full_Adder FA1111 (pp47[33], pp48[32], pp49[31], S[1148], Cout[1148]);
	Full_Adder FA1112 (pp50[30], pp51[29], pp52[28], S[1149], Cout[1149]);
	Full_Adder FA1113 (pp53[27], pp54[26], pp55[25], S[1150], Cout[1150]);
	Full_Adder FA1114 (pp56[24], pp57[23], pp58[22], S[1151], Cout[1151]);
	Full_Adder FA1115 (pp59[21], pp60[20], pp61[19], S[1152], Cout[1152]);
	Full_Adder FA1116 (pp62[18], pp63[17], Cout[479], S[1153], Cout[1153]);
	Full_Adder FA1117 (Cout[480], Cout[481], Cout[482], S[1154], Cout[1154]);
	Full_Adder FA1118 (Cout[483], Cout[484], Cout[485], S[1155], Cout[1155]);
	Full_Adder FA1119 (S[486], S[487], S[488], S[1156], Cout[1156]);
	Full_Adder FA1120 (S[489], S[490], S[491], S[1157], Cout[1157]);
	Full_Adder FA1121 (pp33[48], pp34[47], pp35[46], S[1158], Cout[1158]);
	Full_Adder FA1122 (pp36[45], pp37[44], pp38[43], S[1159], Cout[1159]);
	Full_Adder FA1123 (pp39[42], pp40[41], pp41[40], S[1160], Cout[1160]);
	Full_Adder FA1124 (pp42[39], pp43[38], pp44[37], S[1161], Cout[1161]);
	Full_Adder FA1125 (pp45[36], pp46[35], pp47[34], S[1162], Cout[1162]);
	Full_Adder FA1126 (pp48[33], pp49[32], pp50[31], S[1163], Cout[1163]);
	Full_Adder FA1127 (pp51[30], pp52[29], pp53[28], S[1164], Cout[1164]);
	Full_Adder FA1128 (pp54[27], pp55[26], pp56[25], S[1165], Cout[1165]);
	Full_Adder FA1129 (pp57[24], pp58[23], pp59[22], S[1166], Cout[1166]);
	Full_Adder FA1130 (pp60[21], pp61[20], pp62[19], S[1167], Cout[1167]);
	Full_Adder FA1131 (pp63[18], Cout[486], Cout[487], S[1168], Cout[1168]);
	Full_Adder FA1132 (Cout[488], Cout[489], Cout[490], S[1169], Cout[1169]);
	Full_Adder FA1133 (Cout[491], S[492], S[493], S[1170], Cout[1170]);
	Full_Adder FA1134 (S[494], S[495], S[496], S[1171], Cout[1171]);
	Full_Adder FA1135 (pp31[51], pp32[50], pp33[49], S[1172], Cout[1172]);
	Full_Adder FA1136 (pp34[48], pp35[47], pp36[46], S[1173], Cout[1173]);
	Full_Adder FA1137 (pp37[45], pp38[44], pp39[43], S[1174], Cout[1174]);
	Full_Adder FA1138 (pp40[42], pp41[41], pp42[40], S[1175], Cout[1175]);
	Full_Adder FA1139 (pp43[39], pp44[38], pp45[37], S[1176], Cout[1176]);
	Full_Adder FA1140 (pp46[36], pp47[35], pp48[34], S[1177], Cout[1177]);
	Full_Adder FA1141 (pp49[33], pp50[32], pp51[31], S[1178], Cout[1178]);
	Full_Adder FA1142 (pp52[30], pp53[29], pp54[28], S[1179], Cout[1179]);
	Full_Adder FA1143 (pp55[27], pp56[26], pp57[25], S[1180], Cout[1180]);
	Full_Adder FA1144 (pp58[24], pp59[23], pp60[22], S[1181], Cout[1181]);
	Full_Adder FA1145 (pp61[21], pp62[20], pp63[19], S[1182], Cout[1182]);
	Full_Adder FA1146 (Cout[492], Cout[493], Cout[494], S[1183], Cout[1183]);
	Full_Adder FA1147 (Cout[495], Cout[496], S[497], S[1184], Cout[1184]);
	Full_Adder FA1148 (S[498], S[499], S[500], S[1185], Cout[1185]);
	Full_Adder FA1149 (pp29[54], pp30[53], pp31[52], S[1186], Cout[1186]);
	Full_Adder FA1150 (pp32[51], pp33[50], pp34[49], S[1187], Cout[1187]);
	Full_Adder FA1151 (pp35[48], pp36[47], pp37[46], S[1188], Cout[1188]);
	Full_Adder FA1152 (pp38[45], pp39[44], pp40[43], S[1189], Cout[1189]);
	Full_Adder FA1153 (pp41[42], pp42[41], pp43[40], S[1190], Cout[1190]);
	Full_Adder FA1154 (pp44[39], pp45[38], pp46[37], S[1191], Cout[1191]);
	Full_Adder FA1155 (pp47[36], pp48[35], pp49[34], S[1192], Cout[1192]);
	Full_Adder FA1156 (pp50[33], pp51[32], pp52[31], S[1193], Cout[1193]);
	Full_Adder FA1157 (pp53[30], pp54[29], pp55[28], S[1194], Cout[1194]);
	Full_Adder FA1158 (pp56[27], pp57[26], pp58[25], S[1195], Cout[1195]);
	Full_Adder FA1159 (pp59[24], pp60[23], pp61[22], S[1196], Cout[1196]);
	Full_Adder FA1160 (pp62[21], pp63[20], Cout[497], S[1197], Cout[1197]);
	Full_Adder FA1161 (Cout[498], Cout[499], Cout[500], S[1198], Cout[1198]);
	Full_Adder FA1162 (S[501], S[502], S[503], S[1199], Cout[1199]);
	Full_Adder FA1163 (pp27[57], pp28[56], pp29[55], S[1200], Cout[1200]);
	Full_Adder FA1164 (pp30[54], pp31[53], pp32[52], S[1201], Cout[1201]);
	Full_Adder FA1165 (pp33[51], pp34[50], pp35[49], S[1202], Cout[1202]);
	Full_Adder FA1166 (pp36[48], pp37[47], pp38[46], S[1203], Cout[1203]);
	Full_Adder FA1167 (pp39[45], pp40[44], pp41[43], S[1204], Cout[1204]);
	Full_Adder FA1168 (pp42[42], pp43[41], pp44[40], S[1205], Cout[1205]);
	Full_Adder FA1169 (pp45[39], pp46[38], pp47[37], S[1206], Cout[1206]);
	Full_Adder FA1170 (pp48[36], pp49[35], pp50[34], S[1207], Cout[1207]);
	Full_Adder FA1171 (pp51[33], pp52[32], pp53[31], S[1208], Cout[1208]);
	Full_Adder FA1172 (pp54[30], pp55[29], pp56[28], S[1209], Cout[1209]);
	Full_Adder FA1173 (pp57[27], pp58[26], pp59[25], S[1210], Cout[1210]);
	Full_Adder FA1174 (pp60[24], pp61[23], pp62[22], S[1211], Cout[1211]);
	Full_Adder FA1175 (pp63[21], Cout[501], Cout[502], S[1212], Cout[1212]);
	Full_Adder FA1176 (Cout[503], S[504], S[505], S[1213], Cout[1213]);
	Full_Adder FA1177 (pp25[60], pp26[59], pp27[58], S[1214], Cout[1214]);
	Full_Adder FA1178 (pp28[57], pp29[56], pp30[55], S[1215], Cout[1215]);
	Full_Adder FA1179 (pp31[54], pp32[53], pp33[52], S[1216], Cout[1216]);
	Full_Adder FA1180 (pp34[51], pp35[50], pp36[49], S[1217], Cout[1217]);
	Full_Adder FA1181 (pp37[48], pp38[47], pp39[46], S[1218], Cout[1218]);
	Full_Adder FA1182 (pp40[45], pp41[44], pp42[43], S[1219], Cout[1219]);
	Full_Adder FA1183 (pp43[42], pp44[41], pp45[40], S[1220], Cout[1220]);
	Full_Adder FA1184 (pp46[39], pp47[38], pp48[37], S[1221], Cout[1221]);
	Full_Adder FA1185 (pp49[36], pp50[35], pp51[34], S[1222], Cout[1222]);
	Full_Adder FA1186 (pp52[33], pp53[32], pp54[31], S[1223], Cout[1223]);
	Full_Adder FA1187 (pp55[30], pp56[29], pp57[28], S[1224], Cout[1224]);
	Full_Adder FA1188 (pp58[27], pp59[26], pp60[25], S[1225], Cout[1225]);
	Full_Adder FA1189 (pp61[24], pp62[23], pp63[22], S[1226], Cout[1226]);
	Full_Adder FA1190 (Cout[504], Cout[505], S[506], S[1227], Cout[1227]);
	Full_Adder FA1191 (pp23[63], pp24[62], pp25[61], S[1228], Cout[1228]);
	Full_Adder FA1192 (pp26[60], pp27[59], pp28[58], S[1229], Cout[1229]);
	Full_Adder FA1193 (pp29[57], pp30[56], pp31[55], S[1230], Cout[1230]);
	Full_Adder FA1194 (pp32[54], pp33[53], pp34[52], S[1231], Cout[1231]);
	Full_Adder FA1195 (pp35[51], pp36[50], pp37[49], S[1232], Cout[1232]);
	Full_Adder FA1196 (pp38[48], pp39[47], pp40[46], S[1233], Cout[1233]);
	Full_Adder FA1197 (pp41[45], pp42[44], pp43[43], S[1234], Cout[1234]);
	Full_Adder FA1198 (pp44[42], pp45[41], pp46[40], S[1235], Cout[1235]);
	Full_Adder FA1199 (pp47[39], pp48[38], pp49[37], S[1236], Cout[1236]);
	Full_Adder FA1200 (pp50[36], pp51[35], pp52[34], S[1237], Cout[1237]);
	Full_Adder FA1201 (pp53[33], pp54[32], pp55[31], S[1238], Cout[1238]);
	Full_Adder FA1202 (pp56[30], pp57[29], pp58[28], S[1239], Cout[1239]);
	Full_Adder FA1203 (pp59[27], pp60[26], pp61[25], S[1240], Cout[1240]);
	Full_Adder FA1204 (pp62[24], pp63[23], Cout[506], S[1241], Cout[1241]);
	Full_Adder FA1205 (pp24[63], pp25[62], pp26[61], S[1242], Cout[1242]);
	Full_Adder FA1206 (pp27[60], pp28[59], pp29[58], S[1243], Cout[1243]);
	Full_Adder FA1207 (pp30[57], pp31[56], pp32[55], S[1244], Cout[1244]);
	Full_Adder FA1208 (pp33[54], pp34[53], pp35[52], S[1245], Cout[1245]);
	Full_Adder FA1209 (pp36[51], pp37[50], pp38[49], S[1246], Cout[1246]);
	Full_Adder FA1210 (pp39[48], pp40[47], pp41[46], S[1247], Cout[1247]);
	Full_Adder FA1211 (pp42[45], pp43[44], pp44[43], S[1248], Cout[1248]);
	Full_Adder FA1212 (pp45[42], pp46[41], pp47[40], S[1249], Cout[1249]);
	Full_Adder FA1213 (pp48[39], pp49[38], pp50[37], S[1250], Cout[1250]);
	Full_Adder FA1214 (pp51[36], pp52[35], pp53[34], S[1251], Cout[1251]);
	Full_Adder FA1215 (pp54[33], pp55[32], pp56[31], S[1252], Cout[1252]);
	Full_Adder FA1216 (pp57[30], pp58[29], pp59[28], S[1253], Cout[1253]);
	Full_Adder FA1217 (pp60[27], pp61[26], pp62[25], S[1254], Cout[1254]);
	Full_Adder FA1218 (pp25[63], pp26[62], pp27[61], S[1255], Cout[1255]);
	Full_Adder FA1219 (pp28[60], pp29[59], pp30[58], S[1256], Cout[1256]);
	Full_Adder FA1220 (pp31[57], pp32[56], pp33[55], S[1257], Cout[1257]);
	Full_Adder FA1221 (pp34[54], pp35[53], pp36[52], S[1258], Cout[1258]);
	Full_Adder FA1222 (pp37[51], pp38[50], pp39[49], S[1259], Cout[1259]);
	Full_Adder FA1223 (pp40[48], pp41[47], pp42[46], S[1260], Cout[1260]);
	Full_Adder FA1224 (pp43[45], pp44[44], pp45[43], S[1261], Cout[1261]);
	Full_Adder FA1225 (pp46[42], pp47[41], pp48[40], S[1262], Cout[1262]);
	Full_Adder FA1226 (pp49[39], pp50[38], pp51[37], S[1263], Cout[1263]);
	Full_Adder FA1227 (pp52[36], pp53[35], pp54[34], S[1264], Cout[1264]);
	Full_Adder FA1228 (pp55[33], pp56[32], pp57[31], S[1265], Cout[1265]);
	Full_Adder FA1229 (pp58[30], pp59[29], pp60[28], S[1266], Cout[1266]);
	Full_Adder FA1230 (pp26[63], pp27[62], pp28[61], S[1267], Cout[1267]);
	Full_Adder FA1231 (pp29[60], pp30[59], pp31[58], S[1268], Cout[1268]);
	Full_Adder FA1232 (pp32[57], pp33[56], pp34[55], S[1269], Cout[1269]);
	Full_Adder FA1233 (pp35[54], pp36[53], pp37[52], S[1270], Cout[1270]);
	Full_Adder FA1234 (pp38[51], pp39[50], pp40[49], S[1271], Cout[1271]);
	Full_Adder FA1235 (pp41[48], pp42[47], pp43[46], S[1272], Cout[1272]);
	Full_Adder FA1236 (pp44[45], pp45[44], pp46[43], S[1273], Cout[1273]);
	Full_Adder FA1237 (pp47[42], pp48[41], pp49[40], S[1274], Cout[1274]);
	Full_Adder FA1238 (pp50[39], pp51[38], pp52[37], S[1275], Cout[1275]);
	Full_Adder FA1239 (pp53[36], pp54[35], pp55[34], S[1276], Cout[1276]);
	Full_Adder FA1240 (pp56[33], pp57[32], pp58[31], S[1277], Cout[1277]);
	Full_Adder FA1241 (pp27[63], pp28[62], pp29[61], S[1278], Cout[1278]);
	Full_Adder FA1242 (pp30[60], pp31[59], pp32[58], S[1279], Cout[1279]);
	Full_Adder FA1243 (pp33[57], pp34[56], pp35[55], S[1280], Cout[1280]);
	Full_Adder FA1244 (pp36[54], pp37[53], pp38[52], S[1281], Cout[1281]);
	Full_Adder FA1245 (pp39[51], pp40[50], pp41[49], S[1282], Cout[1282]);
	Full_Adder FA1246 (pp42[48], pp43[47], pp44[46], S[1283], Cout[1283]);
	Full_Adder FA1247 (pp45[45], pp46[44], pp47[43], S[1284], Cout[1284]);
	Full_Adder FA1248 (pp48[42], pp49[41], pp50[40], S[1285], Cout[1285]);
	Full_Adder FA1249 (pp51[39], pp52[38], pp53[37], S[1286], Cout[1286]);
	Full_Adder FA1250 (pp54[36], pp55[35], pp56[34], S[1287], Cout[1287]);
	Full_Adder FA1251 (pp28[63], pp29[62], pp30[61], S[1288], Cout[1288]);
	Full_Adder FA1252 (pp31[60], pp32[59], pp33[58], S[1289], Cout[1289]);
	Full_Adder FA1253 (pp34[57], pp35[56], pp36[55], S[1290], Cout[1290]);
	Full_Adder FA1254 (pp37[54], pp38[53], pp39[52], S[1291], Cout[1291]);
	Full_Adder FA1255 (pp40[51], pp41[50], pp42[49], S[1292], Cout[1292]);
	Full_Adder FA1256 (pp43[48], pp44[47], pp45[46], S[1293], Cout[1293]);
	Full_Adder FA1257 (pp46[45], pp47[44], pp48[43], S[1294], Cout[1294]);
	Full_Adder FA1258 (pp49[42], pp50[41], pp51[40], S[1295], Cout[1295]);
	Full_Adder FA1259 (pp52[39], pp53[38], pp54[37], S[1296], Cout[1296]);
	Full_Adder FA1260 (pp29[63], pp30[62], pp31[61], S[1297], Cout[1297]);
	Full_Adder FA1261 (pp32[60], pp33[59], pp34[58], S[1298], Cout[1298]);
	Full_Adder FA1262 (pp35[57], pp36[56], pp37[55], S[1299], Cout[1299]);
	Full_Adder FA1263 (pp38[54], pp39[53], pp40[52], S[1300], Cout[1300]);
	Full_Adder FA1264 (pp41[51], pp42[50], pp43[49], S[1301], Cout[1301]);
	Full_Adder FA1265 (pp44[48], pp45[47], pp46[46], S[1302], Cout[1302]);
	Full_Adder FA1266 (pp47[45], pp48[44], pp49[43], S[1303], Cout[1303]);
	Full_Adder FA1267 (pp50[42], pp51[41], pp52[40], S[1304], Cout[1304]);
	Full_Adder FA1268 (pp30[63], pp31[62], pp32[61], S[1305], Cout[1305]);
	Full_Adder FA1269 (pp33[60], pp34[59], pp35[58], S[1306], Cout[1306]);
	Full_Adder FA1270 (pp36[57], pp37[56], pp38[55], S[1307], Cout[1307]);
	Full_Adder FA1271 (pp39[54], pp40[53], pp41[52], S[1308], Cout[1308]);
	Full_Adder FA1272 (pp42[51], pp43[50], pp44[49], S[1309], Cout[1309]);
	Full_Adder FA1273 (pp45[48], pp46[47], pp47[46], S[1310], Cout[1310]);
	Full_Adder FA1274 (pp48[45], pp49[44], pp50[43], S[1311], Cout[1311]);
	Full_Adder FA1275 (pp31[63], pp32[62], pp33[61], S[1312], Cout[1312]);
	Full_Adder FA1276 (pp34[60], pp35[59], pp36[58], S[1313], Cout[1313]);
	Full_Adder FA1277 (pp37[57], pp38[56], pp39[55], S[1314], Cout[1314]);
	Full_Adder FA1278 (pp40[54], pp41[53], pp42[52], S[1315], Cout[1315]);
	Full_Adder FA1279 (pp43[51], pp44[50], pp45[49], S[1316], Cout[1316]);
	Full_Adder FA1280 (pp46[48], pp47[47], pp48[46], S[1317], Cout[1317]);
	Full_Adder FA1281 (pp32[63], pp33[62], pp34[61], S[1318], Cout[1318]);
	Full_Adder FA1282 (pp35[60], pp36[59], pp37[58], S[1319], Cout[1319]);
	Full_Adder FA1283 (pp38[57], pp39[56], pp40[55], S[1320], Cout[1320]);
	Full_Adder FA1284 (pp41[54], pp42[53], pp43[52], S[1321], Cout[1321]);
	Full_Adder FA1285 (pp44[51], pp45[50], pp46[49], S[1322], Cout[1322]);
	Full_Adder FA1286 (pp33[63], pp34[62], pp35[61], S[1323], Cout[1323]);
	Full_Adder FA1287 (pp36[60], pp37[59], pp38[58], S[1324], Cout[1324]);
	Full_Adder FA1288 (pp39[57], pp40[56], pp41[55], S[1325], Cout[1325]);
	Full_Adder FA1289 (pp42[54], pp43[53], pp44[52], S[1326], Cout[1326]);
	Full_Adder FA1290 (pp34[63], pp35[62], pp36[61], S[1327], Cout[1327]);
	Full_Adder FA1291 (pp37[60], pp38[59], pp39[58], S[1328], Cout[1328]);
	Full_Adder FA1292 (pp40[57], pp41[56], pp42[55], S[1329], Cout[1329]);
	Full_Adder FA1293 (pp35[63], pp36[62], pp37[61], S[1330], Cout[1330]);
	Full_Adder FA1294 (pp38[60], pp39[59], pp40[58], S[1331], Cout[1331]);
	Full_Adder FA1295 (pp36[63], pp37[62], pp38[61], S[1332], Cout[1332]);
	Half_Adder HA38 (pp0[19], pp1[18], S[1333], Cout[1333]);
	Full_Adder FA1296 (pp0[20], pp1[19], pp2[18], S[1334], Cout[1334]);
	Half_Adder HA39 (pp3[17], pp4[16], S[1335], Cout[1335]);
	Full_Adder FA1297 (pp0[21], pp1[20], pp2[19], S[1336], Cout[1336]);
	Full_Adder FA1298 (pp3[18], pp4[17], pp5[16], S[1337], Cout[1337]);
	Half_Adder HA40 (pp6[15], pp7[14], S[1338], Cout[1338]);
	Full_Adder FA1299 (pp0[22], pp1[21], pp2[20], S[1339], Cout[1339]);
	Full_Adder FA1300 (pp3[19], pp4[18], pp5[17], S[1340], Cout[1340]);
	Full_Adder FA1301 (pp6[16], pp7[15], pp8[14], S[1341], Cout[1341]);
	Half_Adder HA41 (pp9[13], pp10[12], S[1342], Cout[1342]);
	Full_Adder FA1302 (pp0[23], pp1[22], pp2[21], S[1343], Cout[1343]);
	Full_Adder FA1303 (pp3[20], pp4[19], pp5[18], S[1344], Cout[1344]);
	Full_Adder FA1304 (pp6[17], pp7[16], pp8[15], S[1345], Cout[1345]);
	Full_Adder FA1305 (pp9[14], pp10[13], pp11[12], S[1346], Cout[1346]);
	Half_Adder HA42 (pp12[11], pp13[10], S[1347], Cout[1347]);
	Full_Adder FA1306 (pp0[24], pp1[23], pp2[22], S[1348], Cout[1348]);
	Full_Adder FA1307 (pp3[21], pp4[20], pp5[19], S[1349], Cout[1349]);
	Full_Adder FA1308 (pp6[18], pp7[17], pp8[16], S[1350], Cout[1350]);
	Full_Adder FA1309 (pp9[15], pp10[14], pp11[13], S[1351], Cout[1351]);
	Full_Adder FA1310 (pp12[12], pp13[11], pp14[10], S[1352], Cout[1352]);
	Half_Adder HA43 (pp15[9], pp16[8], S[1353], Cout[1353]);
	Full_Adder FA1311 (pp0[25], pp1[24], pp2[23], S[1354], Cout[1354]);
	Full_Adder FA1312 (pp3[22], pp4[21], pp5[20], S[1355], Cout[1355]);
	Full_Adder FA1313 (pp6[19], pp7[18], pp8[17], S[1356], Cout[1356]);
	Full_Adder FA1314 (pp9[16], pp10[15], pp11[14], S[1357], Cout[1357]);
	Full_Adder FA1315 (pp12[13], pp13[12], pp14[11], S[1358], Cout[1358]);
	Full_Adder FA1316 (pp15[10], pp16[9], pp17[8], S[1359], Cout[1359]);
	Half_Adder HA44 (pp18[7], pp19[6], S[1360], Cout[1360]);
	Full_Adder FA1317 (pp0[26], pp1[25], pp2[24], S[1361], Cout[1361]);
	Full_Adder FA1318 (pp3[23], pp4[22], pp5[21], S[1362], Cout[1362]);
	Full_Adder FA1319 (pp6[20], pp7[19], pp8[18], S[1363], Cout[1363]);
	Full_Adder FA1320 (pp9[17], pp10[16], pp11[15], S[1364], Cout[1364]);
	Full_Adder FA1321 (pp12[14], pp13[13], pp14[12], S[1365], Cout[1365]);
	Full_Adder FA1322 (pp15[11], pp16[10], pp17[9], S[1366], Cout[1366]);
	Full_Adder FA1323 (pp18[8], pp19[7], pp20[6], S[1367], Cout[1367]);
	Half_Adder HA45 (pp21[5], pp22[4], S[1368], Cout[1368]);
	Full_Adder FA1324 (pp0[27], pp1[26], pp2[25], S[1369], Cout[1369]);
	Full_Adder FA1325 (pp3[24], pp4[23], pp5[22], S[1370], Cout[1370]);
	Full_Adder FA1326 (pp6[21], pp7[20], pp8[19], S[1371], Cout[1371]);
	Full_Adder FA1327 (pp9[18], pp10[17], pp11[16], S[1372], Cout[1372]);
	Full_Adder FA1328 (pp12[15], pp13[14], pp14[13], S[1373], Cout[1373]);
	Full_Adder FA1329 (pp15[12], pp16[11], pp17[10], S[1374], Cout[1374]);
	Full_Adder FA1330 (pp18[9], pp19[8], pp20[7], S[1375], Cout[1375]);
	Full_Adder FA1331 (pp21[6], pp22[5], pp23[4], S[1376], Cout[1376]);
	Half_Adder HA46 (pp24[3], pp25[2], S[1377], Cout[1377]);
	Full_Adder FA1332 (pp2[26], pp3[25], pp4[24], S[1378], Cout[1378]);
	Full_Adder FA1333 (pp5[23], pp6[22], pp7[21], S[1379], Cout[1379]);
	Full_Adder FA1334 (pp8[20], pp9[19], pp10[18], S[1380], Cout[1380]);
	Full_Adder FA1335 (pp11[17], pp12[16], pp13[15], S[1381], Cout[1381]);
	Full_Adder FA1336 (pp14[14], pp15[13], pp16[12], S[1382], Cout[1382]);
	Full_Adder FA1337 (pp17[11], pp18[10], pp19[9], S[1383], Cout[1383]);
	Full_Adder FA1338 (pp20[8], pp21[7], pp22[6], S[1384], Cout[1384]);
	Full_Adder FA1339 (pp23[5], pp24[4], pp25[3], S[1385], Cout[1385]);
	Full_Adder FA1340 (pp26[2], pp27[1], pp28[0], S[1386], Cout[1386]);
	Full_Adder FA1341 (pp5[24], pp6[23], pp7[22], S[1387], Cout[1387]);
	Full_Adder FA1342 (pp8[21], pp9[20], pp10[19], S[1388], Cout[1388]);
	Full_Adder FA1343 (pp11[18], pp12[17], pp13[16], S[1389], Cout[1389]);
	Full_Adder FA1344 (pp14[15], pp15[14], pp16[13], S[1390], Cout[1390]);
	Full_Adder FA1345 (pp17[12], pp18[11], pp19[10], S[1391], Cout[1391]);
	Full_Adder FA1346 (pp20[9], pp21[8], pp22[7], S[1392], Cout[1392]);
	Full_Adder FA1347 (pp23[6], pp24[5], pp25[4], S[1393], Cout[1393]);
	Full_Adder FA1348 (pp26[3], pp27[2], pp28[1], S[1394], Cout[1394]);
	Full_Adder FA1349 (pp29[0], Cout[507], S[508], S[1395], Cout[1395]);
	Full_Adder FA1350 (pp8[22], pp9[21], pp10[20], S[1396], Cout[1396]);
	Full_Adder FA1351 (pp11[19], pp12[18], pp13[17], S[1397], Cout[1397]);
	Full_Adder FA1352 (pp14[16], pp15[15], pp16[14], S[1398], Cout[1398]);
	Full_Adder FA1353 (pp17[13], pp18[12], pp19[11], S[1399], Cout[1399]);
	Full_Adder FA1354 (pp20[10], pp21[9], pp22[8], S[1400], Cout[1400]);
	Full_Adder FA1355 (pp23[7], pp24[6], pp25[5], S[1401], Cout[1401]);
	Full_Adder FA1356 (pp26[4], pp27[3], pp28[2], S[1402], Cout[1402]);
	Full_Adder FA1357 (pp29[1], pp30[0], Cout[508], S[1403], Cout[1403]);
	Full_Adder FA1358 (Cout[509], S[510], S[511], S[1404], Cout[1404]);
	Full_Adder FA1359 (pp11[20], pp12[19], pp13[18], S[1405], Cout[1405]);
	Full_Adder FA1360 (pp14[17], pp15[16], pp16[15], S[1406], Cout[1406]);
	Full_Adder FA1361 (pp17[14], pp18[13], pp19[12], S[1407], Cout[1407]);
	Full_Adder FA1362 (pp20[11], pp21[10], pp22[9], S[1408], Cout[1408]);
	Full_Adder FA1363 (pp23[8], pp24[7], pp25[6], S[1409], Cout[1409]);
	Full_Adder FA1364 (pp26[5], pp27[4], pp28[3], S[1410], Cout[1410]);
	Full_Adder FA1365 (pp29[2], pp30[1], pp31[0], S[1411], Cout[1411]);
	Full_Adder FA1366 (Cout[510], Cout[511], Cout[512], S[1412], Cout[1412]);
	Full_Adder FA1367 (S[513], S[514], S[515], S[1413], Cout[1413]);
	Full_Adder FA1368 (pp14[18], pp15[17], pp16[16], S[1414], Cout[1414]);
	Full_Adder FA1369 (pp17[15], pp18[14], pp19[13], S[1415], Cout[1415]);
	Full_Adder FA1370 (pp20[12], pp21[11], pp22[10], S[1416], Cout[1416]);
	Full_Adder FA1371 (pp23[9], pp24[8], pp25[7], S[1417], Cout[1417]);
	Full_Adder FA1372 (pp26[6], pp27[5], pp28[4], S[1418], Cout[1418]);
	Full_Adder FA1373 (pp29[3], pp30[2], pp31[1], S[1419], Cout[1419]);
	Full_Adder FA1374 (pp32[0], Cout[513], Cout[514], S[1420], Cout[1420]);
	Full_Adder FA1375 (Cout[515], Cout[516], S[517], S[1421], Cout[1421]);
	Full_Adder FA1376 (S[518], S[519], S[520], S[1422], Cout[1422]);
	Full_Adder FA1377 (pp17[16], pp18[15], pp19[14], S[1423], Cout[1423]);
	Full_Adder FA1378 (pp20[13], pp21[12], pp22[11], S[1424], Cout[1424]);
	Full_Adder FA1379 (pp23[10], pp24[9], pp25[8], S[1425], Cout[1425]);
	Full_Adder FA1380 (pp26[7], pp27[6], pp28[5], S[1426], Cout[1426]);
	Full_Adder FA1381 (pp29[4], pp30[3], pp31[2], S[1427], Cout[1427]);
	Full_Adder FA1382 (pp32[1], pp33[0], Cout[517], S[1428], Cout[1428]);
	Full_Adder FA1383 (Cout[518], Cout[519], Cout[520], S[1429], Cout[1429]);
	Full_Adder FA1384 (Cout[521], S[522], S[523], S[1430], Cout[1430]);
	Full_Adder FA1385 (S[524], S[525], S[526], S[1431], Cout[1431]);
	Full_Adder FA1386 (pp20[14], pp21[13], pp22[12], S[1432], Cout[1432]);
	Full_Adder FA1387 (pp23[11], pp24[10], pp25[9], S[1433], Cout[1433]);
	Full_Adder FA1388 (pp26[8], pp27[7], pp28[6], S[1434], Cout[1434]);
	Full_Adder FA1389 (pp29[5], pp30[4], pp31[3], S[1435], Cout[1435]);
	Full_Adder FA1390 (pp32[2], pp33[1], pp34[0], S[1436], Cout[1436]);
	Full_Adder FA1391 (Cout[522], Cout[523], Cout[524], S[1437], Cout[1437]);
	Full_Adder FA1392 (Cout[525], Cout[526], Cout[527], S[1438], Cout[1438]);
	Full_Adder FA1393 (S[528], S[529], S[530], S[1439], Cout[1439]);
	Full_Adder FA1394 (S[531], S[532], S[533], S[1440], Cout[1440]);
	Full_Adder FA1395 (pp23[12], pp24[11], pp25[10], S[1441], Cout[1441]);
	Full_Adder FA1396 (pp26[9], pp27[8], pp28[7], S[1442], Cout[1442]);
	Full_Adder FA1397 (pp29[6], pp30[5], pp31[4], S[1443], Cout[1443]);
	Full_Adder FA1398 (pp32[3], pp33[2], pp34[1], S[1444], Cout[1444]);
	Full_Adder FA1399 (pp35[0], Cout[528], Cout[529], S[1445], Cout[1445]);
	Full_Adder FA1400 (Cout[530], Cout[531], Cout[532], S[1446], Cout[1446]);
	Full_Adder FA1401 (Cout[533], Cout[534], S[535], S[1447], Cout[1447]);
	Full_Adder FA1402 (S[536], S[537], S[538], S[1448], Cout[1448]);
	Full_Adder FA1403 (S[539], S[540], S[541], S[1449], Cout[1449]);
	Full_Adder FA1404 (pp26[10], pp27[9], pp28[8], S[1450], Cout[1450]);
	Full_Adder FA1405 (pp29[7], pp30[6], pp31[5], S[1451], Cout[1451]);
	Full_Adder FA1406 (pp32[4], pp33[3], pp34[2], S[1452], Cout[1452]);
	Full_Adder FA1407 (pp35[1], pp36[0], Cout[535], S[1453], Cout[1453]);
	Full_Adder FA1408 (Cout[536], Cout[537], Cout[538], S[1454], Cout[1454]);
	Full_Adder FA1409 (Cout[539], Cout[540], Cout[541], S[1455], Cout[1455]);
	Full_Adder FA1410 (Cout[542], S[543], S[544], S[1456], Cout[1456]);
	Full_Adder FA1411 (S[545], S[546], S[547], S[1457], Cout[1457]);
	Full_Adder FA1412 (S[548], S[549], S[550], S[1458], Cout[1458]);
	Full_Adder FA1413 (pp29[8], pp30[7], pp31[6], S[1459], Cout[1459]);
	Full_Adder FA1414 (pp32[5], pp33[4], pp34[3], S[1460], Cout[1460]);
	Full_Adder FA1415 (pp35[2], pp36[1], pp37[0], S[1461], Cout[1461]);
	Full_Adder FA1416 (Cout[543], Cout[544], Cout[545], S[1462], Cout[1462]);
	Full_Adder FA1417 (Cout[546], Cout[547], Cout[548], S[1463], Cout[1463]);
	Full_Adder FA1418 (Cout[549], Cout[550], Cout[551], S[1464], Cout[1464]);
	Full_Adder FA1419 (S[552], S[553], S[554], S[1465], Cout[1465]);
	Full_Adder FA1420 (S[555], S[556], S[557], S[1466], Cout[1466]);
	Full_Adder FA1421 (S[558], S[559], S[560], S[1467], Cout[1467]);
	Full_Adder FA1422 (pp32[6], pp33[5], pp34[4], S[1468], Cout[1468]);
	Full_Adder FA1423 (pp35[3], pp36[2], pp37[1], S[1469], Cout[1469]);
	Full_Adder FA1424 (pp38[0], Cout[552], Cout[553], S[1470], Cout[1470]);
	Full_Adder FA1425 (Cout[554], Cout[555], Cout[556], S[1471], Cout[1471]);
	Full_Adder FA1426 (Cout[557], Cout[558], Cout[559], S[1472], Cout[1472]);
	Full_Adder FA1427 (Cout[560], Cout[561], S[562], S[1473], Cout[1473]);
	Full_Adder FA1428 (S[563], S[564], S[565], S[1474], Cout[1474]);
	Full_Adder FA1429 (S[566], S[567], S[568], S[1475], Cout[1475]);
	Full_Adder FA1430 (S[569], S[570], S[571], S[1476], Cout[1476]);
	Full_Adder FA1431 (pp35[4], pp36[3], pp37[2], S[1477], Cout[1477]);
	Full_Adder FA1432 (pp38[1], pp39[0], Cout[562], S[1478], Cout[1478]);
	Full_Adder FA1433 (Cout[563], Cout[564], Cout[565], S[1479], Cout[1479]);
	Full_Adder FA1434 (Cout[566], Cout[567], Cout[568], S[1480], Cout[1480]);
	Full_Adder FA1435 (Cout[569], Cout[570], Cout[571], S[1481], Cout[1481]);
	Full_Adder FA1436 (Cout[572], S[573], S[574], S[1482], Cout[1482]);
	Full_Adder FA1437 (S[575], S[576], S[577], S[1483], Cout[1483]);
	Full_Adder FA1438 (S[578], S[579], S[580], S[1484], Cout[1484]);
	Full_Adder FA1439 (S[581], S[582], S[583], S[1485], Cout[1485]);
	Full_Adder FA1440 (pp38[2], pp39[1], pp40[0], S[1486], Cout[1486]);
	Full_Adder FA1441 (Cout[573], Cout[574], Cout[575], S[1487], Cout[1487]);
	Full_Adder FA1442 (Cout[576], Cout[577], Cout[578], S[1488], Cout[1488]);
	Full_Adder FA1443 (Cout[579], Cout[580], Cout[581], S[1489], Cout[1489]);
	Full_Adder FA1444 (Cout[582], Cout[583], Cout[584], S[1490], Cout[1490]);
	Full_Adder FA1445 (S[585], S[586], S[587], S[1491], Cout[1491]);
	Full_Adder FA1446 (S[588], S[589], S[590], S[1492], Cout[1492]);
	Full_Adder FA1447 (S[591], S[592], S[593], S[1493], Cout[1493]);
	Full_Adder FA1448 (S[594], S[595], S[596], S[1494], Cout[1494]);
	Full_Adder FA1449 (pp41[0], Cout[585], Cout[586], S[1495], Cout[1495]);
	Full_Adder FA1450 (Cout[587], Cout[588], Cout[589], S[1496], Cout[1496]);
	Full_Adder FA1451 (Cout[590], Cout[591], Cout[592], S[1497], Cout[1497]);
	Full_Adder FA1452 (Cout[593], Cout[594], Cout[595], S[1498], Cout[1498]);
	Full_Adder FA1453 (Cout[596], Cout[597], S[598], S[1499], Cout[1499]);
	Full_Adder FA1454 (S[599], S[600], S[601], S[1500], Cout[1500]);
	Full_Adder FA1455 (S[602], S[603], S[604], S[1501], Cout[1501]);
	Full_Adder FA1456 (S[605], S[606], S[607], S[1502], Cout[1502]);
	Full_Adder FA1457 (S[608], S[609], S[610], S[1503], Cout[1503]);
	Full_Adder FA1458 (Cout[598], Cout[599], Cout[600], S[1504], Cout[1504]);
	Full_Adder FA1459 (Cout[601], Cout[602], Cout[603], S[1505], Cout[1505]);
	Full_Adder FA1460 (Cout[604], Cout[605], Cout[606], S[1506], Cout[1506]);
	Full_Adder FA1461 (Cout[607], Cout[608], Cout[609], S[1507], Cout[1507]);
	Full_Adder FA1462 (Cout[610], Cout[611], S[612], S[1508], Cout[1508]);
	Full_Adder FA1463 (S[613], S[614], S[615], S[1509], Cout[1509]);
	Full_Adder FA1464 (S[616], S[617], S[618], S[1510], Cout[1510]);
	Full_Adder FA1465 (S[619], S[620], S[621], S[1511], Cout[1511]);
	Full_Adder FA1466 (S[622], S[623], S[624], S[1512], Cout[1512]);
	Full_Adder FA1467 (Cout[612], Cout[613], Cout[614], S[1513], Cout[1513]);
	Full_Adder FA1468 (Cout[615], Cout[616], Cout[617], S[1514], Cout[1514]);
	Full_Adder FA1469 (Cout[618], Cout[619], Cout[620], S[1515], Cout[1515]);
	Full_Adder FA1470 (Cout[621], Cout[622], Cout[623], S[1516], Cout[1516]);
	Full_Adder FA1471 (Cout[624], Cout[625], S[626], S[1517], Cout[1517]);
	Full_Adder FA1472 (S[627], S[628], S[629], S[1518], Cout[1518]);
	Full_Adder FA1473 (S[630], S[631], S[632], S[1519], Cout[1519]);
	Full_Adder FA1474 (S[633], S[634], S[635], S[1520], Cout[1520]);
	Full_Adder FA1475 (S[636], S[637], S[638], S[1521], Cout[1521]);
	Full_Adder FA1476 (Cout[626], Cout[627], Cout[628], S[1522], Cout[1522]);
	Full_Adder FA1477 (Cout[629], Cout[630], Cout[631], S[1523], Cout[1523]);
	Full_Adder FA1478 (Cout[632], Cout[633], Cout[634], S[1524], Cout[1524]);
	Full_Adder FA1479 (Cout[635], Cout[636], Cout[637], S[1525], Cout[1525]);
	Full_Adder FA1480 (Cout[638], Cout[639], S[640], S[1526], Cout[1526]);
	Full_Adder FA1481 (S[641], S[642], S[643], S[1527], Cout[1527]);
	Full_Adder FA1482 (S[644], S[645], S[646], S[1528], Cout[1528]);
	Full_Adder FA1483 (S[647], S[648], S[649], S[1529], Cout[1529]);
	Full_Adder FA1484 (S[650], S[651], S[652], S[1530], Cout[1530]);
	Full_Adder FA1485 (Cout[640], Cout[641], Cout[642], S[1531], Cout[1531]);
	Full_Adder FA1486 (Cout[643], Cout[644], Cout[645], S[1532], Cout[1532]);
	Full_Adder FA1487 (Cout[646], Cout[647], Cout[648], S[1533], Cout[1533]);
	Full_Adder FA1488 (Cout[649], Cout[650], Cout[651], S[1534], Cout[1534]);
	Full_Adder FA1489 (Cout[652], Cout[653], S[654], S[1535], Cout[1535]);
	Full_Adder FA1490 (S[655], S[656], S[657], S[1536], Cout[1536]);
	Full_Adder FA1491 (S[658], S[659], S[660], S[1537], Cout[1537]);
	Full_Adder FA1492 (S[661], S[662], S[663], S[1538], Cout[1538]);
	Full_Adder FA1493 (S[664], S[665], S[666], S[1539], Cout[1539]);
	Full_Adder FA1494 (Cout[654], Cout[655], Cout[656], S[1540], Cout[1540]);
	Full_Adder FA1495 (Cout[657], Cout[658], Cout[659], S[1541], Cout[1541]);
	Full_Adder FA1496 (Cout[660], Cout[661], Cout[662], S[1542], Cout[1542]);
	Full_Adder FA1497 (Cout[663], Cout[664], Cout[665], S[1543], Cout[1543]);
	Full_Adder FA1498 (Cout[666], Cout[667], S[668], S[1544], Cout[1544]);
	Full_Adder FA1499 (S[669], S[670], S[671], S[1545], Cout[1545]);
	Full_Adder FA1500 (S[672], S[673], S[674], S[1546], Cout[1546]);
	Full_Adder FA1501 (S[675], S[676], S[677], S[1547], Cout[1547]);
	Full_Adder FA1502 (S[678], S[679], S[680], S[1548], Cout[1548]);
	Full_Adder FA1503 (Cout[668], Cout[669], Cout[670], S[1549], Cout[1549]);
	Full_Adder FA1504 (Cout[671], Cout[672], Cout[673], S[1550], Cout[1550]);
	Full_Adder FA1505 (Cout[674], Cout[675], Cout[676], S[1551], Cout[1551]);
	Full_Adder FA1506 (Cout[677], Cout[678], Cout[679], S[1552], Cout[1552]);
	Full_Adder FA1507 (Cout[680], Cout[681], S[682], S[1553], Cout[1553]);
	Full_Adder FA1508 (S[683], S[684], S[685], S[1554], Cout[1554]);
	Full_Adder FA1509 (S[686], S[687], S[688], S[1555], Cout[1555]);
	Full_Adder FA1510 (S[689], S[690], S[691], S[1556], Cout[1556]);
	Full_Adder FA1511 (S[692], S[693], S[694], S[1557], Cout[1557]);
	Full_Adder FA1512 (Cout[682], Cout[683], Cout[684], S[1558], Cout[1558]);
	Full_Adder FA1513 (Cout[685], Cout[686], Cout[687], S[1559], Cout[1559]);
	Full_Adder FA1514 (Cout[688], Cout[689], Cout[690], S[1560], Cout[1560]);
	Full_Adder FA1515 (Cout[691], Cout[692], Cout[693], S[1561], Cout[1561]);
	Full_Adder FA1516 (Cout[694], Cout[695], S[696], S[1562], Cout[1562]);
	Full_Adder FA1517 (S[697], S[698], S[699], S[1563], Cout[1563]);
	Full_Adder FA1518 (S[700], S[701], S[702], S[1564], Cout[1564]);
	Full_Adder FA1519 (S[703], S[704], S[705], S[1565], Cout[1565]);
	Full_Adder FA1520 (S[706], S[707], S[708], S[1566], Cout[1566]);
	Full_Adder FA1521 (Cout[696], Cout[697], Cout[698], S[1567], Cout[1567]);
	Full_Adder FA1522 (Cout[699], Cout[700], Cout[701], S[1568], Cout[1568]);
	Full_Adder FA1523 (Cout[702], Cout[703], Cout[704], S[1569], Cout[1569]);
	Full_Adder FA1524 (Cout[705], Cout[706], Cout[707], S[1570], Cout[1570]);
	Full_Adder FA1525 (Cout[708], Cout[709], S[710], S[1571], Cout[1571]);
	Full_Adder FA1526 (S[711], S[712], S[713], S[1572], Cout[1572]);
	Full_Adder FA1527 (S[714], S[715], S[716], S[1573], Cout[1573]);
	Full_Adder FA1528 (S[717], S[718], S[719], S[1574], Cout[1574]);
	Full_Adder FA1529 (S[720], S[721], S[722], S[1575], Cout[1575]);
	Full_Adder FA1530 (Cout[710], Cout[711], Cout[712], S[1576], Cout[1576]);
	Full_Adder FA1531 (Cout[713], Cout[714], Cout[715], S[1577], Cout[1577]);
	Full_Adder FA1532 (Cout[716], Cout[717], Cout[718], S[1578], Cout[1578]);
	Full_Adder FA1533 (Cout[719], Cout[720], Cout[721], S[1579], Cout[1579]);
	Full_Adder FA1534 (Cout[722], Cout[723], S[724], S[1580], Cout[1580]);
	Full_Adder FA1535 (S[725], S[726], S[727], S[1581], Cout[1581]);
	Full_Adder FA1536 (S[728], S[729], S[730], S[1582], Cout[1582]);
	Full_Adder FA1537 (S[731], S[732], S[733], S[1583], Cout[1583]);
	Full_Adder FA1538 (S[734], S[735], S[736], S[1584], Cout[1584]);
	Full_Adder FA1539 (Cout[724], Cout[725], Cout[726], S[1585], Cout[1585]);
	Full_Adder FA1540 (Cout[727], Cout[728], Cout[729], S[1586], Cout[1586]);
	Full_Adder FA1541 (Cout[730], Cout[731], Cout[732], S[1587], Cout[1587]);
	Full_Adder FA1542 (Cout[733], Cout[734], Cout[735], S[1588], Cout[1588]);
	Full_Adder FA1543 (Cout[736], Cout[737], S[738], S[1589], Cout[1589]);
	Full_Adder FA1544 (S[739], S[740], S[741], S[1590], Cout[1590]);
	Full_Adder FA1545 (S[742], S[743], S[744], S[1591], Cout[1591]);
	Full_Adder FA1546 (S[745], S[746], S[747], S[1592], Cout[1592]);
	Full_Adder FA1547 (S[748], S[749], S[750], S[1593], Cout[1593]);
	Full_Adder FA1548 (Cout[738], Cout[739], Cout[740], S[1594], Cout[1594]);
	Full_Adder FA1549 (Cout[741], Cout[742], Cout[743], S[1595], Cout[1595]);
	Full_Adder FA1550 (Cout[744], Cout[745], Cout[746], S[1596], Cout[1596]);
	Full_Adder FA1551 (Cout[747], Cout[748], Cout[749], S[1597], Cout[1597]);
	Full_Adder FA1552 (Cout[750], Cout[751], S[752], S[1598], Cout[1598]);
	Full_Adder FA1553 (S[753], S[754], S[755], S[1599], Cout[1599]);
	Full_Adder FA1554 (S[756], S[757], S[758], S[1600], Cout[1600]);
	Full_Adder FA1555 (S[759], S[760], S[761], S[1601], Cout[1601]);
	Full_Adder FA1556 (S[762], S[763], S[764], S[1602], Cout[1602]);
	Full_Adder FA1557 (Cout[752], Cout[753], Cout[754], S[1603], Cout[1603]);
	Full_Adder FA1558 (Cout[755], Cout[756], Cout[757], S[1604], Cout[1604]);
	Full_Adder FA1559 (Cout[758], Cout[759], Cout[760], S[1605], Cout[1605]);
	Full_Adder FA1560 (Cout[761], Cout[762], Cout[763], S[1606], Cout[1606]);
	Full_Adder FA1561 (Cout[764], Cout[765], S[766], S[1607], Cout[1607]);
	Full_Adder FA1562 (S[767], S[768], S[769], S[1608], Cout[1608]);
	Full_Adder FA1563 (S[770], S[771], S[772], S[1609], Cout[1609]);
	Full_Adder FA1564 (S[773], S[774], S[775], S[1610], Cout[1610]);
	Full_Adder FA1565 (S[776], S[777], S[778], S[1611], Cout[1611]);
	Full_Adder FA1566 (Cout[766], Cout[767], Cout[768], S[1612], Cout[1612]);
	Full_Adder FA1567 (Cout[769], Cout[770], Cout[771], S[1613], Cout[1613]);
	Full_Adder FA1568 (Cout[772], Cout[773], Cout[774], S[1614], Cout[1614]);
	Full_Adder FA1569 (Cout[775], Cout[776], Cout[777], S[1615], Cout[1615]);
	Full_Adder FA1570 (Cout[778], Cout[779], S[780], S[1616], Cout[1616]);
	Full_Adder FA1571 (S[781], S[782], S[783], S[1617], Cout[1617]);
	Full_Adder FA1572 (S[784], S[785], S[786], S[1618], Cout[1618]);
	Full_Adder FA1573 (S[787], S[788], S[789], S[1619], Cout[1619]);
	Full_Adder FA1574 (S[790], S[791], S[792], S[1620], Cout[1620]);
	Full_Adder FA1575 (Cout[780], Cout[781], Cout[782], S[1621], Cout[1621]);
	Full_Adder FA1576 (Cout[783], Cout[784], Cout[785], S[1622], Cout[1622]);
	Full_Adder FA1577 (Cout[786], Cout[787], Cout[788], S[1623], Cout[1623]);
	Full_Adder FA1578 (Cout[789], Cout[790], Cout[791], S[1624], Cout[1624]);
	Full_Adder FA1579 (Cout[792], Cout[793], S[794], S[1625], Cout[1625]);
	Full_Adder FA1580 (S[795], S[796], S[797], S[1626], Cout[1626]);
	Full_Adder FA1581 (S[798], S[799], S[800], S[1627], Cout[1627]);
	Full_Adder FA1582 (S[801], S[802], S[803], S[1628], Cout[1628]);
	Full_Adder FA1583 (S[804], S[805], S[806], S[1629], Cout[1629]);
	Full_Adder FA1584 (Cout[794], Cout[795], Cout[796], S[1630], Cout[1630]);
	Full_Adder FA1585 (Cout[797], Cout[798], Cout[799], S[1631], Cout[1631]);
	Full_Adder FA1586 (Cout[800], Cout[801], Cout[802], S[1632], Cout[1632]);
	Full_Adder FA1587 (Cout[803], Cout[804], Cout[805], S[1633], Cout[1633]);
	Full_Adder FA1588 (Cout[806], Cout[807], S[808], S[1634], Cout[1634]);
	Full_Adder FA1589 (S[809], S[810], S[811], S[1635], Cout[1635]);
	Full_Adder FA1590 (S[812], S[813], S[814], S[1636], Cout[1636]);
	Full_Adder FA1591 (S[815], S[816], S[817], S[1637], Cout[1637]);
	Full_Adder FA1592 (S[818], S[819], S[820], S[1638], Cout[1638]);
	Full_Adder FA1593 (Cout[808], Cout[809], Cout[810], S[1639], Cout[1639]);
	Full_Adder FA1594 (Cout[811], Cout[812], Cout[813], S[1640], Cout[1640]);
	Full_Adder FA1595 (Cout[814], Cout[815], Cout[816], S[1641], Cout[1641]);
	Full_Adder FA1596 (Cout[817], Cout[818], Cout[819], S[1642], Cout[1642]);
	Full_Adder FA1597 (Cout[820], Cout[821], S[822], S[1643], Cout[1643]);
	Full_Adder FA1598 (S[823], S[824], S[825], S[1644], Cout[1644]);
	Full_Adder FA1599 (S[826], S[827], S[828], S[1645], Cout[1645]);
	Full_Adder FA1600 (S[829], S[830], S[831], S[1646], Cout[1646]);
	Full_Adder FA1601 (S[832], S[833], S[834], S[1647], Cout[1647]);
	Full_Adder FA1602 (Cout[822], Cout[823], Cout[824], S[1648], Cout[1648]);
	Full_Adder FA1603 (Cout[825], Cout[826], Cout[827], S[1649], Cout[1649]);
	Full_Adder FA1604 (Cout[828], Cout[829], Cout[830], S[1650], Cout[1650]);
	Full_Adder FA1605 (Cout[831], Cout[832], Cout[833], S[1651], Cout[1651]);
	Full_Adder FA1606 (Cout[834], Cout[835], S[836], S[1652], Cout[1652]);
	Full_Adder FA1607 (S[837], S[838], S[839], S[1653], Cout[1653]);
	Full_Adder FA1608 (S[840], S[841], S[842], S[1654], Cout[1654]);
	Full_Adder FA1609 (S[843], S[844], S[845], S[1655], Cout[1655]);
	Full_Adder FA1610 (S[846], S[847], S[848], S[1656], Cout[1656]);
	Full_Adder FA1611 (Cout[836], Cout[837], Cout[838], S[1657], Cout[1657]);
	Full_Adder FA1612 (Cout[839], Cout[840], Cout[841], S[1658], Cout[1658]);
	Full_Adder FA1613 (Cout[842], Cout[843], Cout[844], S[1659], Cout[1659]);
	Full_Adder FA1614 (Cout[845], Cout[846], Cout[847], S[1660], Cout[1660]);
	Full_Adder FA1615 (Cout[848], Cout[849], S[850], S[1661], Cout[1661]);
	Full_Adder FA1616 (S[851], S[852], S[853], S[1662], Cout[1662]);
	Full_Adder FA1617 (S[854], S[855], S[856], S[1663], Cout[1663]);
	Full_Adder FA1618 (S[857], S[858], S[859], S[1664], Cout[1664]);
	Full_Adder FA1619 (S[860], S[861], S[862], S[1665], Cout[1665]);
	Full_Adder FA1620 (Cout[850], Cout[851], Cout[852], S[1666], Cout[1666]);
	Full_Adder FA1621 (Cout[853], Cout[854], Cout[855], S[1667], Cout[1667]);
	Full_Adder FA1622 (Cout[856], Cout[857], Cout[858], S[1668], Cout[1668]);
	Full_Adder FA1623 (Cout[859], Cout[860], Cout[861], S[1669], Cout[1669]);
	Full_Adder FA1624 (Cout[862], Cout[863], S[864], S[1670], Cout[1670]);
	Full_Adder FA1625 (S[865], S[866], S[867], S[1671], Cout[1671]);
	Full_Adder FA1626 (S[868], S[869], S[870], S[1672], Cout[1672]);
	Full_Adder FA1627 (S[871], S[872], S[873], S[1673], Cout[1673]);
	Full_Adder FA1628 (S[874], S[875], S[876], S[1674], Cout[1674]);
	Full_Adder FA1629 (Cout[864], Cout[865], Cout[866], S[1675], Cout[1675]);
	Full_Adder FA1630 (Cout[867], Cout[868], Cout[869], S[1676], Cout[1676]);
	Full_Adder FA1631 (Cout[870], Cout[871], Cout[872], S[1677], Cout[1677]);
	Full_Adder FA1632 (Cout[873], Cout[874], Cout[875], S[1678], Cout[1678]);
	Full_Adder FA1633 (Cout[876], Cout[877], S[878], S[1679], Cout[1679]);
	Full_Adder FA1634 (S[879], S[880], S[881], S[1680], Cout[1680]);
	Full_Adder FA1635 (S[882], S[883], S[884], S[1681], Cout[1681]);
	Full_Adder FA1636 (S[885], S[886], S[887], S[1682], Cout[1682]);
	Full_Adder FA1637 (S[888], S[889], S[890], S[1683], Cout[1683]);
	Full_Adder FA1638 (Cout[878], Cout[879], Cout[880], S[1684], Cout[1684]);
	Full_Adder FA1639 (Cout[881], Cout[882], Cout[883], S[1685], Cout[1685]);
	Full_Adder FA1640 (Cout[884], Cout[885], Cout[886], S[1686], Cout[1686]);
	Full_Adder FA1641 (Cout[887], Cout[888], Cout[889], S[1687], Cout[1687]);
	Full_Adder FA1642 (Cout[890], Cout[891], S[892], S[1688], Cout[1688]);
	Full_Adder FA1643 (S[893], S[894], S[895], S[1689], Cout[1689]);
	Full_Adder FA1644 (S[896], S[897], S[898], S[1690], Cout[1690]);
	Full_Adder FA1645 (S[899], S[900], S[901], S[1691], Cout[1691]);
	Full_Adder FA1646 (S[902], S[903], S[904], S[1692], Cout[1692]);
	Full_Adder FA1647 (Cout[892], Cout[893], Cout[894], S[1693], Cout[1693]);
	Full_Adder FA1648 (Cout[895], Cout[896], Cout[897], S[1694], Cout[1694]);
	Full_Adder FA1649 (Cout[898], Cout[899], Cout[900], S[1695], Cout[1695]);
	Full_Adder FA1650 (Cout[901], Cout[902], Cout[903], S[1696], Cout[1696]);
	Full_Adder FA1651 (Cout[904], Cout[905], S[906], S[1697], Cout[1697]);
	Full_Adder FA1652 (S[907], S[908], S[909], S[1698], Cout[1698]);
	Full_Adder FA1653 (S[910], S[911], S[912], S[1699], Cout[1699]);
	Full_Adder FA1654 (S[913], S[914], S[915], S[1700], Cout[1700]);
	Full_Adder FA1655 (S[916], S[917], S[918], S[1701], Cout[1701]);
	Full_Adder FA1656 (Cout[906], Cout[907], Cout[908], S[1702], Cout[1702]);
	Full_Adder FA1657 (Cout[909], Cout[910], Cout[911], S[1703], Cout[1703]);
	Full_Adder FA1658 (Cout[912], Cout[913], Cout[914], S[1704], Cout[1704]);
	Full_Adder FA1659 (Cout[915], Cout[916], Cout[917], S[1705], Cout[1705]);
	Full_Adder FA1660 (Cout[918], Cout[919], S[920], S[1706], Cout[1706]);
	Full_Adder FA1661 (S[921], S[922], S[923], S[1707], Cout[1707]);
	Full_Adder FA1662 (S[924], S[925], S[926], S[1708], Cout[1708]);
	Full_Adder FA1663 (S[927], S[928], S[929], S[1709], Cout[1709]);
	Full_Adder FA1664 (S[930], S[931], S[932], S[1710], Cout[1710]);
	Full_Adder FA1665 (Cout[920], Cout[921], Cout[922], S[1711], Cout[1711]);
	Full_Adder FA1666 (Cout[923], Cout[924], Cout[925], S[1712], Cout[1712]);
	Full_Adder FA1667 (Cout[926], Cout[927], Cout[928], S[1713], Cout[1713]);
	Full_Adder FA1668 (Cout[929], Cout[930], Cout[931], S[1714], Cout[1714]);
	Full_Adder FA1669 (Cout[932], Cout[933], S[934], S[1715], Cout[1715]);
	Full_Adder FA1670 (S[935], S[936], S[937], S[1716], Cout[1716]);
	Full_Adder FA1671 (S[938], S[939], S[940], S[1717], Cout[1717]);
	Full_Adder FA1672 (S[941], S[942], S[943], S[1718], Cout[1718]);
	Full_Adder FA1673 (S[944], S[945], S[946], S[1719], Cout[1719]);
	Full_Adder FA1674 (Cout[934], Cout[935], Cout[936], S[1720], Cout[1720]);
	Full_Adder FA1675 (Cout[937], Cout[938], Cout[939], S[1721], Cout[1721]);
	Full_Adder FA1676 (Cout[940], Cout[941], Cout[942], S[1722], Cout[1722]);
	Full_Adder FA1677 (Cout[943], Cout[944], Cout[945], S[1723], Cout[1723]);
	Full_Adder FA1678 (Cout[946], Cout[947], S[948], S[1724], Cout[1724]);
	Full_Adder FA1679 (S[949], S[950], S[951], S[1725], Cout[1725]);
	Full_Adder FA1680 (S[952], S[953], S[954], S[1726], Cout[1726]);
	Full_Adder FA1681 (S[955], S[956], S[957], S[1727], Cout[1727]);
	Full_Adder FA1682 (S[958], S[959], S[960], S[1728], Cout[1728]);
	Full_Adder FA1683 (Cout[948], Cout[949], Cout[950], S[1729], Cout[1729]);
	Full_Adder FA1684 (Cout[951], Cout[952], Cout[953], S[1730], Cout[1730]);
	Full_Adder FA1685 (Cout[954], Cout[955], Cout[956], S[1731], Cout[1731]);
	Full_Adder FA1686 (Cout[957], Cout[958], Cout[959], S[1732], Cout[1732]);
	Full_Adder FA1687 (Cout[960], Cout[961], S[962], S[1733], Cout[1733]);
	Full_Adder FA1688 (S[963], S[964], S[965], S[1734], Cout[1734]);
	Full_Adder FA1689 (S[966], S[967], S[968], S[1735], Cout[1735]);
	Full_Adder FA1690 (S[969], S[970], S[971], S[1736], Cout[1736]);
	Full_Adder FA1691 (S[972], S[973], S[974], S[1737], Cout[1737]);
	Full_Adder FA1692 (Cout[962], Cout[963], Cout[964], S[1738], Cout[1738]);
	Full_Adder FA1693 (Cout[965], Cout[966], Cout[967], S[1739], Cout[1739]);
	Full_Adder FA1694 (Cout[968], Cout[969], Cout[970], S[1740], Cout[1740]);
	Full_Adder FA1695 (Cout[971], Cout[972], Cout[973], S[1741], Cout[1741]);
	Full_Adder FA1696 (Cout[974], Cout[975], S[976], S[1742], Cout[1742]);
	Full_Adder FA1697 (S[977], S[978], S[979], S[1743], Cout[1743]);
	Full_Adder FA1698 (S[980], S[981], S[982], S[1744], Cout[1744]);
	Full_Adder FA1699 (S[983], S[984], S[985], S[1745], Cout[1745]);
	Full_Adder FA1700 (S[986], S[987], S[988], S[1746], Cout[1746]);
	Full_Adder FA1701 (Cout[976], Cout[977], Cout[978], S[1747], Cout[1747]);
	Full_Adder FA1702 (Cout[979], Cout[980], Cout[981], S[1748], Cout[1748]);
	Full_Adder FA1703 (Cout[982], Cout[983], Cout[984], S[1749], Cout[1749]);
	Full_Adder FA1704 (Cout[985], Cout[986], Cout[987], S[1750], Cout[1750]);
	Full_Adder FA1705 (Cout[988], Cout[989], S[990], S[1751], Cout[1751]);
	Full_Adder FA1706 (S[991], S[992], S[993], S[1752], Cout[1752]);
	Full_Adder FA1707 (S[994], S[995], S[996], S[1753], Cout[1753]);
	Full_Adder FA1708 (S[997], S[998], S[999], S[1754], Cout[1754]);
	Full_Adder FA1709 (S[1000], S[1001], S[1002], S[1755], Cout[1755]);
	Full_Adder FA1710 (Cout[990], Cout[991], Cout[992], S[1756], Cout[1756]);
	Full_Adder FA1711 (Cout[993], Cout[994], Cout[995], S[1757], Cout[1757]);
	Full_Adder FA1712 (Cout[996], Cout[997], Cout[998], S[1758], Cout[1758]);
	Full_Adder FA1713 (Cout[999], Cout[1000], Cout[1001], S[1759], Cout[1759]);
	Full_Adder FA1714 (Cout[1002], Cout[1003], S[1004], S[1760], Cout[1760]);
	Full_Adder FA1715 (S[1005], S[1006], S[1007], S[1761], Cout[1761]);
	Full_Adder FA1716 (S[1008], S[1009], S[1010], S[1762], Cout[1762]);
	Full_Adder FA1717 (S[1011], S[1012], S[1013], S[1763], Cout[1763]);
	Full_Adder FA1718 (S[1014], S[1015], S[1016], S[1764], Cout[1764]);
	Full_Adder FA1719 (Cout[1004], Cout[1005], Cout[1006], S[1765], Cout[1765]);
	Full_Adder FA1720 (Cout[1007], Cout[1008], Cout[1009], S[1766], Cout[1766]);
	Full_Adder FA1721 (Cout[1010], Cout[1011], Cout[1012], S[1767], Cout[1767]);
	Full_Adder FA1722 (Cout[1013], Cout[1014], Cout[1015], S[1768], Cout[1768]);
	Full_Adder FA1723 (Cout[1016], Cout[1017], S[1018], S[1769], Cout[1769]);
	Full_Adder FA1724 (S[1019], S[1020], S[1021], S[1770], Cout[1770]);
	Full_Adder FA1725 (S[1022], S[1023], S[1024], S[1771], Cout[1771]);
	Full_Adder FA1726 (S[1025], S[1026], S[1027], S[1772], Cout[1772]);
	Full_Adder FA1727 (S[1028], S[1029], S[1030], S[1773], Cout[1773]);
	Full_Adder FA1728 (Cout[1018], Cout[1019], Cout[1020], S[1774], Cout[1774]);
	Full_Adder FA1729 (Cout[1021], Cout[1022], Cout[1023], S[1775], Cout[1775]);
	Full_Adder FA1730 (Cout[1024], Cout[1025], Cout[1026], S[1776], Cout[1776]);
	Full_Adder FA1731 (Cout[1027], Cout[1028], Cout[1029], S[1777], Cout[1777]);
	Full_Adder FA1732 (Cout[1030], Cout[1031], S[1032], S[1778], Cout[1778]);
	Full_Adder FA1733 (S[1033], S[1034], S[1035], S[1779], Cout[1779]);
	Full_Adder FA1734 (S[1036], S[1037], S[1038], S[1780], Cout[1780]);
	Full_Adder FA1735 (S[1039], S[1040], S[1041], S[1781], Cout[1781]);
	Full_Adder FA1736 (S[1042], S[1043], S[1044], S[1782], Cout[1782]);
	Full_Adder FA1737 (Cout[1032], Cout[1033], Cout[1034], S[1783], Cout[1783]);
	Full_Adder FA1738 (Cout[1035], Cout[1036], Cout[1037], S[1784], Cout[1784]);
	Full_Adder FA1739 (Cout[1038], Cout[1039], Cout[1040], S[1785], Cout[1785]);
	Full_Adder FA1740 (Cout[1041], Cout[1042], Cout[1043], S[1786], Cout[1786]);
	Full_Adder FA1741 (Cout[1044], Cout[1045], S[1046], S[1787], Cout[1787]);
	Full_Adder FA1742 (S[1047], S[1048], S[1049], S[1788], Cout[1788]);
	Full_Adder FA1743 (S[1050], S[1051], S[1052], S[1789], Cout[1789]);
	Full_Adder FA1744 (S[1053], S[1054], S[1055], S[1790], Cout[1790]);
	Full_Adder FA1745 (S[1056], S[1057], S[1058], S[1791], Cout[1791]);
	Full_Adder FA1746 (Cout[1046], Cout[1047], Cout[1048], S[1792], Cout[1792]);
	Full_Adder FA1747 (Cout[1049], Cout[1050], Cout[1051], S[1793], Cout[1793]);
	Full_Adder FA1748 (Cout[1052], Cout[1053], Cout[1054], S[1794], Cout[1794]);
	Full_Adder FA1749 (Cout[1055], Cout[1056], Cout[1057], S[1795], Cout[1795]);
	Full_Adder FA1750 (Cout[1058], Cout[1059], S[1060], S[1796], Cout[1796]);
	Full_Adder FA1751 (S[1061], S[1062], S[1063], S[1797], Cout[1797]);
	Full_Adder FA1752 (S[1064], S[1065], S[1066], S[1798], Cout[1798]);
	Full_Adder FA1753 (S[1067], S[1068], S[1069], S[1799], Cout[1799]);
	Full_Adder FA1754 (S[1070], S[1071], S[1072], S[1800], Cout[1800]);
	Full_Adder FA1755 (Cout[1060], Cout[1061], Cout[1062], S[1801], Cout[1801]);
	Full_Adder FA1756 (Cout[1063], Cout[1064], Cout[1065], S[1802], Cout[1802]);
	Full_Adder FA1757 (Cout[1066], Cout[1067], Cout[1068], S[1803], Cout[1803]);
	Full_Adder FA1758 (Cout[1069], Cout[1070], Cout[1071], S[1804], Cout[1804]);
	Full_Adder FA1759 (Cout[1072], Cout[1073], S[1074], S[1805], Cout[1805]);
	Full_Adder FA1760 (S[1075], S[1076], S[1077], S[1806], Cout[1806]);
	Full_Adder FA1761 (S[1078], S[1079], S[1080], S[1807], Cout[1807]);
	Full_Adder FA1762 (S[1081], S[1082], S[1083], S[1808], Cout[1808]);
	Full_Adder FA1763 (S[1084], S[1085], S[1086], S[1809], Cout[1809]);
	Full_Adder FA1764 (Cout[1074], Cout[1075], Cout[1076], S[1810], Cout[1810]);
	Full_Adder FA1765 (Cout[1077], Cout[1078], Cout[1079], S[1811], Cout[1811]);
	Full_Adder FA1766 (Cout[1080], Cout[1081], Cout[1082], S[1812], Cout[1812]);
	Full_Adder FA1767 (Cout[1083], Cout[1084], Cout[1085], S[1813], Cout[1813]);
	Full_Adder FA1768 (Cout[1086], Cout[1087], S[1088], S[1814], Cout[1814]);
	Full_Adder FA1769 (S[1089], S[1090], S[1091], S[1815], Cout[1815]);
	Full_Adder FA1770 (S[1092], S[1093], S[1094], S[1816], Cout[1816]);
	Full_Adder FA1771 (S[1095], S[1096], S[1097], S[1817], Cout[1817]);
	Full_Adder FA1772 (S[1098], S[1099], S[1100], S[1818], Cout[1818]);
	Full_Adder FA1773 (Cout[1088], Cout[1089], Cout[1090], S[1819], Cout[1819]);
	Full_Adder FA1774 (Cout[1091], Cout[1092], Cout[1093], S[1820], Cout[1820]);
	Full_Adder FA1775 (Cout[1094], Cout[1095], Cout[1096], S[1821], Cout[1821]);
	Full_Adder FA1776 (Cout[1097], Cout[1098], Cout[1099], S[1822], Cout[1822]);
	Full_Adder FA1777 (Cout[1100], Cout[1101], S[1102], S[1823], Cout[1823]);
	Full_Adder FA1778 (S[1103], S[1104], S[1105], S[1824], Cout[1824]);
	Full_Adder FA1779 (S[1106], S[1107], S[1108], S[1825], Cout[1825]);
	Full_Adder FA1780 (S[1109], S[1110], S[1111], S[1826], Cout[1826]);
	Full_Adder FA1781 (S[1112], S[1113], S[1114], S[1827], Cout[1827]);
	Full_Adder FA1782 (Cout[1102], Cout[1103], Cout[1104], S[1828], Cout[1828]);
	Full_Adder FA1783 (Cout[1105], Cout[1106], Cout[1107], S[1829], Cout[1829]);
	Full_Adder FA1784 (Cout[1108], Cout[1109], Cout[1110], S[1830], Cout[1830]);
	Full_Adder FA1785 (Cout[1111], Cout[1112], Cout[1113], S[1831], Cout[1831]);
	Full_Adder FA1786 (Cout[1114], Cout[1115], S[1116], S[1832], Cout[1832]);
	Full_Adder FA1787 (S[1117], S[1118], S[1119], S[1833], Cout[1833]);
	Full_Adder FA1788 (S[1120], S[1121], S[1122], S[1834], Cout[1834]);
	Full_Adder FA1789 (S[1123], S[1124], S[1125], S[1835], Cout[1835]);
	Full_Adder FA1790 (S[1126], S[1127], S[1128], S[1836], Cout[1836]);
	Full_Adder FA1791 (Cout[1116], Cout[1117], Cout[1118], S[1837], Cout[1837]);
	Full_Adder FA1792 (Cout[1119], Cout[1120], Cout[1121], S[1838], Cout[1838]);
	Full_Adder FA1793 (Cout[1122], Cout[1123], Cout[1124], S[1839], Cout[1839]);
	Full_Adder FA1794 (Cout[1125], Cout[1126], Cout[1127], S[1840], Cout[1840]);
	Full_Adder FA1795 (Cout[1128], Cout[1129], S[1130], S[1841], Cout[1841]);
	Full_Adder FA1796 (S[1131], S[1132], S[1133], S[1842], Cout[1842]);
	Full_Adder FA1797 (S[1134], S[1135], S[1136], S[1843], Cout[1843]);
	Full_Adder FA1798 (S[1137], S[1138], S[1139], S[1844], Cout[1844]);
	Full_Adder FA1799 (S[1140], S[1141], S[1142], S[1845], Cout[1845]);
	Full_Adder FA1800 (Cout[1130], Cout[1131], Cout[1132], S[1846], Cout[1846]);
	Full_Adder FA1801 (Cout[1133], Cout[1134], Cout[1135], S[1847], Cout[1847]);
	Full_Adder FA1802 (Cout[1136], Cout[1137], Cout[1138], S[1848], Cout[1848]);
	Full_Adder FA1803 (Cout[1139], Cout[1140], Cout[1141], S[1849], Cout[1849]);
	Full_Adder FA1804 (Cout[1142], Cout[1143], S[1144], S[1850], Cout[1850]);
	Full_Adder FA1805 (S[1145], S[1146], S[1147], S[1851], Cout[1851]);
	Full_Adder FA1806 (S[1148], S[1149], S[1150], S[1852], Cout[1852]);
	Full_Adder FA1807 (S[1151], S[1152], S[1153], S[1853], Cout[1853]);
	Full_Adder FA1808 (S[1154], S[1155], S[1156], S[1854], Cout[1854]);
	Full_Adder FA1809 (Cout[1144], Cout[1145], Cout[1146], S[1855], Cout[1855]);
	Full_Adder FA1810 (Cout[1147], Cout[1148], Cout[1149], S[1856], Cout[1856]);
	Full_Adder FA1811 (Cout[1150], Cout[1151], Cout[1152], S[1857], Cout[1857]);
	Full_Adder FA1812 (Cout[1153], Cout[1154], Cout[1155], S[1858], Cout[1858]);
	Full_Adder FA1813 (Cout[1156], Cout[1157], S[1158], S[1859], Cout[1859]);
	Full_Adder FA1814 (S[1159], S[1160], S[1161], S[1860], Cout[1860]);
	Full_Adder FA1815 (S[1162], S[1163], S[1164], S[1861], Cout[1861]);
	Full_Adder FA1816 (S[1165], S[1166], S[1167], S[1862], Cout[1862]);
	Full_Adder FA1817 (S[1168], S[1169], S[1170], S[1863], Cout[1863]);
	Full_Adder FA1818 (Cout[1158], Cout[1159], Cout[1160], S[1864], Cout[1864]);
	Full_Adder FA1819 (Cout[1161], Cout[1162], Cout[1163], S[1865], Cout[1865]);
	Full_Adder FA1820 (Cout[1164], Cout[1165], Cout[1166], S[1866], Cout[1866]);
	Full_Adder FA1821 (Cout[1167], Cout[1168], Cout[1169], S[1867], Cout[1867]);
	Full_Adder FA1822 (Cout[1170], Cout[1171], S[1172], S[1868], Cout[1868]);
	Full_Adder FA1823 (S[1173], S[1174], S[1175], S[1869], Cout[1869]);
	Full_Adder FA1824 (S[1176], S[1177], S[1178], S[1870], Cout[1870]);
	Full_Adder FA1825 (S[1179], S[1180], S[1181], S[1871], Cout[1871]);
	Full_Adder FA1826 (S[1182], S[1183], S[1184], S[1872], Cout[1872]);
	Full_Adder FA1827 (Cout[1172], Cout[1173], Cout[1174], S[1873], Cout[1873]);
	Full_Adder FA1828 (Cout[1175], Cout[1176], Cout[1177], S[1874], Cout[1874]);
	Full_Adder FA1829 (Cout[1178], Cout[1179], Cout[1180], S[1875], Cout[1875]);
	Full_Adder FA1830 (Cout[1181], Cout[1182], Cout[1183], S[1876], Cout[1876]);
	Full_Adder FA1831 (Cout[1184], Cout[1185], S[1186], S[1877], Cout[1877]);
	Full_Adder FA1832 (S[1187], S[1188], S[1189], S[1878], Cout[1878]);
	Full_Adder FA1833 (S[1190], S[1191], S[1192], S[1879], Cout[1879]);
	Full_Adder FA1834 (S[1193], S[1194], S[1195], S[1880], Cout[1880]);
	Full_Adder FA1835 (S[1196], S[1197], S[1198], S[1881], Cout[1881]);
	Full_Adder FA1836 (Cout[1186], Cout[1187], Cout[1188], S[1882], Cout[1882]);
	Full_Adder FA1837 (Cout[1189], Cout[1190], Cout[1191], S[1883], Cout[1883]);
	Full_Adder FA1838 (Cout[1192], Cout[1193], Cout[1194], S[1884], Cout[1884]);
	Full_Adder FA1839 (Cout[1195], Cout[1196], Cout[1197], S[1885], Cout[1885]);
	Full_Adder FA1840 (Cout[1198], Cout[1199], S[1200], S[1886], Cout[1886]);
	Full_Adder FA1841 (S[1201], S[1202], S[1203], S[1887], Cout[1887]);
	Full_Adder FA1842 (S[1204], S[1205], S[1206], S[1888], Cout[1888]);
	Full_Adder FA1843 (S[1207], S[1208], S[1209], S[1889], Cout[1889]);
	Full_Adder FA1844 (S[1210], S[1211], S[1212], S[1890], Cout[1890]);
	Full_Adder FA1845 (Cout[1200], Cout[1201], Cout[1202], S[1891], Cout[1891]);
	Full_Adder FA1846 (Cout[1203], Cout[1204], Cout[1205], S[1892], Cout[1892]);
	Full_Adder FA1847 (Cout[1206], Cout[1207], Cout[1208], S[1893], Cout[1893]);
	Full_Adder FA1848 (Cout[1209], Cout[1210], Cout[1211], S[1894], Cout[1894]);
	Full_Adder FA1849 (Cout[1212], Cout[1213], S[1214], S[1895], Cout[1895]);
	Full_Adder FA1850 (S[1215], S[1216], S[1217], S[1896], Cout[1896]);
	Full_Adder FA1851 (S[1218], S[1219], S[1220], S[1897], Cout[1897]);
	Full_Adder FA1852 (S[1221], S[1222], S[1223], S[1898], Cout[1898]);
	Full_Adder FA1853 (S[1224], S[1225], S[1226], S[1899], Cout[1899]);
	Full_Adder FA1854 (Cout[1214], Cout[1215], Cout[1216], S[1900], Cout[1900]);
	Full_Adder FA1855 (Cout[1217], Cout[1218], Cout[1219], S[1901], Cout[1901]);
	Full_Adder FA1856 (Cout[1220], Cout[1221], Cout[1222], S[1902], Cout[1902]);
	Full_Adder FA1857 (Cout[1223], Cout[1224], Cout[1225], S[1903], Cout[1903]);
	Full_Adder FA1858 (Cout[1226], Cout[1227], S[1228], S[1904], Cout[1904]);
	Full_Adder FA1859 (S[1229], S[1230], S[1231], S[1905], Cout[1905]);
	Full_Adder FA1860 (S[1232], S[1233], S[1234], S[1906], Cout[1906]);
	Full_Adder FA1861 (S[1235], S[1236], S[1237], S[1907], Cout[1907]);
	Full_Adder FA1862 (S[1238], S[1239], S[1240], S[1908], Cout[1908]);
	Full_Adder FA1863 (pp63[24], Cout[1228], Cout[1229], S[1909], Cout[1909]);
	Full_Adder FA1864 (Cout[1230], Cout[1231], Cout[1232], S[1910], Cout[1910]);
	Full_Adder FA1865 (Cout[1233], Cout[1234], Cout[1235], S[1911], Cout[1911]);
	Full_Adder FA1866 (Cout[1236], Cout[1237], Cout[1238], S[1912], Cout[1912]);
	Full_Adder FA1867 (Cout[1239], Cout[1240], Cout[1241], S[1913], Cout[1913]);
	Full_Adder FA1868 (S[1242], S[1243], S[1244], S[1914], Cout[1914]);
	Full_Adder FA1869 (S[1245], S[1246], S[1247], S[1915], Cout[1915]);
	Full_Adder FA1870 (S[1248], S[1249], S[1250], S[1916], Cout[1916]);
	Full_Adder FA1871 (S[1251], S[1252], S[1253], S[1917], Cout[1917]);
	Full_Adder FA1872 (pp61[27], pp62[26], pp63[25], S[1918], Cout[1918]);
	Full_Adder FA1873 (Cout[1242], Cout[1243], Cout[1244], S[1919], Cout[1919]);
	Full_Adder FA1874 (Cout[1245], Cout[1246], Cout[1247], S[1920], Cout[1920]);
	Full_Adder FA1875 (Cout[1248], Cout[1249], Cout[1250], S[1921], Cout[1921]);
	Full_Adder FA1876 (Cout[1251], Cout[1252], Cout[1253], S[1922], Cout[1922]);
	Full_Adder FA1877 (Cout[1254], S[1255], S[1256], S[1923], Cout[1923]);
	Full_Adder FA1878 (S[1257], S[1258], S[1259], S[1924], Cout[1924]);
	Full_Adder FA1879 (S[1260], S[1261], S[1262], S[1925], Cout[1925]);
	Full_Adder FA1880 (S[1263], S[1264], S[1265], S[1926], Cout[1926]);
	Full_Adder FA1881 (pp59[30], pp60[29], pp61[28], S[1927], Cout[1927]);
	Full_Adder FA1882 (pp62[27], pp63[26], Cout[1255], S[1928], Cout[1928]);
	Full_Adder FA1883 (Cout[1256], Cout[1257], Cout[1258], S[1929], Cout[1929]);
	Full_Adder FA1884 (Cout[1259], Cout[1260], Cout[1261], S[1930], Cout[1930]);
	Full_Adder FA1885 (Cout[1262], Cout[1263], Cout[1264], S[1931], Cout[1931]);
	Full_Adder FA1886 (Cout[1265], Cout[1266], S[1267], S[1932], Cout[1932]);
	Full_Adder FA1887 (S[1268], S[1269], S[1270], S[1933], Cout[1933]);
	Full_Adder FA1888 (S[1271], S[1272], S[1273], S[1934], Cout[1934]);
	Full_Adder FA1889 (S[1274], S[1275], S[1276], S[1935], Cout[1935]);
	Full_Adder FA1890 (pp57[33], pp58[32], pp59[31], S[1936], Cout[1936]);
	Full_Adder FA1891 (pp60[30], pp61[29], pp62[28], S[1937], Cout[1937]);
	Full_Adder FA1892 (pp63[27], Cout[1267], Cout[1268], S[1938], Cout[1938]);
	Full_Adder FA1893 (Cout[1269], Cout[1270], Cout[1271], S[1939], Cout[1939]);
	Full_Adder FA1894 (Cout[1272], Cout[1273], Cout[1274], S[1940], Cout[1940]);
	Full_Adder FA1895 (Cout[1275], Cout[1276], Cout[1277], S[1941], Cout[1941]);
	Full_Adder FA1896 (S[1278], S[1279], S[1280], S[1942], Cout[1942]);
	Full_Adder FA1897 (S[1281], S[1282], S[1283], S[1943], Cout[1943]);
	Full_Adder FA1898 (S[1284], S[1285], S[1286], S[1944], Cout[1944]);
	Full_Adder FA1899 (pp55[36], pp56[35], pp57[34], S[1945], Cout[1945]);
	Full_Adder FA1900 (pp58[33], pp59[32], pp60[31], S[1946], Cout[1946]);
	Full_Adder FA1901 (pp61[30], pp62[29], pp63[28], S[1947], Cout[1947]);
	Full_Adder FA1902 (Cout[1278], Cout[1279], Cout[1280], S[1948], Cout[1948]);
	Full_Adder FA1903 (Cout[1281], Cout[1282], Cout[1283], S[1949], Cout[1949]);
	Full_Adder FA1904 (Cout[1284], Cout[1285], Cout[1286], S[1950], Cout[1950]);
	Full_Adder FA1905 (Cout[1287], S[1288], S[1289], S[1951], Cout[1951]);
	Full_Adder FA1906 (S[1290], S[1291], S[1292], S[1952], Cout[1952]);
	Full_Adder FA1907 (S[1293], S[1294], S[1295], S[1953], Cout[1953]);
	Full_Adder FA1908 (pp53[39], pp54[38], pp55[37], S[1954], Cout[1954]);
	Full_Adder FA1909 (pp56[36], pp57[35], pp58[34], S[1955], Cout[1955]);
	Full_Adder FA1910 (pp59[33], pp60[32], pp61[31], S[1956], Cout[1956]);
	Full_Adder FA1911 (pp62[30], pp63[29], Cout[1288], S[1957], Cout[1957]);
	Full_Adder FA1912 (Cout[1289], Cout[1290], Cout[1291], S[1958], Cout[1958]);
	Full_Adder FA1913 (Cout[1292], Cout[1293], Cout[1294], S[1959], Cout[1959]);
	Full_Adder FA1914 (Cout[1295], Cout[1296], S[1297], S[1960], Cout[1960]);
	Full_Adder FA1915 (S[1298], S[1299], S[1300], S[1961], Cout[1961]);
	Full_Adder FA1916 (S[1301], S[1302], S[1303], S[1962], Cout[1962]);
	Full_Adder FA1917 (pp51[42], pp52[41], pp53[40], S[1963], Cout[1963]);
	Full_Adder FA1918 (pp54[39], pp55[38], pp56[37], S[1964], Cout[1964]);
	Full_Adder FA1919 (pp57[36], pp58[35], pp59[34], S[1965], Cout[1965]);
	Full_Adder FA1920 (pp60[33], pp61[32], pp62[31], S[1966], Cout[1966]);
	Full_Adder FA1921 (pp63[30], Cout[1297], Cout[1298], S[1967], Cout[1967]);
	Full_Adder FA1922 (Cout[1299], Cout[1300], Cout[1301], S[1968], Cout[1968]);
	Full_Adder FA1923 (Cout[1302], Cout[1303], Cout[1304], S[1969], Cout[1969]);
	Full_Adder FA1924 (S[1305], S[1306], S[1307], S[1970], Cout[1970]);
	Full_Adder FA1925 (S[1308], S[1309], S[1310], S[1971], Cout[1971]);
	Full_Adder FA1926 (pp49[45], pp50[44], pp51[43], S[1972], Cout[1972]);
	Full_Adder FA1927 (pp52[42], pp53[41], pp54[40], S[1973], Cout[1973]);
	Full_Adder FA1928 (pp55[39], pp56[38], pp57[37], S[1974], Cout[1974]);
	Full_Adder FA1929 (pp58[36], pp59[35], pp60[34], S[1975], Cout[1975]);
	Full_Adder FA1930 (pp61[33], pp62[32], pp63[31], S[1976], Cout[1976]);
	Full_Adder FA1931 (Cout[1305], Cout[1306], Cout[1307], S[1977], Cout[1977]);
	Full_Adder FA1932 (Cout[1308], Cout[1309], Cout[1310], S[1978], Cout[1978]);
	Full_Adder FA1933 (Cout[1311], S[1312], S[1313], S[1979], Cout[1979]);
	Full_Adder FA1934 (S[1314], S[1315], S[1316], S[1980], Cout[1980]);
	Full_Adder FA1935 (pp47[48], pp48[47], pp49[46], S[1981], Cout[1981]);
	Full_Adder FA1936 (pp50[45], pp51[44], pp52[43], S[1982], Cout[1982]);
	Full_Adder FA1937 (pp53[42], pp54[41], pp55[40], S[1983], Cout[1983]);
	Full_Adder FA1938 (pp56[39], pp57[38], pp58[37], S[1984], Cout[1984]);
	Full_Adder FA1939 (pp59[36], pp60[35], pp61[34], S[1985], Cout[1985]);
	Full_Adder FA1940 (pp62[33], pp63[32], Cout[1312], S[1986], Cout[1986]);
	Full_Adder FA1941 (Cout[1313], Cout[1314], Cout[1315], S[1987], Cout[1987]);
	Full_Adder FA1942 (Cout[1316], Cout[1317], S[1318], S[1988], Cout[1988]);
	Full_Adder FA1943 (S[1319], S[1320], S[1321], S[1989], Cout[1989]);
	Full_Adder FA1944 (pp45[51], pp46[50], pp47[49], S[1990], Cout[1990]);
	Full_Adder FA1945 (pp48[48], pp49[47], pp50[46], S[1991], Cout[1991]);
	Full_Adder FA1946 (pp51[45], pp52[44], pp53[43], S[1992], Cout[1992]);
	Full_Adder FA1947 (pp54[42], pp55[41], pp56[40], S[1993], Cout[1993]);
	Full_Adder FA1948 (pp57[39], pp58[38], pp59[37], S[1994], Cout[1994]);
	Full_Adder FA1949 (pp60[36], pp61[35], pp62[34], S[1995], Cout[1995]);
	Full_Adder FA1950 (pp63[33], Cout[1318], Cout[1319], S[1996], Cout[1996]);
	Full_Adder FA1951 (Cout[1320], Cout[1321], Cout[1322], S[1997], Cout[1997]);
	Full_Adder FA1952 (S[1323], S[1324], S[1325], S[1998], Cout[1998]);
	Full_Adder FA1953 (pp43[54], pp44[53], pp45[52], S[1999], Cout[1999]);
	Full_Adder FA1954 (pp46[51], pp47[50], pp48[49], S[2000], Cout[2000]);
	Full_Adder FA1955 (pp49[48], pp50[47], pp51[46], S[2001], Cout[2001]);
	Full_Adder FA1956 (pp52[45], pp53[44], pp54[43], S[2002], Cout[2002]);
	Full_Adder FA1957 (pp55[42], pp56[41], pp57[40], S[2003], Cout[2003]);
	Full_Adder FA1958 (pp58[39], pp59[38], pp60[37], S[2004], Cout[2004]);
	Full_Adder FA1959 (pp61[36], pp62[35], pp63[34], S[2005], Cout[2005]);
	Full_Adder FA1960 (Cout[1323], Cout[1324], Cout[1325], S[2006], Cout[2006]);
	Full_Adder FA1961 (Cout[1326], S[1327], S[1328], S[2007], Cout[2007]);
	Full_Adder FA1962 (pp41[57], pp42[56], pp43[55], S[2008], Cout[2008]);
	Full_Adder FA1963 (pp44[54], pp45[53], pp46[52], S[2009], Cout[2009]);
	Full_Adder FA1964 (pp47[51], pp48[50], pp49[49], S[2010], Cout[2010]);
	Full_Adder FA1965 (pp50[48], pp51[47], pp52[46], S[2011], Cout[2011]);
	Full_Adder FA1966 (pp53[45], pp54[44], pp55[43], S[2012], Cout[2012]);
	Full_Adder FA1967 (pp56[42], pp57[41], pp58[40], S[2013], Cout[2013]);
	Full_Adder FA1968 (pp59[39], pp60[38], pp61[37], S[2014], Cout[2014]);
	Full_Adder FA1969 (pp62[36], pp63[35], Cout[1327], S[2015], Cout[2015]);
	Full_Adder FA1970 (Cout[1328], Cout[1329], S[1330], S[2016], Cout[2016]);
	Full_Adder FA1971 (pp39[60], pp40[59], pp41[58], S[2017], Cout[2017]);
	Full_Adder FA1972 (pp42[57], pp43[56], pp44[55], S[2018], Cout[2018]);
	Full_Adder FA1973 (pp45[54], pp46[53], pp47[52], S[2019], Cout[2019]);
	Full_Adder FA1974 (pp48[51], pp49[50], pp50[49], S[2020], Cout[2020]);
	Full_Adder FA1975 (pp51[48], pp52[47], pp53[46], S[2021], Cout[2021]);
	Full_Adder FA1976 (pp54[45], pp55[44], pp56[43], S[2022], Cout[2022]);
	Full_Adder FA1977 (pp57[42], pp58[41], pp59[40], S[2023], Cout[2023]);
	Full_Adder FA1978 (pp60[39], pp61[38], pp62[37], S[2024], Cout[2024]);
	Full_Adder FA1979 (pp63[36], Cout[1330], Cout[1331], S[2025], Cout[2025]);
	Full_Adder FA1980 (pp37[63], pp38[62], pp39[61], S[2026], Cout[2026]);
	Full_Adder FA1981 (pp40[60], pp41[59], pp42[58], S[2027], Cout[2027]);
	Full_Adder FA1982 (pp43[57], pp44[56], pp45[55], S[2028], Cout[2028]);
	Full_Adder FA1983 (pp46[54], pp47[53], pp48[52], S[2029], Cout[2029]);
	Full_Adder FA1984 (pp49[51], pp50[50], pp51[49], S[2030], Cout[2030]);
	Full_Adder FA1985 (pp52[48], pp53[47], pp54[46], S[2031], Cout[2031]);
	Full_Adder FA1986 (pp55[45], pp56[44], pp57[43], S[2032], Cout[2032]);
	Full_Adder FA1987 (pp58[42], pp59[41], pp60[40], S[2033], Cout[2033]);
	Full_Adder FA1988 (pp61[39], pp62[38], pp63[37], S[2034], Cout[2034]);
	Full_Adder FA1989 (pp38[63], pp39[62], pp40[61], S[2035], Cout[2035]);
	Full_Adder FA1990 (pp41[60], pp42[59], pp43[58], S[2036], Cout[2036]);
	Full_Adder FA1991 (pp44[57], pp45[56], pp46[55], S[2037], Cout[2037]);
	Full_Adder FA1992 (pp47[54], pp48[53], pp49[52], S[2038], Cout[2038]);
	Full_Adder FA1993 (pp50[51], pp51[50], pp52[49], S[2039], Cout[2039]);
	Full_Adder FA1994 (pp53[48], pp54[47], pp55[46], S[2040], Cout[2040]);
	Full_Adder FA1995 (pp56[45], pp57[44], pp58[43], S[2041], Cout[2041]);
	Full_Adder FA1996 (pp59[42], pp60[41], pp61[40], S[2042], Cout[2042]);
	Full_Adder FA1997 (pp39[63], pp40[62], pp41[61], S[2043], Cout[2043]);
	Full_Adder FA1998 (pp42[60], pp43[59], pp44[58], S[2044], Cout[2044]);
	Full_Adder FA1999 (pp45[57], pp46[56], pp47[55], S[2045], Cout[2045]);
	Full_Adder FA2000 (pp48[54], pp49[53], pp50[52], S[2046], Cout[2046]);
	Full_Adder FA2001 (pp51[51], pp52[50], pp53[49], S[2047], Cout[2047]);
	Full_Adder FA2002 (pp54[48], pp55[47], pp56[46], S[2048], Cout[2048]);
	Full_Adder FA2003 (pp57[45], pp58[44], pp59[43], S[2049], Cout[2049]);
	Full_Adder FA2004 (pp40[63], pp41[62], pp42[61], S[2050], Cout[2050]);
	Full_Adder FA2005 (pp43[60], pp44[59], pp45[58], S[2051], Cout[2051]);
	Full_Adder FA2006 (pp46[57], pp47[56], pp48[55], S[2052], Cout[2052]);
	Full_Adder FA2007 (pp49[54], pp50[53], pp51[52], S[2053], Cout[2053]);
	Full_Adder FA2008 (pp52[51], pp53[50], pp54[49], S[2054], Cout[2054]);
	Full_Adder FA2009 (pp55[48], pp56[47], pp57[46], S[2055], Cout[2055]);
	Full_Adder FA2010 (pp41[63], pp42[62], pp43[61], S[2056], Cout[2056]);
	Full_Adder FA2011 (pp44[60], pp45[59], pp46[58], S[2057], Cout[2057]);
	Full_Adder FA2012 (pp47[57], pp48[56], pp49[55], S[2058], Cout[2058]);
	Full_Adder FA2013 (pp50[54], pp51[53], pp52[52], S[2059], Cout[2059]);
	Full_Adder FA2014 (pp53[51], pp54[50], pp55[49], S[2060], Cout[2060]);
	Full_Adder FA2015 (pp42[63], pp43[62], pp44[61], S[2061], Cout[2061]);
	Full_Adder FA2016 (pp45[60], pp46[59], pp47[58], S[2062], Cout[2062]);
	Full_Adder FA2017 (pp48[57], pp49[56], pp50[55], S[2063], Cout[2063]);
	Full_Adder FA2018 (pp51[54], pp52[53], pp53[52], S[2064], Cout[2064]);
	Full_Adder FA2019 (pp43[63], pp44[62], pp45[61], S[2065], Cout[2065]);
	Full_Adder FA2020 (pp46[60], pp47[59], pp48[58], S[2066], Cout[2066]);
	Full_Adder FA2021 (pp49[57], pp50[56], pp51[55], S[2067], Cout[2067]);
	Full_Adder FA2022 (pp44[63], pp45[62], pp46[61], S[2068], Cout[2068]);
	Full_Adder FA2023 (pp47[60], pp48[59], pp49[58], S[2069], Cout[2069]);
	Full_Adder FA2024 (pp45[63], pp46[62], pp47[61], S[2070], Cout[2070]);
	Half_Adder HA47 (pp0[13], pp1[12], S[2071], Cout[2071]);
	Full_Adder FA2025 (pp0[14], pp1[13], pp2[12], S[2072], Cout[2072]);
	Half_Adder HA48 (pp3[11], pp4[10], S[2073], Cout[2073]);
	Full_Adder FA2026 (pp0[15], pp1[14], pp2[13], S[2074], Cout[2074]);
	Full_Adder FA2027 (pp3[12], pp4[11], pp5[10], S[2075], Cout[2075]);
	Half_Adder HA49 (pp6[9], pp7[8], S[2076], Cout[2076]);
	Full_Adder FA2028 (pp0[16], pp1[15], pp2[14], S[2077], Cout[2077]);
	Full_Adder FA2029 (pp3[13], pp4[12], pp5[11], S[2078], Cout[2078]);
	Full_Adder FA2030 (pp6[10], pp7[9], pp8[8], S[2079], Cout[2079]);
	Half_Adder HA50 (pp9[7], pp10[6], S[2080], Cout[2080]);
	Full_Adder FA2031 (pp0[17], pp1[16], pp2[15], S[2081], Cout[2081]);
	Full_Adder FA2032 (pp3[14], pp4[13], pp5[12], S[2082], Cout[2082]);
	Full_Adder FA2033 (pp6[11], pp7[10], pp8[9], S[2083], Cout[2083]);
	Full_Adder FA2034 (pp9[8], pp10[7], pp11[6], S[2084], Cout[2084]);
	Half_Adder HA51 (pp12[5], pp13[4], S[2085], Cout[2085]);
	Full_Adder FA2035 (pp0[18], pp1[17], pp2[16], S[2086], Cout[2086]);
	Full_Adder FA2036 (pp3[15], pp4[14], pp5[13], S[2087], Cout[2087]);
	Full_Adder FA2037 (pp6[12], pp7[11], pp8[10], S[2088], Cout[2088]);
	Full_Adder FA2038 (pp9[9], pp10[8], pp11[7], S[2089], Cout[2089]);
	Full_Adder FA2039 (pp12[6], pp13[5], pp14[4], S[2090], Cout[2090]);
	Half_Adder HA52 (pp15[3], pp16[2], S[2091], Cout[2091]);
	Full_Adder FA2040 (pp2[17], pp3[16], pp4[15], S[2092], Cout[2092]);
	Full_Adder FA2041 (pp5[14], pp6[13], pp7[12], S[2093], Cout[2093]);
	Full_Adder FA2042 (pp8[11], pp9[10], pp10[9], S[2094], Cout[2094]);
	Full_Adder FA2043 (pp11[8], pp12[7], pp13[6], S[2095], Cout[2095]);
	Full_Adder FA2044 (pp14[5], pp15[4], pp16[3], S[2096], Cout[2096]);
	Full_Adder FA2045 (pp17[2], pp18[1], pp19[0], S[2097], Cout[2097]);
	Full_Adder FA2046 (pp5[15], pp6[14], pp7[13], S[2098], Cout[2098]);
	Full_Adder FA2047 (pp8[12], pp9[11], pp10[10], S[2099], Cout[2099]);
	Full_Adder FA2048 (pp11[9], pp12[8], pp13[7], S[2100], Cout[2100]);
	Full_Adder FA2049 (pp14[6], pp15[5], pp16[4], S[2101], Cout[2101]);
	Full_Adder FA2050 (pp17[3], pp18[2], pp19[1], S[2102], Cout[2102]);
	Full_Adder FA2051 (pp20[0], Cout[1333], S[1334], S[2103], Cout[2103]);
	Full_Adder FA2052 (pp8[13], pp9[12], pp10[11], S[2104], Cout[2104]);
	Full_Adder FA2053 (pp11[10], pp12[9], pp13[8], S[2105], Cout[2105]);
	Full_Adder FA2054 (pp14[7], pp15[6], pp16[5], S[2106], Cout[2106]);
	Full_Adder FA2055 (pp17[4], pp18[3], pp19[2], S[2107], Cout[2107]);
	Full_Adder FA2056 (pp20[1], pp21[0], Cout[1334], S[2108], Cout[2108]);
	Full_Adder FA2057 (Cout[1335], S[1336], S[1337], S[2109], Cout[2109]);
	Full_Adder FA2058 (pp11[11], pp12[10], pp13[9], S[2110], Cout[2110]);
	Full_Adder FA2059 (pp14[8], pp15[7], pp16[6], S[2111], Cout[2111]);
	Full_Adder FA2060 (pp17[5], pp18[4], pp19[3], S[2112], Cout[2112]);
	Full_Adder FA2061 (pp20[2], pp21[1], pp22[0], S[2113], Cout[2113]);
	Full_Adder FA2062 (Cout[1336], Cout[1337], Cout[1338], S[2114], Cout[2114]);
	Full_Adder FA2063 (S[1339], S[1340], S[1341], S[2115], Cout[2115]);
	Full_Adder FA2064 (pp14[9], pp15[8], pp16[7], S[2116], Cout[2116]);
	Full_Adder FA2065 (pp17[6], pp18[5], pp19[4], S[2117], Cout[2117]);
	Full_Adder FA2066 (pp20[3], pp21[2], pp22[1], S[2118], Cout[2118]);
	Full_Adder FA2067 (pp23[0], Cout[1339], Cout[1340], S[2119], Cout[2119]);
	Full_Adder FA2068 (Cout[1341], Cout[1342], S[1343], S[2120], Cout[2120]);
	Full_Adder FA2069 (S[1344], S[1345], S[1346], S[2121], Cout[2121]);
	Full_Adder FA2070 (pp17[7], pp18[6], pp19[5], S[2122], Cout[2122]);
	Full_Adder FA2071 (pp20[4], pp21[3], pp22[2], S[2123], Cout[2123]);
	Full_Adder FA2072 (pp23[1], pp24[0], Cout[1343], S[2124], Cout[2124]);
	Full_Adder FA2073 (Cout[1344], Cout[1345], Cout[1346], S[2125], Cout[2125]);
	Full_Adder FA2074 (Cout[1347], S[1348], S[1349], S[2126], Cout[2126]);
	Full_Adder FA2075 (S[1350], S[1351], S[1352], S[2127], Cout[2127]);
	Full_Adder FA2076 (pp20[5], pp21[4], pp22[3], S[2128], Cout[2128]);
	Full_Adder FA2077 (pp23[2], pp24[1], pp25[0], S[2129], Cout[2129]);
	Full_Adder FA2078 (Cout[1348], Cout[1349], Cout[1350], S[2130], Cout[2130]);
	Full_Adder FA2079 (Cout[1351], Cout[1352], Cout[1353], S[2131], Cout[2131]);
	Full_Adder FA2080 (S[1354], S[1355], S[1356], S[2132], Cout[2132]);
	Full_Adder FA2081 (S[1357], S[1358], S[1359], S[2133], Cout[2133]);
	Full_Adder FA2082 (pp23[3], pp24[2], pp25[1], S[2134], Cout[2134]);
	Full_Adder FA2083 (pp26[0], Cout[1354], Cout[1355], S[2135], Cout[2135]);
	Full_Adder FA2084 (Cout[1356], Cout[1357], Cout[1358], S[2136], Cout[2136]);
	Full_Adder FA2085 (Cout[1359], Cout[1360], S[1361], S[2137], Cout[2137]);
	Full_Adder FA2086 (S[1362], S[1363], S[1364], S[2138], Cout[2138]);
	Full_Adder FA2087 (S[1365], S[1366], S[1367], S[2139], Cout[2139]);
	Full_Adder FA2088 (pp26[1], pp27[0], Cout[1361], S[2140], Cout[2140]);
	Full_Adder FA2089 (Cout[1362], Cout[1363], Cout[1364], S[2141], Cout[2141]);
	Full_Adder FA2090 (Cout[1365], Cout[1366], Cout[1367], S[2142], Cout[2142]);
	Full_Adder FA2091 (Cout[1368], S[1369], S[1370], S[2143], Cout[2143]);
	Full_Adder FA2092 (S[1371], S[1372], S[1373], S[2144], Cout[2144]);
	Full_Adder FA2093 (S[1374], S[1375], S[1376], S[2145], Cout[2145]);
	Full_Adder FA2094 (S[507], Cout[1369], Cout[1370], S[2146], Cout[2146]);
	Full_Adder FA2095 (Cout[1371], Cout[1372], Cout[1373], S[2147], Cout[2147]);
	Full_Adder FA2096 (Cout[1374], Cout[1375], Cout[1376], S[2148], Cout[2148]);
	Full_Adder FA2097 (Cout[1377], S[1378], S[1379], S[2149], Cout[2149]);
	Full_Adder FA2098 (S[1380], S[1381], S[1382], S[2150], Cout[2150]);
	Full_Adder FA2099 (S[1383], S[1384], S[1385], S[2151], Cout[2151]);
	Full_Adder FA2100 (S[509], Cout[1378], Cout[1379], S[2152], Cout[2152]);
	Full_Adder FA2101 (Cout[1380], Cout[1381], Cout[1382], S[2153], Cout[2153]);
	Full_Adder FA2102 (Cout[1383], Cout[1384], Cout[1385], S[2154], Cout[2154]);
	Full_Adder FA2103 (Cout[1386], S[1387], S[1388], S[2155], Cout[2155]);
	Full_Adder FA2104 (S[1389], S[1390], S[1391], S[2156], Cout[2156]);
	Full_Adder FA2105 (S[1392], S[1393], S[1394], S[2157], Cout[2157]);
	Full_Adder FA2106 (S[512], Cout[1387], Cout[1388], S[2158], Cout[2158]);
	Full_Adder FA2107 (Cout[1389], Cout[1390], Cout[1391], S[2159], Cout[2159]);
	Full_Adder FA2108 (Cout[1392], Cout[1393], Cout[1394], S[2160], Cout[2160]);
	Full_Adder FA2109 (Cout[1395], S[1396], S[1397], S[2161], Cout[2161]);
	Full_Adder FA2110 (S[1398], S[1399], S[1400], S[2162], Cout[2162]);
	Full_Adder FA2111 (S[1401], S[1402], S[1403], S[2163], Cout[2163]);
	Full_Adder FA2112 (S[516], Cout[1396], Cout[1397], S[2164], Cout[2164]);
	Full_Adder FA2113 (Cout[1398], Cout[1399], Cout[1400], S[2165], Cout[2165]);
	Full_Adder FA2114 (Cout[1401], Cout[1402], Cout[1403], S[2166], Cout[2166]);
	Full_Adder FA2115 (Cout[1404], S[1405], S[1406], S[2167], Cout[2167]);
	Full_Adder FA2116 (S[1407], S[1408], S[1409], S[2168], Cout[2168]);
	Full_Adder FA2117 (S[1410], S[1411], S[1412], S[2169], Cout[2169]);
	Full_Adder FA2118 (S[521], Cout[1405], Cout[1406], S[2170], Cout[2170]);
	Full_Adder FA2119 (Cout[1407], Cout[1408], Cout[1409], S[2171], Cout[2171]);
	Full_Adder FA2120 (Cout[1410], Cout[1411], Cout[1412], S[2172], Cout[2172]);
	Full_Adder FA2121 (Cout[1413], S[1414], S[1415], S[2173], Cout[2173]);
	Full_Adder FA2122 (S[1416], S[1417], S[1418], S[2174], Cout[2174]);
	Full_Adder FA2123 (S[1419], S[1420], S[1421], S[2175], Cout[2175]);
	Full_Adder FA2124 (S[527], Cout[1414], Cout[1415], S[2176], Cout[2176]);
	Full_Adder FA2125 (Cout[1416], Cout[1417], Cout[1418], S[2177], Cout[2177]);
	Full_Adder FA2126 (Cout[1419], Cout[1420], Cout[1421], S[2178], Cout[2178]);
	Full_Adder FA2127 (Cout[1422], S[1423], S[1424], S[2179], Cout[2179]);
	Full_Adder FA2128 (S[1425], S[1426], S[1427], S[2180], Cout[2180]);
	Full_Adder FA2129 (S[1428], S[1429], S[1430], S[2181], Cout[2181]);
	Full_Adder FA2130 (S[534], Cout[1423], Cout[1424], S[2182], Cout[2182]);
	Full_Adder FA2131 (Cout[1425], Cout[1426], Cout[1427], S[2183], Cout[2183]);
	Full_Adder FA2132 (Cout[1428], Cout[1429], Cout[1430], S[2184], Cout[2184]);
	Full_Adder FA2133 (Cout[1431], S[1432], S[1433], S[2185], Cout[2185]);
	Full_Adder FA2134 (S[1434], S[1435], S[1436], S[2186], Cout[2186]);
	Full_Adder FA2135 (S[1437], S[1438], S[1439], S[2187], Cout[2187]);
	Full_Adder FA2136 (S[542], Cout[1432], Cout[1433], S[2188], Cout[2188]);
	Full_Adder FA2137 (Cout[1434], Cout[1435], Cout[1436], S[2189], Cout[2189]);
	Full_Adder FA2138 (Cout[1437], Cout[1438], Cout[1439], S[2190], Cout[2190]);
	Full_Adder FA2139 (Cout[1440], S[1441], S[1442], S[2191], Cout[2191]);
	Full_Adder FA2140 (S[1443], S[1444], S[1445], S[2192], Cout[2192]);
	Full_Adder FA2141 (S[1446], S[1447], S[1448], S[2193], Cout[2193]);
	Full_Adder FA2142 (S[551], Cout[1441], Cout[1442], S[2194], Cout[2194]);
	Full_Adder FA2143 (Cout[1443], Cout[1444], Cout[1445], S[2195], Cout[2195]);
	Full_Adder FA2144 (Cout[1446], Cout[1447], Cout[1448], S[2196], Cout[2196]);
	Full_Adder FA2145 (Cout[1449], S[1450], S[1451], S[2197], Cout[2197]);
	Full_Adder FA2146 (S[1452], S[1453], S[1454], S[2198], Cout[2198]);
	Full_Adder FA2147 (S[1455], S[1456], S[1457], S[2199], Cout[2199]);
	Full_Adder FA2148 (S[561], Cout[1450], Cout[1451], S[2200], Cout[2200]);
	Full_Adder FA2149 (Cout[1452], Cout[1453], Cout[1454], S[2201], Cout[2201]);
	Full_Adder FA2150 (Cout[1455], Cout[1456], Cout[1457], S[2202], Cout[2202]);
	Full_Adder FA2151 (Cout[1458], S[1459], S[1460], S[2203], Cout[2203]);
	Full_Adder FA2152 (S[1461], S[1462], S[1463], S[2204], Cout[2204]);
	Full_Adder FA2153 (S[1464], S[1465], S[1466], S[2205], Cout[2205]);
	Full_Adder FA2154 (S[572], Cout[1459], Cout[1460], S[2206], Cout[2206]);
	Full_Adder FA2155 (Cout[1461], Cout[1462], Cout[1463], S[2207], Cout[2207]);
	Full_Adder FA2156 (Cout[1464], Cout[1465], Cout[1466], S[2208], Cout[2208]);
	Full_Adder FA2157 (Cout[1467], S[1468], S[1469], S[2209], Cout[2209]);
	Full_Adder FA2158 (S[1470], S[1471], S[1472], S[2210], Cout[2210]);
	Full_Adder FA2159 (S[1473], S[1474], S[1475], S[2211], Cout[2211]);
	Full_Adder FA2160 (S[584], Cout[1468], Cout[1469], S[2212], Cout[2212]);
	Full_Adder FA2161 (Cout[1470], Cout[1471], Cout[1472], S[2213], Cout[2213]);
	Full_Adder FA2162 (Cout[1473], Cout[1474], Cout[1475], S[2214], Cout[2214]);
	Full_Adder FA2163 (Cout[1476], S[1477], S[1478], S[2215], Cout[2215]);
	Full_Adder FA2164 (S[1479], S[1480], S[1481], S[2216], Cout[2216]);
	Full_Adder FA2165 (S[1482], S[1483], S[1484], S[2217], Cout[2217]);
	Full_Adder FA2166 (S[597], Cout[1477], Cout[1478], S[2218], Cout[2218]);
	Full_Adder FA2167 (Cout[1479], Cout[1480], Cout[1481], S[2219], Cout[2219]);
	Full_Adder FA2168 (Cout[1482], Cout[1483], Cout[1484], S[2220], Cout[2220]);
	Full_Adder FA2169 (Cout[1485], S[1486], S[1487], S[2221], Cout[2221]);
	Full_Adder FA2170 (S[1488], S[1489], S[1490], S[2222], Cout[2222]);
	Full_Adder FA2171 (S[1491], S[1492], S[1493], S[2223], Cout[2223]);
	Full_Adder FA2172 (S[611], Cout[1486], Cout[1487], S[2224], Cout[2224]);
	Full_Adder FA2173 (Cout[1488], Cout[1489], Cout[1490], S[2225], Cout[2225]);
	Full_Adder FA2174 (Cout[1491], Cout[1492], Cout[1493], S[2226], Cout[2226]);
	Full_Adder FA2175 (Cout[1494], S[1495], S[1496], S[2227], Cout[2227]);
	Full_Adder FA2176 (S[1497], S[1498], S[1499], S[2228], Cout[2228]);
	Full_Adder FA2177 (S[1500], S[1501], S[1502], S[2229], Cout[2229]);
	Full_Adder FA2178 (S[625], Cout[1495], Cout[1496], S[2230], Cout[2230]);
	Full_Adder FA2179 (Cout[1497], Cout[1498], Cout[1499], S[2231], Cout[2231]);
	Full_Adder FA2180 (Cout[1500], Cout[1501], Cout[1502], S[2232], Cout[2232]);
	Full_Adder FA2181 (Cout[1503], S[1504], S[1505], S[2233], Cout[2233]);
	Full_Adder FA2182 (S[1506], S[1507], S[1508], S[2234], Cout[2234]);
	Full_Adder FA2183 (S[1509], S[1510], S[1511], S[2235], Cout[2235]);
	Full_Adder FA2184 (S[639], Cout[1504], Cout[1505], S[2236], Cout[2236]);
	Full_Adder FA2185 (Cout[1506], Cout[1507], Cout[1508], S[2237], Cout[2237]);
	Full_Adder FA2186 (Cout[1509], Cout[1510], Cout[1511], S[2238], Cout[2238]);
	Full_Adder FA2187 (Cout[1512], S[1513], S[1514], S[2239], Cout[2239]);
	Full_Adder FA2188 (S[1515], S[1516], S[1517], S[2240], Cout[2240]);
	Full_Adder FA2189 (S[1518], S[1519], S[1520], S[2241], Cout[2241]);
	Full_Adder FA2190 (S[653], Cout[1513], Cout[1514], S[2242], Cout[2242]);
	Full_Adder FA2191 (Cout[1515], Cout[1516], Cout[1517], S[2243], Cout[2243]);
	Full_Adder FA2192 (Cout[1518], Cout[1519], Cout[1520], S[2244], Cout[2244]);
	Full_Adder FA2193 (Cout[1521], S[1522], S[1523], S[2245], Cout[2245]);
	Full_Adder FA2194 (S[1524], S[1525], S[1526], S[2246], Cout[2246]);
	Full_Adder FA2195 (S[1527], S[1528], S[1529], S[2247], Cout[2247]);
	Full_Adder FA2196 (S[667], Cout[1522], Cout[1523], S[2248], Cout[2248]);
	Full_Adder FA2197 (Cout[1524], Cout[1525], Cout[1526], S[2249], Cout[2249]);
	Full_Adder FA2198 (Cout[1527], Cout[1528], Cout[1529], S[2250], Cout[2250]);
	Full_Adder FA2199 (Cout[1530], S[1531], S[1532], S[2251], Cout[2251]);
	Full_Adder FA2200 (S[1533], S[1534], S[1535], S[2252], Cout[2252]);
	Full_Adder FA2201 (S[1536], S[1537], S[1538], S[2253], Cout[2253]);
	Full_Adder FA2202 (S[681], Cout[1531], Cout[1532], S[2254], Cout[2254]);
	Full_Adder FA2203 (Cout[1533], Cout[1534], Cout[1535], S[2255], Cout[2255]);
	Full_Adder FA2204 (Cout[1536], Cout[1537], Cout[1538], S[2256], Cout[2256]);
	Full_Adder FA2205 (Cout[1539], S[1540], S[1541], S[2257], Cout[2257]);
	Full_Adder FA2206 (S[1542], S[1543], S[1544], S[2258], Cout[2258]);
	Full_Adder FA2207 (S[1545], S[1546], S[1547], S[2259], Cout[2259]);
	Full_Adder FA2208 (S[695], Cout[1540], Cout[1541], S[2260], Cout[2260]);
	Full_Adder FA2209 (Cout[1542], Cout[1543], Cout[1544], S[2261], Cout[2261]);
	Full_Adder FA2210 (Cout[1545], Cout[1546], Cout[1547], S[2262], Cout[2262]);
	Full_Adder FA2211 (Cout[1548], S[1549], S[1550], S[2263], Cout[2263]);
	Full_Adder FA2212 (S[1551], S[1552], S[1553], S[2264], Cout[2264]);
	Full_Adder FA2213 (S[1554], S[1555], S[1556], S[2265], Cout[2265]);
	Full_Adder FA2214 (S[709], Cout[1549], Cout[1550], S[2266], Cout[2266]);
	Full_Adder FA2215 (Cout[1551], Cout[1552], Cout[1553], S[2267], Cout[2267]);
	Full_Adder FA2216 (Cout[1554], Cout[1555], Cout[1556], S[2268], Cout[2268]);
	Full_Adder FA2217 (Cout[1557], S[1558], S[1559], S[2269], Cout[2269]);
	Full_Adder FA2218 (S[1560], S[1561], S[1562], S[2270], Cout[2270]);
	Full_Adder FA2219 (S[1563], S[1564], S[1565], S[2271], Cout[2271]);
	Full_Adder FA2220 (S[723], Cout[1558], Cout[1559], S[2272], Cout[2272]);
	Full_Adder FA2221 (Cout[1560], Cout[1561], Cout[1562], S[2273], Cout[2273]);
	Full_Adder FA2222 (Cout[1563], Cout[1564], Cout[1565], S[2274], Cout[2274]);
	Full_Adder FA2223 (Cout[1566], S[1567], S[1568], S[2275], Cout[2275]);
	Full_Adder FA2224 (S[1569], S[1570], S[1571], S[2276], Cout[2276]);
	Full_Adder FA2225 (S[1572], S[1573], S[1574], S[2277], Cout[2277]);
	Full_Adder FA2226 (S[737], Cout[1567], Cout[1568], S[2278], Cout[2278]);
	Full_Adder FA2227 (Cout[1569], Cout[1570], Cout[1571], S[2279], Cout[2279]);
	Full_Adder FA2228 (Cout[1572], Cout[1573], Cout[1574], S[2280], Cout[2280]);
	Full_Adder FA2229 (Cout[1575], S[1576], S[1577], S[2281], Cout[2281]);
	Full_Adder FA2230 (S[1578], S[1579], S[1580], S[2282], Cout[2282]);
	Full_Adder FA2231 (S[1581], S[1582], S[1583], S[2283], Cout[2283]);
	Full_Adder FA2232 (S[751], Cout[1576], Cout[1577], S[2284], Cout[2284]);
	Full_Adder FA2233 (Cout[1578], Cout[1579], Cout[1580], S[2285], Cout[2285]);
	Full_Adder FA2234 (Cout[1581], Cout[1582], Cout[1583], S[2286], Cout[2286]);
	Full_Adder FA2235 (Cout[1584], S[1585], S[1586], S[2287], Cout[2287]);
	Full_Adder FA2236 (S[1587], S[1588], S[1589], S[2288], Cout[2288]);
	Full_Adder FA2237 (S[1590], S[1591], S[1592], S[2289], Cout[2289]);
	Full_Adder FA2238 (S[765], Cout[1585], Cout[1586], S[2290], Cout[2290]);
	Full_Adder FA2239 (Cout[1587], Cout[1588], Cout[1589], S[2291], Cout[2291]);
	Full_Adder FA2240 (Cout[1590], Cout[1591], Cout[1592], S[2292], Cout[2292]);
	Full_Adder FA2241 (Cout[1593], S[1594], S[1595], S[2293], Cout[2293]);
	Full_Adder FA2242 (S[1596], S[1597], S[1598], S[2294], Cout[2294]);
	Full_Adder FA2243 (S[1599], S[1600], S[1601], S[2295], Cout[2295]);
	Full_Adder FA2244 (S[779], Cout[1594], Cout[1595], S[2296], Cout[2296]);
	Full_Adder FA2245 (Cout[1596], Cout[1597], Cout[1598], S[2297], Cout[2297]);
	Full_Adder FA2246 (Cout[1599], Cout[1600], Cout[1601], S[2298], Cout[2298]);
	Full_Adder FA2247 (Cout[1602], S[1603], S[1604], S[2299], Cout[2299]);
	Full_Adder FA2248 (S[1605], S[1606], S[1607], S[2300], Cout[2300]);
	Full_Adder FA2249 (S[1608], S[1609], S[1610], S[2301], Cout[2301]);
	Full_Adder FA2250 (S[793], Cout[1603], Cout[1604], S[2302], Cout[2302]);
	Full_Adder FA2251 (Cout[1605], Cout[1606], Cout[1607], S[2303], Cout[2303]);
	Full_Adder FA2252 (Cout[1608], Cout[1609], Cout[1610], S[2304], Cout[2304]);
	Full_Adder FA2253 (Cout[1611], S[1612], S[1613], S[2305], Cout[2305]);
	Full_Adder FA2254 (S[1614], S[1615], S[1616], S[2306], Cout[2306]);
	Full_Adder FA2255 (S[1617], S[1618], S[1619], S[2307], Cout[2307]);
	Full_Adder FA2256 (S[807], Cout[1612], Cout[1613], S[2308], Cout[2308]);
	Full_Adder FA2257 (Cout[1614], Cout[1615], Cout[1616], S[2309], Cout[2309]);
	Full_Adder FA2258 (Cout[1617], Cout[1618], Cout[1619], S[2310], Cout[2310]);
	Full_Adder FA2259 (Cout[1620], S[1621], S[1622], S[2311], Cout[2311]);
	Full_Adder FA2260 (S[1623], S[1624], S[1625], S[2312], Cout[2312]);
	Full_Adder FA2261 (S[1626], S[1627], S[1628], S[2313], Cout[2313]);
	Full_Adder FA2262 (S[821], Cout[1621], Cout[1622], S[2314], Cout[2314]);
	Full_Adder FA2263 (Cout[1623], Cout[1624], Cout[1625], S[2315], Cout[2315]);
	Full_Adder FA2264 (Cout[1626], Cout[1627], Cout[1628], S[2316], Cout[2316]);
	Full_Adder FA2265 (Cout[1629], S[1630], S[1631], S[2317], Cout[2317]);
	Full_Adder FA2266 (S[1632], S[1633], S[1634], S[2318], Cout[2318]);
	Full_Adder FA2267 (S[1635], S[1636], S[1637], S[2319], Cout[2319]);
	Full_Adder FA2268 (S[835], Cout[1630], Cout[1631], S[2320], Cout[2320]);
	Full_Adder FA2269 (Cout[1632], Cout[1633], Cout[1634], S[2321], Cout[2321]);
	Full_Adder FA2270 (Cout[1635], Cout[1636], Cout[1637], S[2322], Cout[2322]);
	Full_Adder FA2271 (Cout[1638], S[1639], S[1640], S[2323], Cout[2323]);
	Full_Adder FA2272 (S[1641], S[1642], S[1643], S[2324], Cout[2324]);
	Full_Adder FA2273 (S[1644], S[1645], S[1646], S[2325], Cout[2325]);
	Full_Adder FA2274 (S[849], Cout[1639], Cout[1640], S[2326], Cout[2326]);
	Full_Adder FA2275 (Cout[1641], Cout[1642], Cout[1643], S[2327], Cout[2327]);
	Full_Adder FA2276 (Cout[1644], Cout[1645], Cout[1646], S[2328], Cout[2328]);
	Full_Adder FA2277 (Cout[1647], S[1648], S[1649], S[2329], Cout[2329]);
	Full_Adder FA2278 (S[1650], S[1651], S[1652], S[2330], Cout[2330]);
	Full_Adder FA2279 (S[1653], S[1654], S[1655], S[2331], Cout[2331]);
	Full_Adder FA2280 (S[863], Cout[1648], Cout[1649], S[2332], Cout[2332]);
	Full_Adder FA2281 (Cout[1650], Cout[1651], Cout[1652], S[2333], Cout[2333]);
	Full_Adder FA2282 (Cout[1653], Cout[1654], Cout[1655], S[2334], Cout[2334]);
	Full_Adder FA2283 (Cout[1656], S[1657], S[1658], S[2335], Cout[2335]);
	Full_Adder FA2284 (S[1659], S[1660], S[1661], S[2336], Cout[2336]);
	Full_Adder FA2285 (S[1662], S[1663], S[1664], S[2337], Cout[2337]);
	Full_Adder FA2286 (S[877], Cout[1657], Cout[1658], S[2338], Cout[2338]);
	Full_Adder FA2287 (Cout[1659], Cout[1660], Cout[1661], S[2339], Cout[2339]);
	Full_Adder FA2288 (Cout[1662], Cout[1663], Cout[1664], S[2340], Cout[2340]);
	Full_Adder FA2289 (Cout[1665], S[1666], S[1667], S[2341], Cout[2341]);
	Full_Adder FA2290 (S[1668], S[1669], S[1670], S[2342], Cout[2342]);
	Full_Adder FA2291 (S[1671], S[1672], S[1673], S[2343], Cout[2343]);
	Full_Adder FA2292 (S[891], Cout[1666], Cout[1667], S[2344], Cout[2344]);
	Full_Adder FA2293 (Cout[1668], Cout[1669], Cout[1670], S[2345], Cout[2345]);
	Full_Adder FA2294 (Cout[1671], Cout[1672], Cout[1673], S[2346], Cout[2346]);
	Full_Adder FA2295 (Cout[1674], S[1675], S[1676], S[2347], Cout[2347]);
	Full_Adder FA2296 (S[1677], S[1678], S[1679], S[2348], Cout[2348]);
	Full_Adder FA2297 (S[1680], S[1681], S[1682], S[2349], Cout[2349]);
	Full_Adder FA2298 (S[905], Cout[1675], Cout[1676], S[2350], Cout[2350]);
	Full_Adder FA2299 (Cout[1677], Cout[1678], Cout[1679], S[2351], Cout[2351]);
	Full_Adder FA2300 (Cout[1680], Cout[1681], Cout[1682], S[2352], Cout[2352]);
	Full_Adder FA2301 (Cout[1683], S[1684], S[1685], S[2353], Cout[2353]);
	Full_Adder FA2302 (S[1686], S[1687], S[1688], S[2354], Cout[2354]);
	Full_Adder FA2303 (S[1689], S[1690], S[1691], S[2355], Cout[2355]);
	Full_Adder FA2304 (S[919], Cout[1684], Cout[1685], S[2356], Cout[2356]);
	Full_Adder FA2305 (Cout[1686], Cout[1687], Cout[1688], S[2357], Cout[2357]);
	Full_Adder FA2306 (Cout[1689], Cout[1690], Cout[1691], S[2358], Cout[2358]);
	Full_Adder FA2307 (Cout[1692], S[1693], S[1694], S[2359], Cout[2359]);
	Full_Adder FA2308 (S[1695], S[1696], S[1697], S[2360], Cout[2360]);
	Full_Adder FA2309 (S[1698], S[1699], S[1700], S[2361], Cout[2361]);
	Full_Adder FA2310 (S[933], Cout[1693], Cout[1694], S[2362], Cout[2362]);
	Full_Adder FA2311 (Cout[1695], Cout[1696], Cout[1697], S[2363], Cout[2363]);
	Full_Adder FA2312 (Cout[1698], Cout[1699], Cout[1700], S[2364], Cout[2364]);
	Full_Adder FA2313 (Cout[1701], S[1702], S[1703], S[2365], Cout[2365]);
	Full_Adder FA2314 (S[1704], S[1705], S[1706], S[2366], Cout[2366]);
	Full_Adder FA2315 (S[1707], S[1708], S[1709], S[2367], Cout[2367]);
	Full_Adder FA2316 (S[947], Cout[1702], Cout[1703], S[2368], Cout[2368]);
	Full_Adder FA2317 (Cout[1704], Cout[1705], Cout[1706], S[2369], Cout[2369]);
	Full_Adder FA2318 (Cout[1707], Cout[1708], Cout[1709], S[2370], Cout[2370]);
	Full_Adder FA2319 (Cout[1710], S[1711], S[1712], S[2371], Cout[2371]);
	Full_Adder FA2320 (S[1713], S[1714], S[1715], S[2372], Cout[2372]);
	Full_Adder FA2321 (S[1716], S[1717], S[1718], S[2373], Cout[2373]);
	Full_Adder FA2322 (S[961], Cout[1711], Cout[1712], S[2374], Cout[2374]);
	Full_Adder FA2323 (Cout[1713], Cout[1714], Cout[1715], S[2375], Cout[2375]);
	Full_Adder FA2324 (Cout[1716], Cout[1717], Cout[1718], S[2376], Cout[2376]);
	Full_Adder FA2325 (Cout[1719], S[1720], S[1721], S[2377], Cout[2377]);
	Full_Adder FA2326 (S[1722], S[1723], S[1724], S[2378], Cout[2378]);
	Full_Adder FA2327 (S[1725], S[1726], S[1727], S[2379], Cout[2379]);
	Full_Adder FA2328 (S[975], Cout[1720], Cout[1721], S[2380], Cout[2380]);
	Full_Adder FA2329 (Cout[1722], Cout[1723], Cout[1724], S[2381], Cout[2381]);
	Full_Adder FA2330 (Cout[1725], Cout[1726], Cout[1727], S[2382], Cout[2382]);
	Full_Adder FA2331 (Cout[1728], S[1729], S[1730], S[2383], Cout[2383]);
	Full_Adder FA2332 (S[1731], S[1732], S[1733], S[2384], Cout[2384]);
	Full_Adder FA2333 (S[1734], S[1735], S[1736], S[2385], Cout[2385]);
	Full_Adder FA2334 (S[989], Cout[1729], Cout[1730], S[2386], Cout[2386]);
	Full_Adder FA2335 (Cout[1731], Cout[1732], Cout[1733], S[2387], Cout[2387]);
	Full_Adder FA2336 (Cout[1734], Cout[1735], Cout[1736], S[2388], Cout[2388]);
	Full_Adder FA2337 (Cout[1737], S[1738], S[1739], S[2389], Cout[2389]);
	Full_Adder FA2338 (S[1740], S[1741], S[1742], S[2390], Cout[2390]);
	Full_Adder FA2339 (S[1743], S[1744], S[1745], S[2391], Cout[2391]);
	Full_Adder FA2340 (S[1003], Cout[1738], Cout[1739], S[2392], Cout[2392]);
	Full_Adder FA2341 (Cout[1740], Cout[1741], Cout[1742], S[2393], Cout[2393]);
	Full_Adder FA2342 (Cout[1743], Cout[1744], Cout[1745], S[2394], Cout[2394]);
	Full_Adder FA2343 (Cout[1746], S[1747], S[1748], S[2395], Cout[2395]);
	Full_Adder FA2344 (S[1749], S[1750], S[1751], S[2396], Cout[2396]);
	Full_Adder FA2345 (S[1752], S[1753], S[1754], S[2397], Cout[2397]);
	Full_Adder FA2346 (S[1017], Cout[1747], Cout[1748], S[2398], Cout[2398]);
	Full_Adder FA2347 (Cout[1749], Cout[1750], Cout[1751], S[2399], Cout[2399]);
	Full_Adder FA2348 (Cout[1752], Cout[1753], Cout[1754], S[2400], Cout[2400]);
	Full_Adder FA2349 (Cout[1755], S[1756], S[1757], S[2401], Cout[2401]);
	Full_Adder FA2350 (S[1758], S[1759], S[1760], S[2402], Cout[2402]);
	Full_Adder FA2351 (S[1761], S[1762], S[1763], S[2403], Cout[2403]);
	Full_Adder FA2352 (S[1031], Cout[1756], Cout[1757], S[2404], Cout[2404]);
	Full_Adder FA2353 (Cout[1758], Cout[1759], Cout[1760], S[2405], Cout[2405]);
	Full_Adder FA2354 (Cout[1761], Cout[1762], Cout[1763], S[2406], Cout[2406]);
	Full_Adder FA2355 (Cout[1764], S[1765], S[1766], S[2407], Cout[2407]);
	Full_Adder FA2356 (S[1767], S[1768], S[1769], S[2408], Cout[2408]);
	Full_Adder FA2357 (S[1770], S[1771], S[1772], S[2409], Cout[2409]);
	Full_Adder FA2358 (S[1045], Cout[1765], Cout[1766], S[2410], Cout[2410]);
	Full_Adder FA2359 (Cout[1767], Cout[1768], Cout[1769], S[2411], Cout[2411]);
	Full_Adder FA2360 (Cout[1770], Cout[1771], Cout[1772], S[2412], Cout[2412]);
	Full_Adder FA2361 (Cout[1773], S[1774], S[1775], S[2413], Cout[2413]);
	Full_Adder FA2362 (S[1776], S[1777], S[1778], S[2414], Cout[2414]);
	Full_Adder FA2363 (S[1779], S[1780], S[1781], S[2415], Cout[2415]);
	Full_Adder FA2364 (S[1059], Cout[1774], Cout[1775], S[2416], Cout[2416]);
	Full_Adder FA2365 (Cout[1776], Cout[1777], Cout[1778], S[2417], Cout[2417]);
	Full_Adder FA2366 (Cout[1779], Cout[1780], Cout[1781], S[2418], Cout[2418]);
	Full_Adder FA2367 (Cout[1782], S[1783], S[1784], S[2419], Cout[2419]);
	Full_Adder FA2368 (S[1785], S[1786], S[1787], S[2420], Cout[2420]);
	Full_Adder FA2369 (S[1788], S[1789], S[1790], S[2421], Cout[2421]);
	Full_Adder FA2370 (S[1073], Cout[1783], Cout[1784], S[2422], Cout[2422]);
	Full_Adder FA2371 (Cout[1785], Cout[1786], Cout[1787], S[2423], Cout[2423]);
	Full_Adder FA2372 (Cout[1788], Cout[1789], Cout[1790], S[2424], Cout[2424]);
	Full_Adder FA2373 (Cout[1791], S[1792], S[1793], S[2425], Cout[2425]);
	Full_Adder FA2374 (S[1794], S[1795], S[1796], S[2426], Cout[2426]);
	Full_Adder FA2375 (S[1797], S[1798], S[1799], S[2427], Cout[2427]);
	Full_Adder FA2376 (S[1087], Cout[1792], Cout[1793], S[2428], Cout[2428]);
	Full_Adder FA2377 (Cout[1794], Cout[1795], Cout[1796], S[2429], Cout[2429]);
	Full_Adder FA2378 (Cout[1797], Cout[1798], Cout[1799], S[2430], Cout[2430]);
	Full_Adder FA2379 (Cout[1800], S[1801], S[1802], S[2431], Cout[2431]);
	Full_Adder FA2380 (S[1803], S[1804], S[1805], S[2432], Cout[2432]);
	Full_Adder FA2381 (S[1806], S[1807], S[1808], S[2433], Cout[2433]);
	Full_Adder FA2382 (S[1101], Cout[1801], Cout[1802], S[2434], Cout[2434]);
	Full_Adder FA2383 (Cout[1803], Cout[1804], Cout[1805], S[2435], Cout[2435]);
	Full_Adder FA2384 (Cout[1806], Cout[1807], Cout[1808], S[2436], Cout[2436]);
	Full_Adder FA2385 (Cout[1809], S[1810], S[1811], S[2437], Cout[2437]);
	Full_Adder FA2386 (S[1812], S[1813], S[1814], S[2438], Cout[2438]);
	Full_Adder FA2387 (S[1815], S[1816], S[1817], S[2439], Cout[2439]);
	Full_Adder FA2388 (S[1115], Cout[1810], Cout[1811], S[2440], Cout[2440]);
	Full_Adder FA2389 (Cout[1812], Cout[1813], Cout[1814], S[2441], Cout[2441]);
	Full_Adder FA2390 (Cout[1815], Cout[1816], Cout[1817], S[2442], Cout[2442]);
	Full_Adder FA2391 (Cout[1818], S[1819], S[1820], S[2443], Cout[2443]);
	Full_Adder FA2392 (S[1821], S[1822], S[1823], S[2444], Cout[2444]);
	Full_Adder FA2393 (S[1824], S[1825], S[1826], S[2445], Cout[2445]);
	Full_Adder FA2394 (S[1129], Cout[1819], Cout[1820], S[2446], Cout[2446]);
	Full_Adder FA2395 (Cout[1821], Cout[1822], Cout[1823], S[2447], Cout[2447]);
	Full_Adder FA2396 (Cout[1824], Cout[1825], Cout[1826], S[2448], Cout[2448]);
	Full_Adder FA2397 (Cout[1827], S[1828], S[1829], S[2449], Cout[2449]);
	Full_Adder FA2398 (S[1830], S[1831], S[1832], S[2450], Cout[2450]);
	Full_Adder FA2399 (S[1833], S[1834], S[1835], S[2451], Cout[2451]);
	Full_Adder FA2400 (S[1143], Cout[1828], Cout[1829], S[2452], Cout[2452]);
	Full_Adder FA2401 (Cout[1830], Cout[1831], Cout[1832], S[2453], Cout[2453]);
	Full_Adder FA2402 (Cout[1833], Cout[1834], Cout[1835], S[2454], Cout[2454]);
	Full_Adder FA2403 (Cout[1836], S[1837], S[1838], S[2455], Cout[2455]);
	Full_Adder FA2404 (S[1839], S[1840], S[1841], S[2456], Cout[2456]);
	Full_Adder FA2405 (S[1842], S[1843], S[1844], S[2457], Cout[2457]);
	Full_Adder FA2406 (S[1157], Cout[1837], Cout[1838], S[2458], Cout[2458]);
	Full_Adder FA2407 (Cout[1839], Cout[1840], Cout[1841], S[2459], Cout[2459]);
	Full_Adder FA2408 (Cout[1842], Cout[1843], Cout[1844], S[2460], Cout[2460]);
	Full_Adder FA2409 (Cout[1845], S[1846], S[1847], S[2461], Cout[2461]);
	Full_Adder FA2410 (S[1848], S[1849], S[1850], S[2462], Cout[2462]);
	Full_Adder FA2411 (S[1851], S[1852], S[1853], S[2463], Cout[2463]);
	Full_Adder FA2412 (S[1171], Cout[1846], Cout[1847], S[2464], Cout[2464]);
	Full_Adder FA2413 (Cout[1848], Cout[1849], Cout[1850], S[2465], Cout[2465]);
	Full_Adder FA2414 (Cout[1851], Cout[1852], Cout[1853], S[2466], Cout[2466]);
	Full_Adder FA2415 (Cout[1854], S[1855], S[1856], S[2467], Cout[2467]);
	Full_Adder FA2416 (S[1857], S[1858], S[1859], S[2468], Cout[2468]);
	Full_Adder FA2417 (S[1860], S[1861], S[1862], S[2469], Cout[2469]);
	Full_Adder FA2418 (S[1185], Cout[1855], Cout[1856], S[2470], Cout[2470]);
	Full_Adder FA2419 (Cout[1857], Cout[1858], Cout[1859], S[2471], Cout[2471]);
	Full_Adder FA2420 (Cout[1860], Cout[1861], Cout[1862], S[2472], Cout[2472]);
	Full_Adder FA2421 (Cout[1863], S[1864], S[1865], S[2473], Cout[2473]);
	Full_Adder FA2422 (S[1866], S[1867], S[1868], S[2474], Cout[2474]);
	Full_Adder FA2423 (S[1869], S[1870], S[1871], S[2475], Cout[2475]);
	Full_Adder FA2424 (S[1199], Cout[1864], Cout[1865], S[2476], Cout[2476]);
	Full_Adder FA2425 (Cout[1866], Cout[1867], Cout[1868], S[2477], Cout[2477]);
	Full_Adder FA2426 (Cout[1869], Cout[1870], Cout[1871], S[2478], Cout[2478]);
	Full_Adder FA2427 (Cout[1872], S[1873], S[1874], S[2479], Cout[2479]);
	Full_Adder FA2428 (S[1875], S[1876], S[1877], S[2480], Cout[2480]);
	Full_Adder FA2429 (S[1878], S[1879], S[1880], S[2481], Cout[2481]);
	Full_Adder FA2430 (S[1213], Cout[1873], Cout[1874], S[2482], Cout[2482]);
	Full_Adder FA2431 (Cout[1875], Cout[1876], Cout[1877], S[2483], Cout[2483]);
	Full_Adder FA2432 (Cout[1878], Cout[1879], Cout[1880], S[2484], Cout[2484]);
	Full_Adder FA2433 (Cout[1881], S[1882], S[1883], S[2485], Cout[2485]);
	Full_Adder FA2434 (S[1884], S[1885], S[1886], S[2486], Cout[2486]);
	Full_Adder FA2435 (S[1887], S[1888], S[1889], S[2487], Cout[2487]);
	Full_Adder FA2436 (S[1227], Cout[1882], Cout[1883], S[2488], Cout[2488]);
	Full_Adder FA2437 (Cout[1884], Cout[1885], Cout[1886], S[2489], Cout[2489]);
	Full_Adder FA2438 (Cout[1887], Cout[1888], Cout[1889], S[2490], Cout[2490]);
	Full_Adder FA2439 (Cout[1890], S[1891], S[1892], S[2491], Cout[2491]);
	Full_Adder FA2440 (S[1893], S[1894], S[1895], S[2492], Cout[2492]);
	Full_Adder FA2441 (S[1896], S[1897], S[1898], S[2493], Cout[2493]);
	Full_Adder FA2442 (S[1241], Cout[1891], Cout[1892], S[2494], Cout[2494]);
	Full_Adder FA2443 (Cout[1893], Cout[1894], Cout[1895], S[2495], Cout[2495]);
	Full_Adder FA2444 (Cout[1896], Cout[1897], Cout[1898], S[2496], Cout[2496]);
	Full_Adder FA2445 (Cout[1899], S[1900], S[1901], S[2497], Cout[2497]);
	Full_Adder FA2446 (S[1902], S[1903], S[1904], S[2498], Cout[2498]);
	Full_Adder FA2447 (S[1905], S[1906], S[1907], S[2499], Cout[2499]);
	Full_Adder FA2448 (S[1254], Cout[1900], Cout[1901], S[2500], Cout[2500]);
	Full_Adder FA2449 (Cout[1902], Cout[1903], Cout[1904], S[2501], Cout[2501]);
	Full_Adder FA2450 (Cout[1905], Cout[1906], Cout[1907], S[2502], Cout[2502]);
	Full_Adder FA2451 (Cout[1908], S[1909], S[1910], S[2503], Cout[2503]);
	Full_Adder FA2452 (S[1911], S[1912], S[1913], S[2504], Cout[2504]);
	Full_Adder FA2453 (S[1914], S[1915], S[1916], S[2505], Cout[2505]);
	Full_Adder FA2454 (S[1266], Cout[1909], Cout[1910], S[2506], Cout[2506]);
	Full_Adder FA2455 (Cout[1911], Cout[1912], Cout[1913], S[2507], Cout[2507]);
	Full_Adder FA2456 (Cout[1914], Cout[1915], Cout[1916], S[2508], Cout[2508]);
	Full_Adder FA2457 (Cout[1917], S[1918], S[1919], S[2509], Cout[2509]);
	Full_Adder FA2458 (S[1920], S[1921], S[1922], S[2510], Cout[2510]);
	Full_Adder FA2459 (S[1923], S[1924], S[1925], S[2511], Cout[2511]);
	Full_Adder FA2460 (S[1277], Cout[1918], Cout[1919], S[2512], Cout[2512]);
	Full_Adder FA2461 (Cout[1920], Cout[1921], Cout[1922], S[2513], Cout[2513]);
	Full_Adder FA2462 (Cout[1923], Cout[1924], Cout[1925], S[2514], Cout[2514]);
	Full_Adder FA2463 (Cout[1926], S[1927], S[1928], S[2515], Cout[2515]);
	Full_Adder FA2464 (S[1929], S[1930], S[1931], S[2516], Cout[2516]);
	Full_Adder FA2465 (S[1932], S[1933], S[1934], S[2517], Cout[2517]);
	Full_Adder FA2466 (S[1287], Cout[1927], Cout[1928], S[2518], Cout[2518]);
	Full_Adder FA2467 (Cout[1929], Cout[1930], Cout[1931], S[2519], Cout[2519]);
	Full_Adder FA2468 (Cout[1932], Cout[1933], Cout[1934], S[2520], Cout[2520]);
	Full_Adder FA2469 (Cout[1935], S[1936], S[1937], S[2521], Cout[2521]);
	Full_Adder FA2470 (S[1938], S[1939], S[1940], S[2522], Cout[2522]);
	Full_Adder FA2471 (S[1941], S[1942], S[1943], S[2523], Cout[2523]);
	Full_Adder FA2472 (S[1296], Cout[1936], Cout[1937], S[2524], Cout[2524]);
	Full_Adder FA2473 (Cout[1938], Cout[1939], Cout[1940], S[2525], Cout[2525]);
	Full_Adder FA2474 (Cout[1941], Cout[1942], Cout[1943], S[2526], Cout[2526]);
	Full_Adder FA2475 (Cout[1944], S[1945], S[1946], S[2527], Cout[2527]);
	Full_Adder FA2476 (S[1947], S[1948], S[1949], S[2528], Cout[2528]);
	Full_Adder FA2477 (S[1950], S[1951], S[1952], S[2529], Cout[2529]);
	Full_Adder FA2478 (S[1304], Cout[1945], Cout[1946], S[2530], Cout[2530]);
	Full_Adder FA2479 (Cout[1947], Cout[1948], Cout[1949], S[2531], Cout[2531]);
	Full_Adder FA2480 (Cout[1950], Cout[1951], Cout[1952], S[2532], Cout[2532]);
	Full_Adder FA2481 (Cout[1953], S[1954], S[1955], S[2533], Cout[2533]);
	Full_Adder FA2482 (S[1956], S[1957], S[1958], S[2534], Cout[2534]);
	Full_Adder FA2483 (S[1959], S[1960], S[1961], S[2535], Cout[2535]);
	Full_Adder FA2484 (S[1311], Cout[1954], Cout[1955], S[2536], Cout[2536]);
	Full_Adder FA2485 (Cout[1956], Cout[1957], Cout[1958], S[2537], Cout[2537]);
	Full_Adder FA2486 (Cout[1959], Cout[1960], Cout[1961], S[2538], Cout[2538]);
	Full_Adder FA2487 (Cout[1962], S[1963], S[1964], S[2539], Cout[2539]);
	Full_Adder FA2488 (S[1965], S[1966], S[1967], S[2540], Cout[2540]);
	Full_Adder FA2489 (S[1968], S[1969], S[1970], S[2541], Cout[2541]);
	Full_Adder FA2490 (S[1317], Cout[1963], Cout[1964], S[2542], Cout[2542]);
	Full_Adder FA2491 (Cout[1965], Cout[1966], Cout[1967], S[2543], Cout[2543]);
	Full_Adder FA2492 (Cout[1968], Cout[1969], Cout[1970], S[2544], Cout[2544]);
	Full_Adder FA2493 (Cout[1971], S[1972], S[1973], S[2545], Cout[2545]);
	Full_Adder FA2494 (S[1974], S[1975], S[1976], S[2546], Cout[2546]);
	Full_Adder FA2495 (S[1977], S[1978], S[1979], S[2547], Cout[2547]);
	Full_Adder FA2496 (S[1322], Cout[1972], Cout[1973], S[2548], Cout[2548]);
	Full_Adder FA2497 (Cout[1974], Cout[1975], Cout[1976], S[2549], Cout[2549]);
	Full_Adder FA2498 (Cout[1977], Cout[1978], Cout[1979], S[2550], Cout[2550]);
	Full_Adder FA2499 (Cout[1980], S[1981], S[1982], S[2551], Cout[2551]);
	Full_Adder FA2500 (S[1983], S[1984], S[1985], S[2552], Cout[2552]);
	Full_Adder FA2501 (S[1986], S[1987], S[1988], S[2553], Cout[2553]);
	Full_Adder FA2502 (S[1326], Cout[1981], Cout[1982], S[2554], Cout[2554]);
	Full_Adder FA2503 (Cout[1983], Cout[1984], Cout[1985], S[2555], Cout[2555]);
	Full_Adder FA2504 (Cout[1986], Cout[1987], Cout[1988], S[2556], Cout[2556]);
	Full_Adder FA2505 (Cout[1989], S[1990], S[1991], S[2557], Cout[2557]);
	Full_Adder FA2506 (S[1992], S[1993], S[1994], S[2558], Cout[2558]);
	Full_Adder FA2507 (S[1995], S[1996], S[1997], S[2559], Cout[2559]);
	Full_Adder FA2508 (S[1329], Cout[1990], Cout[1991], S[2560], Cout[2560]);
	Full_Adder FA2509 (Cout[1992], Cout[1993], Cout[1994], S[2561], Cout[2561]);
	Full_Adder FA2510 (Cout[1995], Cout[1996], Cout[1997], S[2562], Cout[2562]);
	Full_Adder FA2511 (Cout[1998], S[1999], S[2000], S[2563], Cout[2563]);
	Full_Adder FA2512 (S[2001], S[2002], S[2003], S[2564], Cout[2564]);
	Full_Adder FA2513 (S[2004], S[2005], S[2006], S[2565], Cout[2565]);
	Full_Adder FA2514 (S[1331], Cout[1999], Cout[2000], S[2566], Cout[2566]);
	Full_Adder FA2515 (Cout[2001], Cout[2002], Cout[2003], S[2567], Cout[2567]);
	Full_Adder FA2516 (Cout[2004], Cout[2005], Cout[2006], S[2568], Cout[2568]);
	Full_Adder FA2517 (Cout[2007], S[2008], S[2009], S[2569], Cout[2569]);
	Full_Adder FA2518 (S[2010], S[2011], S[2012], S[2570], Cout[2570]);
	Full_Adder FA2519 (S[2013], S[2014], S[2015], S[2571], Cout[2571]);
	Full_Adder FA2520 (S[1332], Cout[2008], Cout[2009], S[2572], Cout[2572]);
	Full_Adder FA2521 (Cout[2010], Cout[2011], Cout[2012], S[2573], Cout[2573]);
	Full_Adder FA2522 (Cout[2013], Cout[2014], Cout[2015], S[2574], Cout[2574]);
	Full_Adder FA2523 (Cout[2016], S[2017], S[2018], S[2575], Cout[2575]);
	Full_Adder FA2524 (S[2019], S[2020], S[2021], S[2576], Cout[2576]);
	Full_Adder FA2525 (S[2022], S[2023], S[2024], S[2577], Cout[2577]);
	Full_Adder FA2526 (Cout[1332], Cout[2017], Cout[2018], S[2578], Cout[2578]);
	Full_Adder FA2527 (Cout[2019], Cout[2020], Cout[2021], S[2579], Cout[2579]);
	Full_Adder FA2528 (Cout[2022], Cout[2023], Cout[2024], S[2580], Cout[2580]);
	Full_Adder FA2529 (Cout[2025], S[2026], S[2027], S[2581], Cout[2581]);
	Full_Adder FA2530 (S[2028], S[2029], S[2030], S[2582], Cout[2582]);
	Full_Adder FA2531 (S[2031], S[2032], S[2033], S[2583], Cout[2583]);
	Full_Adder FA2532 (pp62[39], pp63[38], Cout[2026], S[2584], Cout[2584]);
	Full_Adder FA2533 (Cout[2027], Cout[2028], Cout[2029], S[2585], Cout[2585]);
	Full_Adder FA2534 (Cout[2030], Cout[2031], Cout[2032], S[2586], Cout[2586]);
	Full_Adder FA2535 (Cout[2033], Cout[2034], S[2035], S[2587], Cout[2587]);
	Full_Adder FA2536 (S[2036], S[2037], S[2038], S[2588], Cout[2588]);
	Full_Adder FA2537 (S[2039], S[2040], S[2041], S[2589], Cout[2589]);
	Full_Adder FA2538 (pp60[42], pp61[41], pp62[40], S[2590], Cout[2590]);
	Full_Adder FA2539 (pp63[39], Cout[2035], Cout[2036], S[2591], Cout[2591]);
	Full_Adder FA2540 (Cout[2037], Cout[2038], Cout[2039], S[2592], Cout[2592]);
	Full_Adder FA2541 (Cout[2040], Cout[2041], Cout[2042], S[2593], Cout[2593]);
	Full_Adder FA2542 (S[2043], S[2044], S[2045], S[2594], Cout[2594]);
	Full_Adder FA2543 (S[2046], S[2047], S[2048], S[2595], Cout[2595]);
	Full_Adder FA2544 (pp58[45], pp59[44], pp60[43], S[2596], Cout[2596]);
	Full_Adder FA2545 (pp61[42], pp62[41], pp63[40], S[2597], Cout[2597]);
	Full_Adder FA2546 (Cout[2043], Cout[2044], Cout[2045], S[2598], Cout[2598]);
	Full_Adder FA2547 (Cout[2046], Cout[2047], Cout[2048], S[2599], Cout[2599]);
	Full_Adder FA2548 (Cout[2049], S[2050], S[2051], S[2600], Cout[2600]);
	Full_Adder FA2549 (S[2052], S[2053], S[2054], S[2601], Cout[2601]);
	Full_Adder FA2550 (pp56[48], pp57[47], pp58[46], S[2602], Cout[2602]);
	Full_Adder FA2551 (pp59[45], pp60[44], pp61[43], S[2603], Cout[2603]);
	Full_Adder FA2552 (pp62[42], pp63[41], Cout[2050], S[2604], Cout[2604]);
	Full_Adder FA2553 (Cout[2051], Cout[2052], Cout[2053], S[2605], Cout[2605]);
	Full_Adder FA2554 (Cout[2054], Cout[2055], S[2056], S[2606], Cout[2606]);
	Full_Adder FA2555 (S[2057], S[2058], S[2059], S[2607], Cout[2607]);
	Full_Adder FA2556 (pp54[51], pp55[50], pp56[49], S[2608], Cout[2608]);
	Full_Adder FA2557 (pp57[48], pp58[47], pp59[46], S[2609], Cout[2609]);
	Full_Adder FA2558 (pp60[45], pp61[44], pp62[43], S[2610], Cout[2610]);
	Full_Adder FA2559 (pp63[42], Cout[2056], Cout[2057], S[2611], Cout[2611]);
	Full_Adder FA2560 (Cout[2058], Cout[2059], Cout[2060], S[2612], Cout[2612]);
	Full_Adder FA2561 (S[2061], S[2062], S[2063], S[2613], Cout[2613]);
	Full_Adder FA2562 (pp52[54], pp53[53], pp54[52], S[2614], Cout[2614]);
	Full_Adder FA2563 (pp55[51], pp56[50], pp57[49], S[2615], Cout[2615]);
	Full_Adder FA2564 (pp58[48], pp59[47], pp60[46], S[2616], Cout[2616]);
	Full_Adder FA2565 (pp61[45], pp62[44], pp63[43], S[2617], Cout[2617]);
	Full_Adder FA2566 (Cout[2061], Cout[2062], Cout[2063], S[2618], Cout[2618]);
	Full_Adder FA2567 (Cout[2064], S[2065], S[2066], S[2619], Cout[2619]);
	Full_Adder FA2568 (pp50[57], pp51[56], pp52[55], S[2620], Cout[2620]);
	Full_Adder FA2569 (pp53[54], pp54[53], pp55[52], S[2621], Cout[2621]);
	Full_Adder FA2570 (pp56[51], pp57[50], pp58[49], S[2622], Cout[2622]);
	Full_Adder FA2571 (pp59[48], pp60[47], pp61[46], S[2623], Cout[2623]);
	Full_Adder FA2572 (pp62[45], pp63[44], Cout[2065], S[2624], Cout[2624]);
	Full_Adder FA2573 (Cout[2066], Cout[2067], S[2068], S[2625], Cout[2625]);
	Full_Adder FA2574 (pp48[60], pp49[59], pp50[58], S[2626], Cout[2626]);
	Full_Adder FA2575 (pp51[57], pp52[56], pp53[55], S[2627], Cout[2627]);
	Full_Adder FA2576 (pp54[54], pp55[53], pp56[52], S[2628], Cout[2628]);
	Full_Adder FA2577 (pp57[51], pp58[50], pp59[49], S[2629], Cout[2629]);
	Full_Adder FA2578 (pp60[48], pp61[47], pp62[46], S[2630], Cout[2630]);
	Full_Adder FA2579 (pp63[45], Cout[2068], Cout[2069], S[2631], Cout[2631]);
	Full_Adder FA2580 (pp46[63], pp47[62], pp48[61], S[2632], Cout[2632]);
	Full_Adder FA2581 (pp49[60], pp50[59], pp51[58], S[2633], Cout[2633]);
	Full_Adder FA2582 (pp52[57], pp53[56], pp54[55], S[2634], Cout[2634]);
	Full_Adder FA2583 (pp55[54], pp56[53], pp57[52], S[2635], Cout[2635]);
	Full_Adder FA2584 (pp58[51], pp59[50], pp60[49], S[2636], Cout[2636]);
	Full_Adder FA2585 (pp61[48], pp62[47], pp63[46], S[2637], Cout[2637]);
	Full_Adder FA2586 (pp47[63], pp48[62], pp49[61], S[2638], Cout[2638]);
	Full_Adder FA2587 (pp50[60], pp51[59], pp52[58], S[2639], Cout[2639]);
	Full_Adder FA2588 (pp53[57], pp54[56], pp55[55], S[2640], Cout[2640]);
	Full_Adder FA2589 (pp56[54], pp57[53], pp58[52], S[2641], Cout[2641]);
	Full_Adder FA2590 (pp59[51], pp60[50], pp61[49], S[2642], Cout[2642]);
	Full_Adder FA2591 (pp48[63], pp49[62], pp50[61], S[2643], Cout[2643]);
	Full_Adder FA2592 (pp51[60], pp52[59], pp53[58], S[2644], Cout[2644]);
	Full_Adder FA2593 (pp54[57], pp55[56], pp56[55], S[2645], Cout[2645]);
	Full_Adder FA2594 (pp57[54], pp58[53], pp59[52], S[2646], Cout[2646]);
	Full_Adder FA2595 (pp49[63], pp50[62], pp51[61], S[2647], Cout[2647]);
	Full_Adder FA2596 (pp52[60], pp53[59], pp54[58], S[2648], Cout[2648]);
	Full_Adder FA2597 (pp55[57], pp56[56], pp57[55], S[2649], Cout[2649]);
	Full_Adder FA2598 (pp50[63], pp51[62], pp52[61], S[2650], Cout[2650]);
	Full_Adder FA2599 (pp53[60], pp54[59], pp55[58], S[2651], Cout[2651]);
	Full_Adder FA2600 (pp51[63], pp52[62], pp53[61], S[2652], Cout[2652]);
	Half_Adder HA53 (pp0[9], pp1[8], S[2653], Cout[2653]);
	Full_Adder FA2601 (pp0[10], pp1[9], pp2[8], S[2654], Cout[2654]);
	Half_Adder HA54 (pp3[7], pp4[6], S[2655], Cout[2655]);
	Full_Adder FA2602 (pp0[11], pp1[10], pp2[9], S[2656], Cout[2656]);
	Full_Adder FA2603 (pp3[8], pp4[7], pp5[6], S[2657], Cout[2657]);
	Half_Adder HA55 (pp6[5], pp7[4], S[2658], Cout[2658]);
	Full_Adder FA2604 (pp0[12], pp1[11], pp2[10], S[2659], Cout[2659]);
	Full_Adder FA2605 (pp3[9], pp4[8], pp5[7], S[2660], Cout[2660]);
	Full_Adder FA2606 (pp6[6], pp7[5], pp8[4], S[2661], Cout[2661]);
	Half_Adder HA56 (pp9[3], pp10[2], S[2662], Cout[2662]);
	Full_Adder FA2607 (pp2[11], pp3[10], pp4[9], S[2663], Cout[2663]);
	Full_Adder FA2608 (pp5[8], pp6[7], pp7[6], S[2664], Cout[2664]);
	Full_Adder FA2609 (pp8[5], pp9[4], pp10[3], S[2665], Cout[2665]);
	Full_Adder FA2610 (pp11[2], pp12[1], pp13[0], S[2666], Cout[2666]);
	Full_Adder FA2611 (pp5[9], pp6[8], pp7[7], S[2667], Cout[2667]);
	Full_Adder FA2612 (pp8[6], pp9[5], pp10[4], S[2668], Cout[2668]);
	Full_Adder FA2613 (pp11[3], pp12[2], pp13[1], S[2669], Cout[2669]);
	Full_Adder FA2614 (pp14[0], Cout[2071], S[2072], S[2670], Cout[2670]);
	Full_Adder FA2615 (pp8[7], pp9[6], pp10[5], S[2671], Cout[2671]);
	Full_Adder FA2616 (pp11[4], pp12[3], pp13[2], S[2672], Cout[2672]);
	Full_Adder FA2617 (pp14[1], pp15[0], Cout[2072], S[2673], Cout[2673]);
	Full_Adder FA2618 (Cout[2073], S[2074], S[2075], S[2674], Cout[2674]);
	Full_Adder FA2619 (pp11[5], pp12[4], pp13[3], S[2675], Cout[2675]);
	Full_Adder FA2620 (pp14[2], pp15[1], pp16[0], S[2676], Cout[2676]);
	Full_Adder FA2621 (Cout[2074], Cout[2075], Cout[2076], S[2677], Cout[2677]);
	Full_Adder FA2622 (S[2077], S[2078], S[2079], S[2678], Cout[2678]);
	Full_Adder FA2623 (pp14[3], pp15[2], pp16[1], S[2679], Cout[2679]);
	Full_Adder FA2624 (pp17[0], Cout[2077], Cout[2078], S[2680], Cout[2680]);
	Full_Adder FA2625 (Cout[2079], Cout[2080], S[2081], S[2681], Cout[2681]);
	Full_Adder FA2626 (S[2082], S[2083], S[2084], S[2682], Cout[2682]);
	Full_Adder FA2627 (pp17[1], pp18[0], Cout[2081], S[2683], Cout[2683]);
	Full_Adder FA2628 (Cout[2082], Cout[2083], Cout[2084], S[2684], Cout[2684]);
	Full_Adder FA2629 (Cout[2085], S[2086], S[2087], S[2685], Cout[2685]);
	Full_Adder FA2630 (S[2088], S[2089], S[2090], S[2686], Cout[2686]);
	Full_Adder FA2631 (S[1333], Cout[2086], Cout[2087], S[2687], Cout[2687]);
	Full_Adder FA2632 (Cout[2088], Cout[2089], Cout[2090], S[2688], Cout[2688]);
	Full_Adder FA2633 (Cout[2091], S[2092], S[2093], S[2689], Cout[2689]);
	Full_Adder FA2634 (S[2094], S[2095], S[2096], S[2690], Cout[2690]);
	Full_Adder FA2635 (S[1335], Cout[2092], Cout[2093], S[2691], Cout[2691]);
	Full_Adder FA2636 (Cout[2094], Cout[2095], Cout[2096], S[2692], Cout[2692]);
	Full_Adder FA2637 (Cout[2097], S[2098], S[2099], S[2693], Cout[2693]);
	Full_Adder FA2638 (S[2100], S[2101], S[2102], S[2694], Cout[2694]);
	Full_Adder FA2639 (S[1338], Cout[2098], Cout[2099], S[2695], Cout[2695]);
	Full_Adder FA2640 (Cout[2100], Cout[2101], Cout[2102], S[2696], Cout[2696]);
	Full_Adder FA2641 (Cout[2103], S[2104], S[2105], S[2697], Cout[2697]);
	Full_Adder FA2642 (S[2106], S[2107], S[2108], S[2698], Cout[2698]);
	Full_Adder FA2643 (S[1342], Cout[2104], Cout[2105], S[2699], Cout[2699]);
	Full_Adder FA2644 (Cout[2106], Cout[2107], Cout[2108], S[2700], Cout[2700]);
	Full_Adder FA2645 (Cout[2109], S[2110], S[2111], S[2701], Cout[2701]);
	Full_Adder FA2646 (S[2112], S[2113], S[2114], S[2702], Cout[2702]);
	Full_Adder FA2647 (S[1347], Cout[2110], Cout[2111], S[2703], Cout[2703]);
	Full_Adder FA2648 (Cout[2112], Cout[2113], Cout[2114], S[2704], Cout[2704]);
	Full_Adder FA2649 (Cout[2115], S[2116], S[2117], S[2705], Cout[2705]);
	Full_Adder FA2650 (S[2118], S[2119], S[2120], S[2706], Cout[2706]);
	Full_Adder FA2651 (S[1353], Cout[2116], Cout[2117], S[2707], Cout[2707]);
	Full_Adder FA2652 (Cout[2118], Cout[2119], Cout[2120], S[2708], Cout[2708]);
	Full_Adder FA2653 (Cout[2121], S[2122], S[2123], S[2709], Cout[2709]);
	Full_Adder FA2654 (S[2124], S[2125], S[2126], S[2710], Cout[2710]);
	Full_Adder FA2655 (S[1360], Cout[2122], Cout[2123], S[2711], Cout[2711]);
	Full_Adder FA2656 (Cout[2124], Cout[2125], Cout[2126], S[2712], Cout[2712]);
	Full_Adder FA2657 (Cout[2127], S[2128], S[2129], S[2713], Cout[2713]);
	Full_Adder FA2658 (S[2130], S[2131], S[2132], S[2714], Cout[2714]);
	Full_Adder FA2659 (S[1368], Cout[2128], Cout[2129], S[2715], Cout[2715]);
	Full_Adder FA2660 (Cout[2130], Cout[2131], Cout[2132], S[2716], Cout[2716]);
	Full_Adder FA2661 (Cout[2133], S[2134], S[2135], S[2717], Cout[2717]);
	Full_Adder FA2662 (S[2136], S[2137], S[2138], S[2718], Cout[2718]);
	Full_Adder FA2663 (S[1377], Cout[2134], Cout[2135], S[2719], Cout[2719]);
	Full_Adder FA2664 (Cout[2136], Cout[2137], Cout[2138], S[2720], Cout[2720]);
	Full_Adder FA2665 (Cout[2139], S[2140], S[2141], S[2721], Cout[2721]);
	Full_Adder FA2666 (S[2142], S[2143], S[2144], S[2722], Cout[2722]);
	Full_Adder FA2667 (S[1386], Cout[2140], Cout[2141], S[2723], Cout[2723]);
	Full_Adder FA2668 (Cout[2142], Cout[2143], Cout[2144], S[2724], Cout[2724]);
	Full_Adder FA2669 (Cout[2145], S[2146], S[2147], S[2725], Cout[2725]);
	Full_Adder FA2670 (S[2148], S[2149], S[2150], S[2726], Cout[2726]);
	Full_Adder FA2671 (S[1395], Cout[2146], Cout[2147], S[2727], Cout[2727]);
	Full_Adder FA2672 (Cout[2148], Cout[2149], Cout[2150], S[2728], Cout[2728]);
	Full_Adder FA2673 (Cout[2151], S[2152], S[2153], S[2729], Cout[2729]);
	Full_Adder FA2674 (S[2154], S[2155], S[2156], S[2730], Cout[2730]);
	Full_Adder FA2675 (S[1404], Cout[2152], Cout[2153], S[2731], Cout[2731]);
	Full_Adder FA2676 (Cout[2154], Cout[2155], Cout[2156], S[2732], Cout[2732]);
	Full_Adder FA2677 (Cout[2157], S[2158], S[2159], S[2733], Cout[2733]);
	Full_Adder FA2678 (S[2160], S[2161], S[2162], S[2734], Cout[2734]);
	Full_Adder FA2679 (S[1413], Cout[2158], Cout[2159], S[2735], Cout[2735]);
	Full_Adder FA2680 (Cout[2160], Cout[2161], Cout[2162], S[2736], Cout[2736]);
	Full_Adder FA2681 (Cout[2163], S[2164], S[2165], S[2737], Cout[2737]);
	Full_Adder FA2682 (S[2166], S[2167], S[2168], S[2738], Cout[2738]);
	Full_Adder FA2683 (S[1422], Cout[2164], Cout[2165], S[2739], Cout[2739]);
	Full_Adder FA2684 (Cout[2166], Cout[2167], Cout[2168], S[2740], Cout[2740]);
	Full_Adder FA2685 (Cout[2169], S[2170], S[2171], S[2741], Cout[2741]);
	Full_Adder FA2686 (S[2172], S[2173], S[2174], S[2742], Cout[2742]);
	Full_Adder FA2687 (S[1431], Cout[2170], Cout[2171], S[2743], Cout[2743]);
	Full_Adder FA2688 (Cout[2172], Cout[2173], Cout[2174], S[2744], Cout[2744]);
	Full_Adder FA2689 (Cout[2175], S[2176], S[2177], S[2745], Cout[2745]);
	Full_Adder FA2690 (S[2178], S[2179], S[2180], S[2746], Cout[2746]);
	Full_Adder FA2691 (S[1440], Cout[2176], Cout[2177], S[2747], Cout[2747]);
	Full_Adder FA2692 (Cout[2178], Cout[2179], Cout[2180], S[2748], Cout[2748]);
	Full_Adder FA2693 (Cout[2181], S[2182], S[2183], S[2749], Cout[2749]);
	Full_Adder FA2694 (S[2184], S[2185], S[2186], S[2750], Cout[2750]);
	Full_Adder FA2695 (S[1449], Cout[2182], Cout[2183], S[2751], Cout[2751]);
	Full_Adder FA2696 (Cout[2184], Cout[2185], Cout[2186], S[2752], Cout[2752]);
	Full_Adder FA2697 (Cout[2187], S[2188], S[2189], S[2753], Cout[2753]);
	Full_Adder FA2698 (S[2190], S[2191], S[2192], S[2754], Cout[2754]);
	Full_Adder FA2699 (S[1458], Cout[2188], Cout[2189], S[2755], Cout[2755]);
	Full_Adder FA2700 (Cout[2190], Cout[2191], Cout[2192], S[2756], Cout[2756]);
	Full_Adder FA2701 (Cout[2193], S[2194], S[2195], S[2757], Cout[2757]);
	Full_Adder FA2702 (S[2196], S[2197], S[2198], S[2758], Cout[2758]);
	Full_Adder FA2703 (S[1467], Cout[2194], Cout[2195], S[2759], Cout[2759]);
	Full_Adder FA2704 (Cout[2196], Cout[2197], Cout[2198], S[2760], Cout[2760]);
	Full_Adder FA2705 (Cout[2199], S[2200], S[2201], S[2761], Cout[2761]);
	Full_Adder FA2706 (S[2202], S[2203], S[2204], S[2762], Cout[2762]);
	Full_Adder FA2707 (S[1476], Cout[2200], Cout[2201], S[2763], Cout[2763]);
	Full_Adder FA2708 (Cout[2202], Cout[2203], Cout[2204], S[2764], Cout[2764]);
	Full_Adder FA2709 (Cout[2205], S[2206], S[2207], S[2765], Cout[2765]);
	Full_Adder FA2710 (S[2208], S[2209], S[2210], S[2766], Cout[2766]);
	Full_Adder FA2711 (S[1485], Cout[2206], Cout[2207], S[2767], Cout[2767]);
	Full_Adder FA2712 (Cout[2208], Cout[2209], Cout[2210], S[2768], Cout[2768]);
	Full_Adder FA2713 (Cout[2211], S[2212], S[2213], S[2769], Cout[2769]);
	Full_Adder FA2714 (S[2214], S[2215], S[2216], S[2770], Cout[2770]);
	Full_Adder FA2715 (S[1494], Cout[2212], Cout[2213], S[2771], Cout[2771]);
	Full_Adder FA2716 (Cout[2214], Cout[2215], Cout[2216], S[2772], Cout[2772]);
	Full_Adder FA2717 (Cout[2217], S[2218], S[2219], S[2773], Cout[2773]);
	Full_Adder FA2718 (S[2220], S[2221], S[2222], S[2774], Cout[2774]);
	Full_Adder FA2719 (S[1503], Cout[2218], Cout[2219], S[2775], Cout[2775]);
	Full_Adder FA2720 (Cout[2220], Cout[2221], Cout[2222], S[2776], Cout[2776]);
	Full_Adder FA2721 (Cout[2223], S[2224], S[2225], S[2777], Cout[2777]);
	Full_Adder FA2722 (S[2226], S[2227], S[2228], S[2778], Cout[2778]);
	Full_Adder FA2723 (S[1512], Cout[2224], Cout[2225], S[2779], Cout[2779]);
	Full_Adder FA2724 (Cout[2226], Cout[2227], Cout[2228], S[2780], Cout[2780]);
	Full_Adder FA2725 (Cout[2229], S[2230], S[2231], S[2781], Cout[2781]);
	Full_Adder FA2726 (S[2232], S[2233], S[2234], S[2782], Cout[2782]);
	Full_Adder FA2727 (S[1521], Cout[2230], Cout[2231], S[2783], Cout[2783]);
	Full_Adder FA2728 (Cout[2232], Cout[2233], Cout[2234], S[2784], Cout[2784]);
	Full_Adder FA2729 (Cout[2235], S[2236], S[2237], S[2785], Cout[2785]);
	Full_Adder FA2730 (S[2238], S[2239], S[2240], S[2786], Cout[2786]);
	Full_Adder FA2731 (S[1530], Cout[2236], Cout[2237], S[2787], Cout[2787]);
	Full_Adder FA2732 (Cout[2238], Cout[2239], Cout[2240], S[2788], Cout[2788]);
	Full_Adder FA2733 (Cout[2241], S[2242], S[2243], S[2789], Cout[2789]);
	Full_Adder FA2734 (S[2244], S[2245], S[2246], S[2790], Cout[2790]);
	Full_Adder FA2735 (S[1539], Cout[2242], Cout[2243], S[2791], Cout[2791]);
	Full_Adder FA2736 (Cout[2244], Cout[2245], Cout[2246], S[2792], Cout[2792]);
	Full_Adder FA2737 (Cout[2247], S[2248], S[2249], S[2793], Cout[2793]);
	Full_Adder FA2738 (S[2250], S[2251], S[2252], S[2794], Cout[2794]);
	Full_Adder FA2739 (S[1548], Cout[2248], Cout[2249], S[2795], Cout[2795]);
	Full_Adder FA2740 (Cout[2250], Cout[2251], Cout[2252], S[2796], Cout[2796]);
	Full_Adder FA2741 (Cout[2253], S[2254], S[2255], S[2797], Cout[2797]);
	Full_Adder FA2742 (S[2256], S[2257], S[2258], S[2798], Cout[2798]);
	Full_Adder FA2743 (S[1557], Cout[2254], Cout[2255], S[2799], Cout[2799]);
	Full_Adder FA2744 (Cout[2256], Cout[2257], Cout[2258], S[2800], Cout[2800]);
	Full_Adder FA2745 (Cout[2259], S[2260], S[2261], S[2801], Cout[2801]);
	Full_Adder FA2746 (S[2262], S[2263], S[2264], S[2802], Cout[2802]);
	Full_Adder FA2747 (S[1566], Cout[2260], Cout[2261], S[2803], Cout[2803]);
	Full_Adder FA2748 (Cout[2262], Cout[2263], Cout[2264], S[2804], Cout[2804]);
	Full_Adder FA2749 (Cout[2265], S[2266], S[2267], S[2805], Cout[2805]);
	Full_Adder FA2750 (S[2268], S[2269], S[2270], S[2806], Cout[2806]);
	Full_Adder FA2751 (S[1575], Cout[2266], Cout[2267], S[2807], Cout[2807]);
	Full_Adder FA2752 (Cout[2268], Cout[2269], Cout[2270], S[2808], Cout[2808]);
	Full_Adder FA2753 (Cout[2271], S[2272], S[2273], S[2809], Cout[2809]);
	Full_Adder FA2754 (S[2274], S[2275], S[2276], S[2810], Cout[2810]);
	Full_Adder FA2755 (S[1584], Cout[2272], Cout[2273], S[2811], Cout[2811]);
	Full_Adder FA2756 (Cout[2274], Cout[2275], Cout[2276], S[2812], Cout[2812]);
	Full_Adder FA2757 (Cout[2277], S[2278], S[2279], S[2813], Cout[2813]);
	Full_Adder FA2758 (S[2280], S[2281], S[2282], S[2814], Cout[2814]);
	Full_Adder FA2759 (S[1593], Cout[2278], Cout[2279], S[2815], Cout[2815]);
	Full_Adder FA2760 (Cout[2280], Cout[2281], Cout[2282], S[2816], Cout[2816]);
	Full_Adder FA2761 (Cout[2283], S[2284], S[2285], S[2817], Cout[2817]);
	Full_Adder FA2762 (S[2286], S[2287], S[2288], S[2818], Cout[2818]);
	Full_Adder FA2763 (S[1602], Cout[2284], Cout[2285], S[2819], Cout[2819]);
	Full_Adder FA2764 (Cout[2286], Cout[2287], Cout[2288], S[2820], Cout[2820]);
	Full_Adder FA2765 (Cout[2289], S[2290], S[2291], S[2821], Cout[2821]);
	Full_Adder FA2766 (S[2292], S[2293], S[2294], S[2822], Cout[2822]);
	Full_Adder FA2767 (S[1611], Cout[2290], Cout[2291], S[2823], Cout[2823]);
	Full_Adder FA2768 (Cout[2292], Cout[2293], Cout[2294], S[2824], Cout[2824]);
	Full_Adder FA2769 (Cout[2295], S[2296], S[2297], S[2825], Cout[2825]);
	Full_Adder FA2770 (S[2298], S[2299], S[2300], S[2826], Cout[2826]);
	Full_Adder FA2771 (S[1620], Cout[2296], Cout[2297], S[2827], Cout[2827]);
	Full_Adder FA2772 (Cout[2298], Cout[2299], Cout[2300], S[2828], Cout[2828]);
	Full_Adder FA2773 (Cout[2301], S[2302], S[2303], S[2829], Cout[2829]);
	Full_Adder FA2774 (S[2304], S[2305], S[2306], S[2830], Cout[2830]);
	Full_Adder FA2775 (S[1629], Cout[2302], Cout[2303], S[2831], Cout[2831]);
	Full_Adder FA2776 (Cout[2304], Cout[2305], Cout[2306], S[2832], Cout[2832]);
	Full_Adder FA2777 (Cout[2307], S[2308], S[2309], S[2833], Cout[2833]);
	Full_Adder FA2778 (S[2310], S[2311], S[2312], S[2834], Cout[2834]);
	Full_Adder FA2779 (S[1638], Cout[2308], Cout[2309], S[2835], Cout[2835]);
	Full_Adder FA2780 (Cout[2310], Cout[2311], Cout[2312], S[2836], Cout[2836]);
	Full_Adder FA2781 (Cout[2313], S[2314], S[2315], S[2837], Cout[2837]);
	Full_Adder FA2782 (S[2316], S[2317], S[2318], S[2838], Cout[2838]);
	Full_Adder FA2783 (S[1647], Cout[2314], Cout[2315], S[2839], Cout[2839]);
	Full_Adder FA2784 (Cout[2316], Cout[2317], Cout[2318], S[2840], Cout[2840]);
	Full_Adder FA2785 (Cout[2319], S[2320], S[2321], S[2841], Cout[2841]);
	Full_Adder FA2786 (S[2322], S[2323], S[2324], S[2842], Cout[2842]);
	Full_Adder FA2787 (S[1656], Cout[2320], Cout[2321], S[2843], Cout[2843]);
	Full_Adder FA2788 (Cout[2322], Cout[2323], Cout[2324], S[2844], Cout[2844]);
	Full_Adder FA2789 (Cout[2325], S[2326], S[2327], S[2845], Cout[2845]);
	Full_Adder FA2790 (S[2328], S[2329], S[2330], S[2846], Cout[2846]);
	Full_Adder FA2791 (S[1665], Cout[2326], Cout[2327], S[2847], Cout[2847]);
	Full_Adder FA2792 (Cout[2328], Cout[2329], Cout[2330], S[2848], Cout[2848]);
	Full_Adder FA2793 (Cout[2331], S[2332], S[2333], S[2849], Cout[2849]);
	Full_Adder FA2794 (S[2334], S[2335], S[2336], S[2850], Cout[2850]);
	Full_Adder FA2795 (S[1674], Cout[2332], Cout[2333], S[2851], Cout[2851]);
	Full_Adder FA2796 (Cout[2334], Cout[2335], Cout[2336], S[2852], Cout[2852]);
	Full_Adder FA2797 (Cout[2337], S[2338], S[2339], S[2853], Cout[2853]);
	Full_Adder FA2798 (S[2340], S[2341], S[2342], S[2854], Cout[2854]);
	Full_Adder FA2799 (S[1683], Cout[2338], Cout[2339], S[2855], Cout[2855]);
	Full_Adder FA2800 (Cout[2340], Cout[2341], Cout[2342], S[2856], Cout[2856]);
	Full_Adder FA2801 (Cout[2343], S[2344], S[2345], S[2857], Cout[2857]);
	Full_Adder FA2802 (S[2346], S[2347], S[2348], S[2858], Cout[2858]);
	Full_Adder FA2803 (S[1692], Cout[2344], Cout[2345], S[2859], Cout[2859]);
	Full_Adder FA2804 (Cout[2346], Cout[2347], Cout[2348], S[2860], Cout[2860]);
	Full_Adder FA2805 (Cout[2349], S[2350], S[2351], S[2861], Cout[2861]);
	Full_Adder FA2806 (S[2352], S[2353], S[2354], S[2862], Cout[2862]);
	Full_Adder FA2807 (S[1701], Cout[2350], Cout[2351], S[2863], Cout[2863]);
	Full_Adder FA2808 (Cout[2352], Cout[2353], Cout[2354], S[2864], Cout[2864]);
	Full_Adder FA2809 (Cout[2355], S[2356], S[2357], S[2865], Cout[2865]);
	Full_Adder FA2810 (S[2358], S[2359], S[2360], S[2866], Cout[2866]);
	Full_Adder FA2811 (S[1710], Cout[2356], Cout[2357], S[2867], Cout[2867]);
	Full_Adder FA2812 (Cout[2358], Cout[2359], Cout[2360], S[2868], Cout[2868]);
	Full_Adder FA2813 (Cout[2361], S[2362], S[2363], S[2869], Cout[2869]);
	Full_Adder FA2814 (S[2364], S[2365], S[2366], S[2870], Cout[2870]);
	Full_Adder FA2815 (S[1719], Cout[2362], Cout[2363], S[2871], Cout[2871]);
	Full_Adder FA2816 (Cout[2364], Cout[2365], Cout[2366], S[2872], Cout[2872]);
	Full_Adder FA2817 (Cout[2367], S[2368], S[2369], S[2873], Cout[2873]);
	Full_Adder FA2818 (S[2370], S[2371], S[2372], S[2874], Cout[2874]);
	Full_Adder FA2819 (S[1728], Cout[2368], Cout[2369], S[2875], Cout[2875]);
	Full_Adder FA2820 (Cout[2370], Cout[2371], Cout[2372], S[2876], Cout[2876]);
	Full_Adder FA2821 (Cout[2373], S[2374], S[2375], S[2877], Cout[2877]);
	Full_Adder FA2822 (S[2376], S[2377], S[2378], S[2878], Cout[2878]);
	Full_Adder FA2823 (S[1737], Cout[2374], Cout[2375], S[2879], Cout[2879]);
	Full_Adder FA2824 (Cout[2376], Cout[2377], Cout[2378], S[2880], Cout[2880]);
	Full_Adder FA2825 (Cout[2379], S[2380], S[2381], S[2881], Cout[2881]);
	Full_Adder FA2826 (S[2382], S[2383], S[2384], S[2882], Cout[2882]);
	Full_Adder FA2827 (S[1746], Cout[2380], Cout[2381], S[2883], Cout[2883]);
	Full_Adder FA2828 (Cout[2382], Cout[2383], Cout[2384], S[2884], Cout[2884]);
	Full_Adder FA2829 (Cout[2385], S[2386], S[2387], S[2885], Cout[2885]);
	Full_Adder FA2830 (S[2388], S[2389], S[2390], S[2886], Cout[2886]);
	Full_Adder FA2831 (S[1755], Cout[2386], Cout[2387], S[2887], Cout[2887]);
	Full_Adder FA2832 (Cout[2388], Cout[2389], Cout[2390], S[2888], Cout[2888]);
	Full_Adder FA2833 (Cout[2391], S[2392], S[2393], S[2889], Cout[2889]);
	Full_Adder FA2834 (S[2394], S[2395], S[2396], S[2890], Cout[2890]);
	Full_Adder FA2835 (S[1764], Cout[2392], Cout[2393], S[2891], Cout[2891]);
	Full_Adder FA2836 (Cout[2394], Cout[2395], Cout[2396], S[2892], Cout[2892]);
	Full_Adder FA2837 (Cout[2397], S[2398], S[2399], S[2893], Cout[2893]);
	Full_Adder FA2838 (S[2400], S[2401], S[2402], S[2894], Cout[2894]);
	Full_Adder FA2839 (S[1773], Cout[2398], Cout[2399], S[2895], Cout[2895]);
	Full_Adder FA2840 (Cout[2400], Cout[2401], Cout[2402], S[2896], Cout[2896]);
	Full_Adder FA2841 (Cout[2403], S[2404], S[2405], S[2897], Cout[2897]);
	Full_Adder FA2842 (S[2406], S[2407], S[2408], S[2898], Cout[2898]);
	Full_Adder FA2843 (S[1782], Cout[2404], Cout[2405], S[2899], Cout[2899]);
	Full_Adder FA2844 (Cout[2406], Cout[2407], Cout[2408], S[2900], Cout[2900]);
	Full_Adder FA2845 (Cout[2409], S[2410], S[2411], S[2901], Cout[2901]);
	Full_Adder FA2846 (S[2412], S[2413], S[2414], S[2902], Cout[2902]);
	Full_Adder FA2847 (S[1791], Cout[2410], Cout[2411], S[2903], Cout[2903]);
	Full_Adder FA2848 (Cout[2412], Cout[2413], Cout[2414], S[2904], Cout[2904]);
	Full_Adder FA2849 (Cout[2415], S[2416], S[2417], S[2905], Cout[2905]);
	Full_Adder FA2850 (S[2418], S[2419], S[2420], S[2906], Cout[2906]);
	Full_Adder FA2851 (S[1800], Cout[2416], Cout[2417], S[2907], Cout[2907]);
	Full_Adder FA2852 (Cout[2418], Cout[2419], Cout[2420], S[2908], Cout[2908]);
	Full_Adder FA2853 (Cout[2421], S[2422], S[2423], S[2909], Cout[2909]);
	Full_Adder FA2854 (S[2424], S[2425], S[2426], S[2910], Cout[2910]);
	Full_Adder FA2855 (S[1809], Cout[2422], Cout[2423], S[2911], Cout[2911]);
	Full_Adder FA2856 (Cout[2424], Cout[2425], Cout[2426], S[2912], Cout[2912]);
	Full_Adder FA2857 (Cout[2427], S[2428], S[2429], S[2913], Cout[2913]);
	Full_Adder FA2858 (S[2430], S[2431], S[2432], S[2914], Cout[2914]);
	Full_Adder FA2859 (S[1818], Cout[2428], Cout[2429], S[2915], Cout[2915]);
	Full_Adder FA2860 (Cout[2430], Cout[2431], Cout[2432], S[2916], Cout[2916]);
	Full_Adder FA2861 (Cout[2433], S[2434], S[2435], S[2917], Cout[2917]);
	Full_Adder FA2862 (S[2436], S[2437], S[2438], S[2918], Cout[2918]);
	Full_Adder FA2863 (S[1827], Cout[2434], Cout[2435], S[2919], Cout[2919]);
	Full_Adder FA2864 (Cout[2436], Cout[2437], Cout[2438], S[2920], Cout[2920]);
	Full_Adder FA2865 (Cout[2439], S[2440], S[2441], S[2921], Cout[2921]);
	Full_Adder FA2866 (S[2442], S[2443], S[2444], S[2922], Cout[2922]);
	Full_Adder FA2867 (S[1836], Cout[2440], Cout[2441], S[2923], Cout[2923]);
	Full_Adder FA2868 (Cout[2442], Cout[2443], Cout[2444], S[2924], Cout[2924]);
	Full_Adder FA2869 (Cout[2445], S[2446], S[2447], S[2925], Cout[2925]);
	Full_Adder FA2870 (S[2448], S[2449], S[2450], S[2926], Cout[2926]);
	Full_Adder FA2871 (S[1845], Cout[2446], Cout[2447], S[2927], Cout[2927]);
	Full_Adder FA2872 (Cout[2448], Cout[2449], Cout[2450], S[2928], Cout[2928]);
	Full_Adder FA2873 (Cout[2451], S[2452], S[2453], S[2929], Cout[2929]);
	Full_Adder FA2874 (S[2454], S[2455], S[2456], S[2930], Cout[2930]);
	Full_Adder FA2875 (S[1854], Cout[2452], Cout[2453], S[2931], Cout[2931]);
	Full_Adder FA2876 (Cout[2454], Cout[2455], Cout[2456], S[2932], Cout[2932]);
	Full_Adder FA2877 (Cout[2457], S[2458], S[2459], S[2933], Cout[2933]);
	Full_Adder FA2878 (S[2460], S[2461], S[2462], S[2934], Cout[2934]);
	Full_Adder FA2879 (S[1863], Cout[2458], Cout[2459], S[2935], Cout[2935]);
	Full_Adder FA2880 (Cout[2460], Cout[2461], Cout[2462], S[2936], Cout[2936]);
	Full_Adder FA2881 (Cout[2463], S[2464], S[2465], S[2937], Cout[2937]);
	Full_Adder FA2882 (S[2466], S[2467], S[2468], S[2938], Cout[2938]);
	Full_Adder FA2883 (S[1872], Cout[2464], Cout[2465], S[2939], Cout[2939]);
	Full_Adder FA2884 (Cout[2466], Cout[2467], Cout[2468], S[2940], Cout[2940]);
	Full_Adder FA2885 (Cout[2469], S[2470], S[2471], S[2941], Cout[2941]);
	Full_Adder FA2886 (S[2472], S[2473], S[2474], S[2942], Cout[2942]);
	Full_Adder FA2887 (S[1881], Cout[2470], Cout[2471], S[2943], Cout[2943]);
	Full_Adder FA2888 (Cout[2472], Cout[2473], Cout[2474], S[2944], Cout[2944]);
	Full_Adder FA2889 (Cout[2475], S[2476], S[2477], S[2945], Cout[2945]);
	Full_Adder FA2890 (S[2478], S[2479], S[2480], S[2946], Cout[2946]);
	Full_Adder FA2891 (S[1890], Cout[2476], Cout[2477], S[2947], Cout[2947]);
	Full_Adder FA2892 (Cout[2478], Cout[2479], Cout[2480], S[2948], Cout[2948]);
	Full_Adder FA2893 (Cout[2481], S[2482], S[2483], S[2949], Cout[2949]);
	Full_Adder FA2894 (S[2484], S[2485], S[2486], S[2950], Cout[2950]);
	Full_Adder FA2895 (S[1899], Cout[2482], Cout[2483], S[2951], Cout[2951]);
	Full_Adder FA2896 (Cout[2484], Cout[2485], Cout[2486], S[2952], Cout[2952]);
	Full_Adder FA2897 (Cout[2487], S[2488], S[2489], S[2953], Cout[2953]);
	Full_Adder FA2898 (S[2490], S[2491], S[2492], S[2954], Cout[2954]);
	Full_Adder FA2899 (S[1908], Cout[2488], Cout[2489], S[2955], Cout[2955]);
	Full_Adder FA2900 (Cout[2490], Cout[2491], Cout[2492], S[2956], Cout[2956]);
	Full_Adder FA2901 (Cout[2493], S[2494], S[2495], S[2957], Cout[2957]);
	Full_Adder FA2902 (S[2496], S[2497], S[2498], S[2958], Cout[2958]);
	Full_Adder FA2903 (S[1917], Cout[2494], Cout[2495], S[2959], Cout[2959]);
	Full_Adder FA2904 (Cout[2496], Cout[2497], Cout[2498], S[2960], Cout[2960]);
	Full_Adder FA2905 (Cout[2499], S[2500], S[2501], S[2961], Cout[2961]);
	Full_Adder FA2906 (S[2502], S[2503], S[2504], S[2962], Cout[2962]);
	Full_Adder FA2907 (S[1926], Cout[2500], Cout[2501], S[2963], Cout[2963]);
	Full_Adder FA2908 (Cout[2502], Cout[2503], Cout[2504], S[2964], Cout[2964]);
	Full_Adder FA2909 (Cout[2505], S[2506], S[2507], S[2965], Cout[2965]);
	Full_Adder FA2910 (S[2508], S[2509], S[2510], S[2966], Cout[2966]);
	Full_Adder FA2911 (S[1935], Cout[2506], Cout[2507], S[2967], Cout[2967]);
	Full_Adder FA2912 (Cout[2508], Cout[2509], Cout[2510], S[2968], Cout[2968]);
	Full_Adder FA2913 (Cout[2511], S[2512], S[2513], S[2969], Cout[2969]);
	Full_Adder FA2914 (S[2514], S[2515], S[2516], S[2970], Cout[2970]);
	Full_Adder FA2915 (S[1944], Cout[2512], Cout[2513], S[2971], Cout[2971]);
	Full_Adder FA2916 (Cout[2514], Cout[2515], Cout[2516], S[2972], Cout[2972]);
	Full_Adder FA2917 (Cout[2517], S[2518], S[2519], S[2973], Cout[2973]);
	Full_Adder FA2918 (S[2520], S[2521], S[2522], S[2974], Cout[2974]);
	Full_Adder FA2919 (S[1953], Cout[2518], Cout[2519], S[2975], Cout[2975]);
	Full_Adder FA2920 (Cout[2520], Cout[2521], Cout[2522], S[2976], Cout[2976]);
	Full_Adder FA2921 (Cout[2523], S[2524], S[2525], S[2977], Cout[2977]);
	Full_Adder FA2922 (S[2526], S[2527], S[2528], S[2978], Cout[2978]);
	Full_Adder FA2923 (S[1962], Cout[2524], Cout[2525], S[2979], Cout[2979]);
	Full_Adder FA2924 (Cout[2526], Cout[2527], Cout[2528], S[2980], Cout[2980]);
	Full_Adder FA2925 (Cout[2529], S[2530], S[2531], S[2981], Cout[2981]);
	Full_Adder FA2926 (S[2532], S[2533], S[2534], S[2982], Cout[2982]);
	Full_Adder FA2927 (S[1971], Cout[2530], Cout[2531], S[2983], Cout[2983]);
	Full_Adder FA2928 (Cout[2532], Cout[2533], Cout[2534], S[2984], Cout[2984]);
	Full_Adder FA2929 (Cout[2535], S[2536], S[2537], S[2985], Cout[2985]);
	Full_Adder FA2930 (S[2538], S[2539], S[2540], S[2986], Cout[2986]);
	Full_Adder FA2931 (S[1980], Cout[2536], Cout[2537], S[2987], Cout[2987]);
	Full_Adder FA2932 (Cout[2538], Cout[2539], Cout[2540], S[2988], Cout[2988]);
	Full_Adder FA2933 (Cout[2541], S[2542], S[2543], S[2989], Cout[2989]);
	Full_Adder FA2934 (S[2544], S[2545], S[2546], S[2990], Cout[2990]);
	Full_Adder FA2935 (S[1989], Cout[2542], Cout[2543], S[2991], Cout[2991]);
	Full_Adder FA2936 (Cout[2544], Cout[2545], Cout[2546], S[2992], Cout[2992]);
	Full_Adder FA2937 (Cout[2547], S[2548], S[2549], S[2993], Cout[2993]);
	Full_Adder FA2938 (S[2550], S[2551], S[2552], S[2994], Cout[2994]);
	Full_Adder FA2939 (S[1998], Cout[2548], Cout[2549], S[2995], Cout[2995]);
	Full_Adder FA2940 (Cout[2550], Cout[2551], Cout[2552], S[2996], Cout[2996]);
	Full_Adder FA2941 (Cout[2553], S[2554], S[2555], S[2997], Cout[2997]);
	Full_Adder FA2942 (S[2556], S[2557], S[2558], S[2998], Cout[2998]);
	Full_Adder FA2943 (S[2007], Cout[2554], Cout[2555], S[2999], Cout[2999]);
	Full_Adder FA2944 (Cout[2556], Cout[2557], Cout[2558], S[3000], Cout[3000]);
	Full_Adder FA2945 (Cout[2559], S[2560], S[2561], S[3001], Cout[3001]);
	Full_Adder FA2946 (S[2562], S[2563], S[2564], S[3002], Cout[3002]);
	Full_Adder FA2947 (S[2016], Cout[2560], Cout[2561], S[3003], Cout[3003]);
	Full_Adder FA2948 (Cout[2562], Cout[2563], Cout[2564], S[3004], Cout[3004]);
	Full_Adder FA2949 (Cout[2565], S[2566], S[2567], S[3005], Cout[3005]);
	Full_Adder FA2950 (S[2568], S[2569], S[2570], S[3006], Cout[3006]);
	Full_Adder FA2951 (S[2025], Cout[2566], Cout[2567], S[3007], Cout[3007]);
	Full_Adder FA2952 (Cout[2568], Cout[2569], Cout[2570], S[3008], Cout[3008]);
	Full_Adder FA2953 (Cout[2571], S[2572], S[2573], S[3009], Cout[3009]);
	Full_Adder FA2954 (S[2574], S[2575], S[2576], S[3010], Cout[3010]);
	Full_Adder FA2955 (S[2034], Cout[2572], Cout[2573], S[3011], Cout[3011]);
	Full_Adder FA2956 (Cout[2574], Cout[2575], Cout[2576], S[3012], Cout[3012]);
	Full_Adder FA2957 (Cout[2577], S[2578], S[2579], S[3013], Cout[3013]);
	Full_Adder FA2958 (S[2580], S[2581], S[2582], S[3014], Cout[3014]);
	Full_Adder FA2959 (S[2042], Cout[2578], Cout[2579], S[3015], Cout[3015]);
	Full_Adder FA2960 (Cout[2580], Cout[2581], Cout[2582], S[3016], Cout[3016]);
	Full_Adder FA2961 (Cout[2583], S[2584], S[2585], S[3017], Cout[3017]);
	Full_Adder FA2962 (S[2586], S[2587], S[2588], S[3018], Cout[3018]);
	Full_Adder FA2963 (S[2049], Cout[2584], Cout[2585], S[3019], Cout[3019]);
	Full_Adder FA2964 (Cout[2586], Cout[2587], Cout[2588], S[3020], Cout[3020]);
	Full_Adder FA2965 (Cout[2589], S[2590], S[2591], S[3021], Cout[3021]);
	Full_Adder FA2966 (S[2592], S[2593], S[2594], S[3022], Cout[3022]);
	Full_Adder FA2967 (S[2055], Cout[2590], Cout[2591], S[3023], Cout[3023]);
	Full_Adder FA2968 (Cout[2592], Cout[2593], Cout[2594], S[3024], Cout[3024]);
	Full_Adder FA2969 (Cout[2595], S[2596], S[2597], S[3025], Cout[3025]);
	Full_Adder FA2970 (S[2598], S[2599], S[2600], S[3026], Cout[3026]);
	Full_Adder FA2971 (S[2060], Cout[2596], Cout[2597], S[3027], Cout[3027]);
	Full_Adder FA2972 (Cout[2598], Cout[2599], Cout[2600], S[3028], Cout[3028]);
	Full_Adder FA2973 (Cout[2601], S[2602], S[2603], S[3029], Cout[3029]);
	Full_Adder FA2974 (S[2604], S[2605], S[2606], S[3030], Cout[3030]);
	Full_Adder FA2975 (S[2064], Cout[2602], Cout[2603], S[3031], Cout[3031]);
	Full_Adder FA2976 (Cout[2604], Cout[2605], Cout[2606], S[3032], Cout[3032]);
	Full_Adder FA2977 (Cout[2607], S[2608], S[2609], S[3033], Cout[3033]);
	Full_Adder FA2978 (S[2610], S[2611], S[2612], S[3034], Cout[3034]);
	Full_Adder FA2979 (S[2067], Cout[2608], Cout[2609], S[3035], Cout[3035]);
	Full_Adder FA2980 (Cout[2610], Cout[2611], Cout[2612], S[3036], Cout[3036]);
	Full_Adder FA2981 (Cout[2613], S[2614], S[2615], S[3037], Cout[3037]);
	Full_Adder FA2982 (S[2616], S[2617], S[2618], S[3038], Cout[3038]);
	Full_Adder FA2983 (S[2069], Cout[2614], Cout[2615], S[3039], Cout[3039]);
	Full_Adder FA2984 (Cout[2616], Cout[2617], Cout[2618], S[3040], Cout[3040]);
	Full_Adder FA2985 (Cout[2619], S[2620], S[2621], S[3041], Cout[3041]);
	Full_Adder FA2986 (S[2622], S[2623], S[2624], S[3042], Cout[3042]);
	Full_Adder FA2987 (S[2070], Cout[2620], Cout[2621], S[3043], Cout[3043]);
	Full_Adder FA2988 (Cout[2622], Cout[2623], Cout[2624], S[3044], Cout[3044]);
	Full_Adder FA2989 (Cout[2625], S[2626], S[2627], S[3045], Cout[3045]);
	Full_Adder FA2990 (S[2628], S[2629], S[2630], S[3046], Cout[3046]);
	Full_Adder FA2991 (Cout[2070], Cout[2626], Cout[2627], S[3047], Cout[3047]);
	Full_Adder FA2992 (Cout[2628], Cout[2629], Cout[2630], S[3048], Cout[3048]);
	Full_Adder FA2993 (Cout[2631], S[2632], S[2633], S[3049], Cout[3049]);
	Full_Adder FA2994 (S[2634], S[2635], S[2636], S[3050], Cout[3050]);
	Full_Adder FA2995 (pp62[48], pp63[47], Cout[2632], S[3051], Cout[3051]);
	Full_Adder FA2996 (Cout[2633], Cout[2634], Cout[2635], S[3052], Cout[3052]);
	Full_Adder FA2997 (Cout[2636], Cout[2637], S[2638], S[3053], Cout[3053]);
	Full_Adder FA2998 (S[2639], S[2640], S[2641], S[3054], Cout[3054]);
	Full_Adder FA2999 (pp60[51], pp61[50], pp62[49], S[3055], Cout[3055]);
	Full_Adder FA3000 (pp63[48], Cout[2638], Cout[2639], S[3056], Cout[3056]);
	Full_Adder FA3001 (Cout[2640], Cout[2641], Cout[2642], S[3057], Cout[3057]);
	Full_Adder FA3002 (S[2643], S[2644], S[2645], S[3058], Cout[3058]);
	Full_Adder FA3003 (pp58[54], pp59[53], pp60[52], S[3059], Cout[3059]);
	Full_Adder FA3004 (pp61[51], pp62[50], pp63[49], S[3060], Cout[3060]);
	Full_Adder FA3005 (Cout[2643], Cout[2644], Cout[2645], S[3061], Cout[3061]);
	Full_Adder FA3006 (Cout[2646], S[2647], S[2648], S[3062], Cout[3062]);
	Full_Adder FA3007 (pp56[57], pp57[56], pp58[55], S[3063], Cout[3063]);
	Full_Adder FA3008 (pp59[54], pp60[53], pp61[52], S[3064], Cout[3064]);
	Full_Adder FA3009 (pp62[51], pp63[50], Cout[2647], S[3065], Cout[3065]);
	Full_Adder FA3010 (Cout[2648], Cout[2649], S[2650], S[3066], Cout[3066]);
	Full_Adder FA3011 (pp54[60], pp55[59], pp56[58], S[3067], Cout[3067]);
	Full_Adder FA3012 (pp57[57], pp58[56], pp59[55], S[3068], Cout[3068]);
	Full_Adder FA3013 (pp60[54], pp61[53], pp62[52], S[3069], Cout[3069]);
	Full_Adder FA3014 (pp63[51], Cout[2650], Cout[2651], S[3070], Cout[3070]);
	Full_Adder FA3015 (pp52[63], pp53[62], pp54[61], S[3071], Cout[3071]);
	Full_Adder FA3016 (pp55[60], pp56[59], pp57[58], S[3072], Cout[3072]);
	Full_Adder FA3017 (pp58[57], pp59[56], pp60[55], S[3073], Cout[3073]);
	Full_Adder FA3018 (pp61[54], pp62[53], pp63[52], S[3074], Cout[3074]);
	Full_Adder FA3019 (pp53[63], pp54[62], pp55[61], S[3075], Cout[3075]);
	Full_Adder FA3020 (pp56[60], pp57[59], pp58[58], S[3076], Cout[3076]);
	Full_Adder FA3021 (pp59[57], pp60[56], pp61[55], S[3077], Cout[3077]);
	Full_Adder FA3022 (pp54[63], pp55[62], pp56[61], S[3078], Cout[3078]);
	Full_Adder FA3023 (pp57[60], pp58[59], pp59[58], S[3079], Cout[3079]);
	Full_Adder FA3024 (pp55[63], pp56[62], pp57[61], S[3080], Cout[3080]);
	Half_Adder HA57 (pp0[6], pp1[5], S[3081], Cout[3081]);
	Full_Adder FA3025 (pp0[7], pp1[6], pp2[5], S[3082], Cout[3082]);
	Half_Adder HA58 (pp3[4], pp4[3], S[3083], Cout[3083]);
	Full_Adder FA3026 (pp0[8], pp1[7], pp2[6], S[3084], Cout[3084]);
	Full_Adder FA3027 (pp3[5], pp4[4], pp5[3], S[3085], Cout[3085]);
	Half_Adder HA59 (pp6[2], pp7[1], S[3086], Cout[3086]);
	Full_Adder FA3028 (pp2[7], pp3[6], pp4[5], S[3087], Cout[3087]);
	Full_Adder FA3029 (pp5[4], pp6[3], pp7[2], S[3088], Cout[3088]);
	Full_Adder FA3030 (pp8[1], pp9[0], S[2653], S[3089], Cout[3089]);
	Full_Adder FA3031 (pp5[5], pp6[4], pp7[3], S[3090], Cout[3090]);
	Full_Adder FA3032 (pp8[2], pp9[1], pp10[0], S[3091], Cout[3091]);
	Full_Adder FA3033 (Cout[2653], S[2654], S[2655], S[3092], Cout[3092]);
	Full_Adder FA3034 (pp8[3], pp9[2], pp10[1], S[3093], Cout[3093]);
	Full_Adder FA3035 (pp11[0], Cout[2654], Cout[2655], S[3094], Cout[3094]);
	Full_Adder FA3036 (S[2656], S[2657], S[2658], S[3095], Cout[3095]);
	Full_Adder FA3037 (pp11[1], pp12[0], Cout[2656], S[3096], Cout[3096]);
	Full_Adder FA3038 (Cout[2657], Cout[2658], S[2659], S[3097], Cout[3097]);
	Full_Adder FA3039 (S[2660], S[2661], S[2662], S[3098], Cout[3098]);
	Full_Adder FA3040 (S[2071], Cout[2659], Cout[2660], S[3099], Cout[3099]);
	Full_Adder FA3041 (Cout[2661], Cout[2662], S[2663], S[3100], Cout[3100]);
	Full_Adder FA3042 (S[2664], S[2665], S[2666], S[3101], Cout[3101]);
	Full_Adder FA3043 (S[2073], Cout[2663], Cout[2664], S[3102], Cout[3102]);
	Full_Adder FA3044 (Cout[2665], Cout[2666], S[2667], S[3103], Cout[3103]);
	Full_Adder FA3045 (S[2668], S[2669], S[2670], S[3104], Cout[3104]);
	Full_Adder FA3046 (S[2076], Cout[2667], Cout[2668], S[3105], Cout[3105]);
	Full_Adder FA3047 (Cout[2669], Cout[2670], S[2671], S[3106], Cout[3106]);
	Full_Adder FA3048 (S[2672], S[2673], S[2674], S[3107], Cout[3107]);
	Full_Adder FA3049 (S[2080], Cout[2671], Cout[2672], S[3108], Cout[3108]);
	Full_Adder FA3050 (Cout[2673], Cout[2674], S[2675], S[3109], Cout[3109]);
	Full_Adder FA3051 (S[2676], S[2677], S[2678], S[3110], Cout[3110]);
	Full_Adder FA3052 (S[2085], Cout[2675], Cout[2676], S[3111], Cout[3111]);
	Full_Adder FA3053 (Cout[2677], Cout[2678], S[2679], S[3112], Cout[3112]);
	Full_Adder FA3054 (S[2680], S[2681], S[2682], S[3113], Cout[3113]);
	Full_Adder FA3055 (S[2091], Cout[2679], Cout[2680], S[3114], Cout[3114]);
	Full_Adder FA3056 (Cout[2681], Cout[2682], S[2683], S[3115], Cout[3115]);
	Full_Adder FA3057 (S[2684], S[2685], S[2686], S[3116], Cout[3116]);
	Full_Adder FA3058 (S[2097], Cout[2683], Cout[2684], S[3117], Cout[3117]);
	Full_Adder FA3059 (Cout[2685], Cout[2686], S[2687], S[3118], Cout[3118]);
	Full_Adder FA3060 (S[2688], S[2689], S[2690], S[3119], Cout[3119]);
	Full_Adder FA3061 (S[2103], Cout[2687], Cout[2688], S[3120], Cout[3120]);
	Full_Adder FA3062 (Cout[2689], Cout[2690], S[2691], S[3121], Cout[3121]);
	Full_Adder FA3063 (S[2692], S[2693], S[2694], S[3122], Cout[3122]);
	Full_Adder FA3064 (S[2109], Cout[2691], Cout[2692], S[3123], Cout[3123]);
	Full_Adder FA3065 (Cout[2693], Cout[2694], S[2695], S[3124], Cout[3124]);
	Full_Adder FA3066 (S[2696], S[2697], S[2698], S[3125], Cout[3125]);
	Full_Adder FA3067 (S[2115], Cout[2695], Cout[2696], S[3126], Cout[3126]);
	Full_Adder FA3068 (Cout[2697], Cout[2698], S[2699], S[3127], Cout[3127]);
	Full_Adder FA3069 (S[2700], S[2701], S[2702], S[3128], Cout[3128]);
	Full_Adder FA3070 (S[2121], Cout[2699], Cout[2700], S[3129], Cout[3129]);
	Full_Adder FA3071 (Cout[2701], Cout[2702], S[2703], S[3130], Cout[3130]);
	Full_Adder FA3072 (S[2704], S[2705], S[2706], S[3131], Cout[3131]);
	Full_Adder FA3073 (S[2127], Cout[2703], Cout[2704], S[3132], Cout[3132]);
	Full_Adder FA3074 (Cout[2705], Cout[2706], S[2707], S[3133], Cout[3133]);
	Full_Adder FA3075 (S[2708], S[2709], S[2710], S[3134], Cout[3134]);
	Full_Adder FA3076 (S[2133], Cout[2707], Cout[2708], S[3135], Cout[3135]);
	Full_Adder FA3077 (Cout[2709], Cout[2710], S[2711], S[3136], Cout[3136]);
	Full_Adder FA3078 (S[2712], S[2713], S[2714], S[3137], Cout[3137]);
	Full_Adder FA3079 (S[2139], Cout[2711], Cout[2712], S[3138], Cout[3138]);
	Full_Adder FA3080 (Cout[2713], Cout[2714], S[2715], S[3139], Cout[3139]);
	Full_Adder FA3081 (S[2716], S[2717], S[2718], S[3140], Cout[3140]);
	Full_Adder FA3082 (S[2145], Cout[2715], Cout[2716], S[3141], Cout[3141]);
	Full_Adder FA3083 (Cout[2717], Cout[2718], S[2719], S[3142], Cout[3142]);
	Full_Adder FA3084 (S[2720], S[2721], S[2722], S[3143], Cout[3143]);
	Full_Adder FA3085 (S[2151], Cout[2719], Cout[2720], S[3144], Cout[3144]);
	Full_Adder FA3086 (Cout[2721], Cout[2722], S[2723], S[3145], Cout[3145]);
	Full_Adder FA3087 (S[2724], S[2725], S[2726], S[3146], Cout[3146]);
	Full_Adder FA3088 (S[2157], Cout[2723], Cout[2724], S[3147], Cout[3147]);
	Full_Adder FA3089 (Cout[2725], Cout[2726], S[2727], S[3148], Cout[3148]);
	Full_Adder FA3090 (S[2728], S[2729], S[2730], S[3149], Cout[3149]);
	Full_Adder FA3091 (S[2163], Cout[2727], Cout[2728], S[3150], Cout[3150]);
	Full_Adder FA3092 (Cout[2729], Cout[2730], S[2731], S[3151], Cout[3151]);
	Full_Adder FA3093 (S[2732], S[2733], S[2734], S[3152], Cout[3152]);
	Full_Adder FA3094 (S[2169], Cout[2731], Cout[2732], S[3153], Cout[3153]);
	Full_Adder FA3095 (Cout[2733], Cout[2734], S[2735], S[3154], Cout[3154]);
	Full_Adder FA3096 (S[2736], S[2737], S[2738], S[3155], Cout[3155]);
	Full_Adder FA3097 (S[2175], Cout[2735], Cout[2736], S[3156], Cout[3156]);
	Full_Adder FA3098 (Cout[2737], Cout[2738], S[2739], S[3157], Cout[3157]);
	Full_Adder FA3099 (S[2740], S[2741], S[2742], S[3158], Cout[3158]);
	Full_Adder FA3100 (S[2181], Cout[2739], Cout[2740], S[3159], Cout[3159]);
	Full_Adder FA3101 (Cout[2741], Cout[2742], S[2743], S[3160], Cout[3160]);
	Full_Adder FA3102 (S[2744], S[2745], S[2746], S[3161], Cout[3161]);
	Full_Adder FA3103 (S[2187], Cout[2743], Cout[2744], S[3162], Cout[3162]);
	Full_Adder FA3104 (Cout[2745], Cout[2746], S[2747], S[3163], Cout[3163]);
	Full_Adder FA3105 (S[2748], S[2749], S[2750], S[3164], Cout[3164]);
	Full_Adder FA3106 (S[2193], Cout[2747], Cout[2748], S[3165], Cout[3165]);
	Full_Adder FA3107 (Cout[2749], Cout[2750], S[2751], S[3166], Cout[3166]);
	Full_Adder FA3108 (S[2752], S[2753], S[2754], S[3167], Cout[3167]);
	Full_Adder FA3109 (S[2199], Cout[2751], Cout[2752], S[3168], Cout[3168]);
	Full_Adder FA3110 (Cout[2753], Cout[2754], S[2755], S[3169], Cout[3169]);
	Full_Adder FA3111 (S[2756], S[2757], S[2758], S[3170], Cout[3170]);
	Full_Adder FA3112 (S[2205], Cout[2755], Cout[2756], S[3171], Cout[3171]);
	Full_Adder FA3113 (Cout[2757], Cout[2758], S[2759], S[3172], Cout[3172]);
	Full_Adder FA3114 (S[2760], S[2761], S[2762], S[3173], Cout[3173]);
	Full_Adder FA3115 (S[2211], Cout[2759], Cout[2760], S[3174], Cout[3174]);
	Full_Adder FA3116 (Cout[2761], Cout[2762], S[2763], S[3175], Cout[3175]);
	Full_Adder FA3117 (S[2764], S[2765], S[2766], S[3176], Cout[3176]);
	Full_Adder FA3118 (S[2217], Cout[2763], Cout[2764], S[3177], Cout[3177]);
	Full_Adder FA3119 (Cout[2765], Cout[2766], S[2767], S[3178], Cout[3178]);
	Full_Adder FA3120 (S[2768], S[2769], S[2770], S[3179], Cout[3179]);
	Full_Adder FA3121 (S[2223], Cout[2767], Cout[2768], S[3180], Cout[3180]);
	Full_Adder FA3122 (Cout[2769], Cout[2770], S[2771], S[3181], Cout[3181]);
	Full_Adder FA3123 (S[2772], S[2773], S[2774], S[3182], Cout[3182]);
	Full_Adder FA3124 (S[2229], Cout[2771], Cout[2772], S[3183], Cout[3183]);
	Full_Adder FA3125 (Cout[2773], Cout[2774], S[2775], S[3184], Cout[3184]);
	Full_Adder FA3126 (S[2776], S[2777], S[2778], S[3185], Cout[3185]);
	Full_Adder FA3127 (S[2235], Cout[2775], Cout[2776], S[3186], Cout[3186]);
	Full_Adder FA3128 (Cout[2777], Cout[2778], S[2779], S[3187], Cout[3187]);
	Full_Adder FA3129 (S[2780], S[2781], S[2782], S[3188], Cout[3188]);
	Full_Adder FA3130 (S[2241], Cout[2779], Cout[2780], S[3189], Cout[3189]);
	Full_Adder FA3131 (Cout[2781], Cout[2782], S[2783], S[3190], Cout[3190]);
	Full_Adder FA3132 (S[2784], S[2785], S[2786], S[3191], Cout[3191]);
	Full_Adder FA3133 (S[2247], Cout[2783], Cout[2784], S[3192], Cout[3192]);
	Full_Adder FA3134 (Cout[2785], Cout[2786], S[2787], S[3193], Cout[3193]);
	Full_Adder FA3135 (S[2788], S[2789], S[2790], S[3194], Cout[3194]);
	Full_Adder FA3136 (S[2253], Cout[2787], Cout[2788], S[3195], Cout[3195]);
	Full_Adder FA3137 (Cout[2789], Cout[2790], S[2791], S[3196], Cout[3196]);
	Full_Adder FA3138 (S[2792], S[2793], S[2794], S[3197], Cout[3197]);
	Full_Adder FA3139 (S[2259], Cout[2791], Cout[2792], S[3198], Cout[3198]);
	Full_Adder FA3140 (Cout[2793], Cout[2794], S[2795], S[3199], Cout[3199]);
	Full_Adder FA3141 (S[2796], S[2797], S[2798], S[3200], Cout[3200]);
	Full_Adder FA3142 (S[2265], Cout[2795], Cout[2796], S[3201], Cout[3201]);
	Full_Adder FA3143 (Cout[2797], Cout[2798], S[2799], S[3202], Cout[3202]);
	Full_Adder FA3144 (S[2800], S[2801], S[2802], S[3203], Cout[3203]);
	Full_Adder FA3145 (S[2271], Cout[2799], Cout[2800], S[3204], Cout[3204]);
	Full_Adder FA3146 (Cout[2801], Cout[2802], S[2803], S[3205], Cout[3205]);
	Full_Adder FA3147 (S[2804], S[2805], S[2806], S[3206], Cout[3206]);
	Full_Adder FA3148 (S[2277], Cout[2803], Cout[2804], S[3207], Cout[3207]);
	Full_Adder FA3149 (Cout[2805], Cout[2806], S[2807], S[3208], Cout[3208]);
	Full_Adder FA3150 (S[2808], S[2809], S[2810], S[3209], Cout[3209]);
	Full_Adder FA3151 (S[2283], Cout[2807], Cout[2808], S[3210], Cout[3210]);
	Full_Adder FA3152 (Cout[2809], Cout[2810], S[2811], S[3211], Cout[3211]);
	Full_Adder FA3153 (S[2812], S[2813], S[2814], S[3212], Cout[3212]);
	Full_Adder FA3154 (S[2289], Cout[2811], Cout[2812], S[3213], Cout[3213]);
	Full_Adder FA3155 (Cout[2813], Cout[2814], S[2815], S[3214], Cout[3214]);
	Full_Adder FA3156 (S[2816], S[2817], S[2818], S[3215], Cout[3215]);
	Full_Adder FA3157 (S[2295], Cout[2815], Cout[2816], S[3216], Cout[3216]);
	Full_Adder FA3158 (Cout[2817], Cout[2818], S[2819], S[3217], Cout[3217]);
	Full_Adder FA3159 (S[2820], S[2821], S[2822], S[3218], Cout[3218]);
	Full_Adder FA3160 (S[2301], Cout[2819], Cout[2820], S[3219], Cout[3219]);
	Full_Adder FA3161 (Cout[2821], Cout[2822], S[2823], S[3220], Cout[3220]);
	Full_Adder FA3162 (S[2824], S[2825], S[2826], S[3221], Cout[3221]);
	Full_Adder FA3163 (S[2307], Cout[2823], Cout[2824], S[3222], Cout[3222]);
	Full_Adder FA3164 (Cout[2825], Cout[2826], S[2827], S[3223], Cout[3223]);
	Full_Adder FA3165 (S[2828], S[2829], S[2830], S[3224], Cout[3224]);
	Full_Adder FA3166 (S[2313], Cout[2827], Cout[2828], S[3225], Cout[3225]);
	Full_Adder FA3167 (Cout[2829], Cout[2830], S[2831], S[3226], Cout[3226]);
	Full_Adder FA3168 (S[2832], S[2833], S[2834], S[3227], Cout[3227]);
	Full_Adder FA3169 (S[2319], Cout[2831], Cout[2832], S[3228], Cout[3228]);
	Full_Adder FA3170 (Cout[2833], Cout[2834], S[2835], S[3229], Cout[3229]);
	Full_Adder FA3171 (S[2836], S[2837], S[2838], S[3230], Cout[3230]);
	Full_Adder FA3172 (S[2325], Cout[2835], Cout[2836], S[3231], Cout[3231]);
	Full_Adder FA3173 (Cout[2837], Cout[2838], S[2839], S[3232], Cout[3232]);
	Full_Adder FA3174 (S[2840], S[2841], S[2842], S[3233], Cout[3233]);
	Full_Adder FA3175 (S[2331], Cout[2839], Cout[2840], S[3234], Cout[3234]);
	Full_Adder FA3176 (Cout[2841], Cout[2842], S[2843], S[3235], Cout[3235]);
	Full_Adder FA3177 (S[2844], S[2845], S[2846], S[3236], Cout[3236]);
	Full_Adder FA3178 (S[2337], Cout[2843], Cout[2844], S[3237], Cout[3237]);
	Full_Adder FA3179 (Cout[2845], Cout[2846], S[2847], S[3238], Cout[3238]);
	Full_Adder FA3180 (S[2848], S[2849], S[2850], S[3239], Cout[3239]);
	Full_Adder FA3181 (S[2343], Cout[2847], Cout[2848], S[3240], Cout[3240]);
	Full_Adder FA3182 (Cout[2849], Cout[2850], S[2851], S[3241], Cout[3241]);
	Full_Adder FA3183 (S[2852], S[2853], S[2854], S[3242], Cout[3242]);
	Full_Adder FA3184 (S[2349], Cout[2851], Cout[2852], S[3243], Cout[3243]);
	Full_Adder FA3185 (Cout[2853], Cout[2854], S[2855], S[3244], Cout[3244]);
	Full_Adder FA3186 (S[2856], S[2857], S[2858], S[3245], Cout[3245]);
	Full_Adder FA3187 (S[2355], Cout[2855], Cout[2856], S[3246], Cout[3246]);
	Full_Adder FA3188 (Cout[2857], Cout[2858], S[2859], S[3247], Cout[3247]);
	Full_Adder FA3189 (S[2860], S[2861], S[2862], S[3248], Cout[3248]);
	Full_Adder FA3190 (S[2361], Cout[2859], Cout[2860], S[3249], Cout[3249]);
	Full_Adder FA3191 (Cout[2861], Cout[2862], S[2863], S[3250], Cout[3250]);
	Full_Adder FA3192 (S[2864], S[2865], S[2866], S[3251], Cout[3251]);
	Full_Adder FA3193 (S[2367], Cout[2863], Cout[2864], S[3252], Cout[3252]);
	Full_Adder FA3194 (Cout[2865], Cout[2866], S[2867], S[3253], Cout[3253]);
	Full_Adder FA3195 (S[2868], S[2869], S[2870], S[3254], Cout[3254]);
	Full_Adder FA3196 (S[2373], Cout[2867], Cout[2868], S[3255], Cout[3255]);
	Full_Adder FA3197 (Cout[2869], Cout[2870], S[2871], S[3256], Cout[3256]);
	Full_Adder FA3198 (S[2872], S[2873], S[2874], S[3257], Cout[3257]);
	Full_Adder FA3199 (S[2379], Cout[2871], Cout[2872], S[3258], Cout[3258]);
	Full_Adder FA3200 (Cout[2873], Cout[2874], S[2875], S[3259], Cout[3259]);
	Full_Adder FA3201 (S[2876], S[2877], S[2878], S[3260], Cout[3260]);
	Full_Adder FA3202 (S[2385], Cout[2875], Cout[2876], S[3261], Cout[3261]);
	Full_Adder FA3203 (Cout[2877], Cout[2878], S[2879], S[3262], Cout[3262]);
	Full_Adder FA3204 (S[2880], S[2881], S[2882], S[3263], Cout[3263]);
	Full_Adder FA3205 (S[2391], Cout[2879], Cout[2880], S[3264], Cout[3264]);
	Full_Adder FA3206 (Cout[2881], Cout[2882], S[2883], S[3265], Cout[3265]);
	Full_Adder FA3207 (S[2884], S[2885], S[2886], S[3266], Cout[3266]);
	Full_Adder FA3208 (S[2397], Cout[2883], Cout[2884], S[3267], Cout[3267]);
	Full_Adder FA3209 (Cout[2885], Cout[2886], S[2887], S[3268], Cout[3268]);
	Full_Adder FA3210 (S[2888], S[2889], S[2890], S[3269], Cout[3269]);
	Full_Adder FA3211 (S[2403], Cout[2887], Cout[2888], S[3270], Cout[3270]);
	Full_Adder FA3212 (Cout[2889], Cout[2890], S[2891], S[3271], Cout[3271]);
	Full_Adder FA3213 (S[2892], S[2893], S[2894], S[3272], Cout[3272]);
	Full_Adder FA3214 (S[2409], Cout[2891], Cout[2892], S[3273], Cout[3273]);
	Full_Adder FA3215 (Cout[2893], Cout[2894], S[2895], S[3274], Cout[3274]);
	Full_Adder FA3216 (S[2896], S[2897], S[2898], S[3275], Cout[3275]);
	Full_Adder FA3217 (S[2415], Cout[2895], Cout[2896], S[3276], Cout[3276]);
	Full_Adder FA3218 (Cout[2897], Cout[2898], S[2899], S[3277], Cout[3277]);
	Full_Adder FA3219 (S[2900], S[2901], S[2902], S[3278], Cout[3278]);
	Full_Adder FA3220 (S[2421], Cout[2899], Cout[2900], S[3279], Cout[3279]);
	Full_Adder FA3221 (Cout[2901], Cout[2902], S[2903], S[3280], Cout[3280]);
	Full_Adder FA3222 (S[2904], S[2905], S[2906], S[3281], Cout[3281]);
	Full_Adder FA3223 (S[2427], Cout[2903], Cout[2904], S[3282], Cout[3282]);
	Full_Adder FA3224 (Cout[2905], Cout[2906], S[2907], S[3283], Cout[3283]);
	Full_Adder FA3225 (S[2908], S[2909], S[2910], S[3284], Cout[3284]);
	Full_Adder FA3226 (S[2433], Cout[2907], Cout[2908], S[3285], Cout[3285]);
	Full_Adder FA3227 (Cout[2909], Cout[2910], S[2911], S[3286], Cout[3286]);
	Full_Adder FA3228 (S[2912], S[2913], S[2914], S[3287], Cout[3287]);
	Full_Adder FA3229 (S[2439], Cout[2911], Cout[2912], S[3288], Cout[3288]);
	Full_Adder FA3230 (Cout[2913], Cout[2914], S[2915], S[3289], Cout[3289]);
	Full_Adder FA3231 (S[2916], S[2917], S[2918], S[3290], Cout[3290]);
	Full_Adder FA3232 (S[2445], Cout[2915], Cout[2916], S[3291], Cout[3291]);
	Full_Adder FA3233 (Cout[2917], Cout[2918], S[2919], S[3292], Cout[3292]);
	Full_Adder FA3234 (S[2920], S[2921], S[2922], S[3293], Cout[3293]);
	Full_Adder FA3235 (S[2451], Cout[2919], Cout[2920], S[3294], Cout[3294]);
	Full_Adder FA3236 (Cout[2921], Cout[2922], S[2923], S[3295], Cout[3295]);
	Full_Adder FA3237 (S[2924], S[2925], S[2926], S[3296], Cout[3296]);
	Full_Adder FA3238 (S[2457], Cout[2923], Cout[2924], S[3297], Cout[3297]);
	Full_Adder FA3239 (Cout[2925], Cout[2926], S[2927], S[3298], Cout[3298]);
	Full_Adder FA3240 (S[2928], S[2929], S[2930], S[3299], Cout[3299]);
	Full_Adder FA3241 (S[2463], Cout[2927], Cout[2928], S[3300], Cout[3300]);
	Full_Adder FA3242 (Cout[2929], Cout[2930], S[2931], S[3301], Cout[3301]);
	Full_Adder FA3243 (S[2932], S[2933], S[2934], S[3302], Cout[3302]);
	Full_Adder FA3244 (S[2469], Cout[2931], Cout[2932], S[3303], Cout[3303]);
	Full_Adder FA3245 (Cout[2933], Cout[2934], S[2935], S[3304], Cout[3304]);
	Full_Adder FA3246 (S[2936], S[2937], S[2938], S[3305], Cout[3305]);
	Full_Adder FA3247 (S[2475], Cout[2935], Cout[2936], S[3306], Cout[3306]);
	Full_Adder FA3248 (Cout[2937], Cout[2938], S[2939], S[3307], Cout[3307]);
	Full_Adder FA3249 (S[2940], S[2941], S[2942], S[3308], Cout[3308]);
	Full_Adder FA3250 (S[2481], Cout[2939], Cout[2940], S[3309], Cout[3309]);
	Full_Adder FA3251 (Cout[2941], Cout[2942], S[2943], S[3310], Cout[3310]);
	Full_Adder FA3252 (S[2944], S[2945], S[2946], S[3311], Cout[3311]);
	Full_Adder FA3253 (S[2487], Cout[2943], Cout[2944], S[3312], Cout[3312]);
	Full_Adder FA3254 (Cout[2945], Cout[2946], S[2947], S[3313], Cout[3313]);
	Full_Adder FA3255 (S[2948], S[2949], S[2950], S[3314], Cout[3314]);
	Full_Adder FA3256 (S[2493], Cout[2947], Cout[2948], S[3315], Cout[3315]);
	Full_Adder FA3257 (Cout[2949], Cout[2950], S[2951], S[3316], Cout[3316]);
	Full_Adder FA3258 (S[2952], S[2953], S[2954], S[3317], Cout[3317]);
	Full_Adder FA3259 (S[2499], Cout[2951], Cout[2952], S[3318], Cout[3318]);
	Full_Adder FA3260 (Cout[2953], Cout[2954], S[2955], S[3319], Cout[3319]);
	Full_Adder FA3261 (S[2956], S[2957], S[2958], S[3320], Cout[3320]);
	Full_Adder FA3262 (S[2505], Cout[2955], Cout[2956], S[3321], Cout[3321]);
	Full_Adder FA3263 (Cout[2957], Cout[2958], S[2959], S[3322], Cout[3322]);
	Full_Adder FA3264 (S[2960], S[2961], S[2962], S[3323], Cout[3323]);
	Full_Adder FA3265 (S[2511], Cout[2959], Cout[2960], S[3324], Cout[3324]);
	Full_Adder FA3266 (Cout[2961], Cout[2962], S[2963], S[3325], Cout[3325]);
	Full_Adder FA3267 (S[2964], S[2965], S[2966], S[3326], Cout[3326]);
	Full_Adder FA3268 (S[2517], Cout[2963], Cout[2964], S[3327], Cout[3327]);
	Full_Adder FA3269 (Cout[2965], Cout[2966], S[2967], S[3328], Cout[3328]);
	Full_Adder FA3270 (S[2968], S[2969], S[2970], S[3329], Cout[3329]);
	Full_Adder FA3271 (S[2523], Cout[2967], Cout[2968], S[3330], Cout[3330]);
	Full_Adder FA3272 (Cout[2969], Cout[2970], S[2971], S[3331], Cout[3331]);
	Full_Adder FA3273 (S[2972], S[2973], S[2974], S[3332], Cout[3332]);
	Full_Adder FA3274 (S[2529], Cout[2971], Cout[2972], S[3333], Cout[3333]);
	Full_Adder FA3275 (Cout[2973], Cout[2974], S[2975], S[3334], Cout[3334]);
	Full_Adder FA3276 (S[2976], S[2977], S[2978], S[3335], Cout[3335]);
	Full_Adder FA3277 (S[2535], Cout[2975], Cout[2976], S[3336], Cout[3336]);
	Full_Adder FA3278 (Cout[2977], Cout[2978], S[2979], S[3337], Cout[3337]);
	Full_Adder FA3279 (S[2980], S[2981], S[2982], S[3338], Cout[3338]);
	Full_Adder FA3280 (S[2541], Cout[2979], Cout[2980], S[3339], Cout[3339]);
	Full_Adder FA3281 (Cout[2981], Cout[2982], S[2983], S[3340], Cout[3340]);
	Full_Adder FA3282 (S[2984], S[2985], S[2986], S[3341], Cout[3341]);
	Full_Adder FA3283 (S[2547], Cout[2983], Cout[2984], S[3342], Cout[3342]);
	Full_Adder FA3284 (Cout[2985], Cout[2986], S[2987], S[3343], Cout[3343]);
	Full_Adder FA3285 (S[2988], S[2989], S[2990], S[3344], Cout[3344]);
	Full_Adder FA3286 (S[2553], Cout[2987], Cout[2988], S[3345], Cout[3345]);
	Full_Adder FA3287 (Cout[2989], Cout[2990], S[2991], S[3346], Cout[3346]);
	Full_Adder FA3288 (S[2992], S[2993], S[2994], S[3347], Cout[3347]);
	Full_Adder FA3289 (S[2559], Cout[2991], Cout[2992], S[3348], Cout[3348]);
	Full_Adder FA3290 (Cout[2993], Cout[2994], S[2995], S[3349], Cout[3349]);
	Full_Adder FA3291 (S[2996], S[2997], S[2998], S[3350], Cout[3350]);
	Full_Adder FA3292 (S[2565], Cout[2995], Cout[2996], S[3351], Cout[3351]);
	Full_Adder FA3293 (Cout[2997], Cout[2998], S[2999], S[3352], Cout[3352]);
	Full_Adder FA3294 (S[3000], S[3001], S[3002], S[3353], Cout[3353]);
	Full_Adder FA3295 (S[2571], Cout[2999], Cout[3000], S[3354], Cout[3354]);
	Full_Adder FA3296 (Cout[3001], Cout[3002], S[3003], S[3355], Cout[3355]);
	Full_Adder FA3297 (S[3004], S[3005], S[3006], S[3356], Cout[3356]);
	Full_Adder FA3298 (S[2577], Cout[3003], Cout[3004], S[3357], Cout[3357]);
	Full_Adder FA3299 (Cout[3005], Cout[3006], S[3007], S[3358], Cout[3358]);
	Full_Adder FA3300 (S[3008], S[3009], S[3010], S[3359], Cout[3359]);
	Full_Adder FA3301 (S[2583], Cout[3007], Cout[3008], S[3360], Cout[3360]);
	Full_Adder FA3302 (Cout[3009], Cout[3010], S[3011], S[3361], Cout[3361]);
	Full_Adder FA3303 (S[3012], S[3013], S[3014], S[3362], Cout[3362]);
	Full_Adder FA3304 (S[2589], Cout[3011], Cout[3012], S[3363], Cout[3363]);
	Full_Adder FA3305 (Cout[3013], Cout[3014], S[3015], S[3364], Cout[3364]);
	Full_Adder FA3306 (S[3016], S[3017], S[3018], S[3365], Cout[3365]);
	Full_Adder FA3307 (S[2595], Cout[3015], Cout[3016], S[3366], Cout[3366]);
	Full_Adder FA3308 (Cout[3017], Cout[3018], S[3019], S[3367], Cout[3367]);
	Full_Adder FA3309 (S[3020], S[3021], S[3022], S[3368], Cout[3368]);
	Full_Adder FA3310 (S[2601], Cout[3019], Cout[3020], S[3369], Cout[3369]);
	Full_Adder FA3311 (Cout[3021], Cout[3022], S[3023], S[3370], Cout[3370]);
	Full_Adder FA3312 (S[3024], S[3025], S[3026], S[3371], Cout[3371]);
	Full_Adder FA3313 (S[2607], Cout[3023], Cout[3024], S[3372], Cout[3372]);
	Full_Adder FA3314 (Cout[3025], Cout[3026], S[3027], S[3373], Cout[3373]);
	Full_Adder FA3315 (S[3028], S[3029], S[3030], S[3374], Cout[3374]);
	Full_Adder FA3316 (S[2613], Cout[3027], Cout[3028], S[3375], Cout[3375]);
	Full_Adder FA3317 (Cout[3029], Cout[3030], S[3031], S[3376], Cout[3376]);
	Full_Adder FA3318 (S[3032], S[3033], S[3034], S[3377], Cout[3377]);
	Full_Adder FA3319 (S[2619], Cout[3031], Cout[3032], S[3378], Cout[3378]);
	Full_Adder FA3320 (Cout[3033], Cout[3034], S[3035], S[3379], Cout[3379]);
	Full_Adder FA3321 (S[3036], S[3037], S[3038], S[3380], Cout[3380]);
	Full_Adder FA3322 (S[2625], Cout[3035], Cout[3036], S[3381], Cout[3381]);
	Full_Adder FA3323 (Cout[3037], Cout[3038], S[3039], S[3382], Cout[3382]);
	Full_Adder FA3324 (S[3040], S[3041], S[3042], S[3383], Cout[3383]);
	Full_Adder FA3325 (S[2631], Cout[3039], Cout[3040], S[3384], Cout[3384]);
	Full_Adder FA3326 (Cout[3041], Cout[3042], S[3043], S[3385], Cout[3385]);
	Full_Adder FA3327 (S[3044], S[3045], S[3046], S[3386], Cout[3386]);
	Full_Adder FA3328 (S[2637], Cout[3043], Cout[3044], S[3387], Cout[3387]);
	Full_Adder FA3329 (Cout[3045], Cout[3046], S[3047], S[3388], Cout[3388]);
	Full_Adder FA3330 (S[3048], S[3049], S[3050], S[3389], Cout[3389]);
	Full_Adder FA3331 (S[2642], Cout[3047], Cout[3048], S[3390], Cout[3390]);
	Full_Adder FA3332 (Cout[3049], Cout[3050], S[3051], S[3391], Cout[3391]);
	Full_Adder FA3333 (S[3052], S[3053], S[3054], S[3392], Cout[3392]);
	Full_Adder FA3334 (S[2646], Cout[3051], Cout[3052], S[3393], Cout[3393]);
	Full_Adder FA3335 (Cout[3053], Cout[3054], S[3055], S[3394], Cout[3394]);
	Full_Adder FA3336 (S[3056], S[3057], S[3058], S[3395], Cout[3395]);
	Full_Adder FA3337 (S[2649], Cout[3055], Cout[3056], S[3396], Cout[3396]);
	Full_Adder FA3338 (Cout[3057], Cout[3058], S[3059], S[3397], Cout[3397]);
	Full_Adder FA3339 (S[3060], S[3061], S[3062], S[3398], Cout[3398]);
	Full_Adder FA3340 (S[2651], Cout[3059], Cout[3060], S[3399], Cout[3399]);
	Full_Adder FA3341 (Cout[3061], Cout[3062], S[3063], S[3400], Cout[3400]);
	Full_Adder FA3342 (S[3064], S[3065], S[3066], S[3401], Cout[3401]);
	Full_Adder FA3343 (S[2652], Cout[3063], Cout[3064], S[3402], Cout[3402]);
	Full_Adder FA3344 (Cout[3065], Cout[3066], S[3067], S[3403], Cout[3403]);
	Full_Adder FA3345 (S[3068], S[3069], S[3070], S[3404], Cout[3404]);
	Full_Adder FA3346 (Cout[2652], Cout[3067], Cout[3068], S[3405], Cout[3405]);
	Full_Adder FA3347 (Cout[3069], Cout[3070], S[3071], S[3406], Cout[3406]);
	Full_Adder FA3348 (S[3072], S[3073], S[3074], S[3407], Cout[3407]);
	Full_Adder FA3349 (pp62[54], pp63[53], Cout[3071], S[3408], Cout[3408]);
	Full_Adder FA3350 (Cout[3072], Cout[3073], Cout[3074], S[3409], Cout[3409]);
	Full_Adder FA3351 (S[3075], S[3076], S[3077], S[3410], Cout[3410]);
	Full_Adder FA3352 (pp60[57], pp61[56], pp62[55], S[3411], Cout[3411]);
	Full_Adder FA3353 (pp63[54], Cout[3075], Cout[3076], S[3412], Cout[3412]);
	Full_Adder FA3354 (Cout[3077], S[3078], S[3079], S[3413], Cout[3413]);
	Full_Adder FA3355 (pp58[60], pp59[59], pp60[58], S[3414], Cout[3414]);
	Full_Adder FA3356 (pp61[57], pp62[56], pp63[55], S[3415], Cout[3415]);
	Full_Adder FA3357 (Cout[3078], Cout[3079], S[3080], S[3416], Cout[3416]);
	Full_Adder FA3358 (pp56[63], pp57[62], pp58[61], S[3417], Cout[3417]);
	Full_Adder FA3359 (pp59[60], pp60[59], pp61[58], S[3418], Cout[3418]);
	Full_Adder FA3360 (pp62[57], pp63[56], Cout[3080], S[3419], Cout[3419]);
	Full_Adder FA3361 (pp57[63], pp58[62], pp59[61], S[3420], Cout[3420]);
	Full_Adder FA3362 (pp60[60], pp61[59], pp62[58], S[3421], Cout[3421]);
	Full_Adder FA3363 (pp58[63], pp59[62], pp60[61], S[3422], Cout[3422]);
	Half_Adder HA60 (pp0[4], pp1[3], S[3423], Cout[3423]);
	Full_Adder FA3364 (pp0[5], pp1[4], pp2[3], S[3424], Cout[3424]);
	Half_Adder HA61 (pp3[2], pp4[1], S[3425], Cout[3425]);
	Full_Adder FA3365 (pp2[4], pp3[3], pp4[2], S[3426], Cout[3426]);
	Full_Adder FA3366 (pp5[1], pp6[0], S[3081], S[3427], Cout[3427]);
	Full_Adder FA3367 (pp5[2], pp6[1], pp7[0], S[3428], Cout[3428]);
	Full_Adder FA3368 (Cout[3081], S[3082], S[3083], S[3429], Cout[3429]);
	Full_Adder FA3369 (pp8[0], Cout[3082], Cout[3083], S[3430], Cout[3430]);
	Full_Adder FA3370 (S[3084], S[3085], S[3086], S[3431], Cout[3431]);
	Full_Adder FA3371 (Cout[3084], Cout[3085], Cout[3086], S[3432], Cout[3432]);
	Full_Adder FA3372 (S[3087], S[3088], S[3089], S[3433], Cout[3433]);
	Full_Adder FA3373 (Cout[3087], Cout[3088], Cout[3089], S[3434], Cout[3434]);
	Full_Adder FA3374 (S[3090], S[3091], S[3092], S[3435], Cout[3435]);
	Full_Adder FA3375 (Cout[3090], Cout[3091], Cout[3092], S[3436], Cout[3436]);
	Full_Adder FA3376 (S[3093], S[3094], S[3095], S[3437], Cout[3437]);
	Full_Adder FA3377 (Cout[3093], Cout[3094], Cout[3095], S[3438], Cout[3438]);
	Full_Adder FA3378 (S[3096], S[3097], S[3098], S[3439], Cout[3439]);
	Full_Adder FA3379 (Cout[3096], Cout[3097], Cout[3098], S[3440], Cout[3440]);
	Full_Adder FA3380 (S[3099], S[3100], S[3101], S[3441], Cout[3441]);
	Full_Adder FA3381 (Cout[3099], Cout[3100], Cout[3101], S[3442], Cout[3442]);
	Full_Adder FA3382 (S[3102], S[3103], S[3104], S[3443], Cout[3443]);
	Full_Adder FA3383 (Cout[3102], Cout[3103], Cout[3104], S[3444], Cout[3444]);
	Full_Adder FA3384 (S[3105], S[3106], S[3107], S[3445], Cout[3445]);
	Full_Adder FA3385 (Cout[3105], Cout[3106], Cout[3107], S[3446], Cout[3446]);
	Full_Adder FA3386 (S[3108], S[3109], S[3110], S[3447], Cout[3447]);
	Full_Adder FA3387 (Cout[3108], Cout[3109], Cout[3110], S[3448], Cout[3448]);
	Full_Adder FA3388 (S[3111], S[3112], S[3113], S[3449], Cout[3449]);
	Full_Adder FA3389 (Cout[3111], Cout[3112], Cout[3113], S[3450], Cout[3450]);
	Full_Adder FA3390 (S[3114], S[3115], S[3116], S[3451], Cout[3451]);
	Full_Adder FA3391 (Cout[3114], Cout[3115], Cout[3116], S[3452], Cout[3452]);
	Full_Adder FA3392 (S[3117], S[3118], S[3119], S[3453], Cout[3453]);
	Full_Adder FA3393 (Cout[3117], Cout[3118], Cout[3119], S[3454], Cout[3454]);
	Full_Adder FA3394 (S[3120], S[3121], S[3122], S[3455], Cout[3455]);
	Full_Adder FA3395 (Cout[3120], Cout[3121], Cout[3122], S[3456], Cout[3456]);
	Full_Adder FA3396 (S[3123], S[3124], S[3125], S[3457], Cout[3457]);
	Full_Adder FA3397 (Cout[3123], Cout[3124], Cout[3125], S[3458], Cout[3458]);
	Full_Adder FA3398 (S[3126], S[3127], S[3128], S[3459], Cout[3459]);
	Full_Adder FA3399 (Cout[3126], Cout[3127], Cout[3128], S[3460], Cout[3460]);
	Full_Adder FA3400 (S[3129], S[3130], S[3131], S[3461], Cout[3461]);
	Full_Adder FA3401 (Cout[3129], Cout[3130], Cout[3131], S[3462], Cout[3462]);
	Full_Adder FA3402 (S[3132], S[3133], S[3134], S[3463], Cout[3463]);
	Full_Adder FA3403 (Cout[3132], Cout[3133], Cout[3134], S[3464], Cout[3464]);
	Full_Adder FA3404 (S[3135], S[3136], S[3137], S[3465], Cout[3465]);
	Full_Adder FA3405 (Cout[3135], Cout[3136], Cout[3137], S[3466], Cout[3466]);
	Full_Adder FA3406 (S[3138], S[3139], S[3140], S[3467], Cout[3467]);
	Full_Adder FA3407 (Cout[3138], Cout[3139], Cout[3140], S[3468], Cout[3468]);
	Full_Adder FA3408 (S[3141], S[3142], S[3143], S[3469], Cout[3469]);
	Full_Adder FA3409 (Cout[3141], Cout[3142], Cout[3143], S[3470], Cout[3470]);
	Full_Adder FA3410 (S[3144], S[3145], S[3146], S[3471], Cout[3471]);
	Full_Adder FA3411 (Cout[3144], Cout[3145], Cout[3146], S[3472], Cout[3472]);
	Full_Adder FA3412 (S[3147], S[3148], S[3149], S[3473], Cout[3473]);
	Full_Adder FA3413 (Cout[3147], Cout[3148], Cout[3149], S[3474], Cout[3474]);
	Full_Adder FA3414 (S[3150], S[3151], S[3152], S[3475], Cout[3475]);
	Full_Adder FA3415 (Cout[3150], Cout[3151], Cout[3152], S[3476], Cout[3476]);
	Full_Adder FA3416 (S[3153], S[3154], S[3155], S[3477], Cout[3477]);
	Full_Adder FA3417 (Cout[3153], Cout[3154], Cout[3155], S[3478], Cout[3478]);
	Full_Adder FA3418 (S[3156], S[3157], S[3158], S[3479], Cout[3479]);
	Full_Adder FA3419 (Cout[3156], Cout[3157], Cout[3158], S[3480], Cout[3480]);
	Full_Adder FA3420 (S[3159], S[3160], S[3161], S[3481], Cout[3481]);
	Full_Adder FA3421 (Cout[3159], Cout[3160], Cout[3161], S[3482], Cout[3482]);
	Full_Adder FA3422 (S[3162], S[3163], S[3164], S[3483], Cout[3483]);
	Full_Adder FA3423 (Cout[3162], Cout[3163], Cout[3164], S[3484], Cout[3484]);
	Full_Adder FA3424 (S[3165], S[3166], S[3167], S[3485], Cout[3485]);
	Full_Adder FA3425 (Cout[3165], Cout[3166], Cout[3167], S[3486], Cout[3486]);
	Full_Adder FA3426 (S[3168], S[3169], S[3170], S[3487], Cout[3487]);
	Full_Adder FA3427 (Cout[3168], Cout[3169], Cout[3170], S[3488], Cout[3488]);
	Full_Adder FA3428 (S[3171], S[3172], S[3173], S[3489], Cout[3489]);
	Full_Adder FA3429 (Cout[3171], Cout[3172], Cout[3173], S[3490], Cout[3490]);
	Full_Adder FA3430 (S[3174], S[3175], S[3176], S[3491], Cout[3491]);
	Full_Adder FA3431 (Cout[3174], Cout[3175], Cout[3176], S[3492], Cout[3492]);
	Full_Adder FA3432 (S[3177], S[3178], S[3179], S[3493], Cout[3493]);
	Full_Adder FA3433 (Cout[3177], Cout[3178], Cout[3179], S[3494], Cout[3494]);
	Full_Adder FA3434 (S[3180], S[3181], S[3182], S[3495], Cout[3495]);
	Full_Adder FA3435 (Cout[3180], Cout[3181], Cout[3182], S[3496], Cout[3496]);
	Full_Adder FA3436 (S[3183], S[3184], S[3185], S[3497], Cout[3497]);
	Full_Adder FA3437 (Cout[3183], Cout[3184], Cout[3185], S[3498], Cout[3498]);
	Full_Adder FA3438 (S[3186], S[3187], S[3188], S[3499], Cout[3499]);
	Full_Adder FA3439 (Cout[3186], Cout[3187], Cout[3188], S[3500], Cout[3500]);
	Full_Adder FA3440 (S[3189], S[3190], S[3191], S[3501], Cout[3501]);
	Full_Adder FA3441 (Cout[3189], Cout[3190], Cout[3191], S[3502], Cout[3502]);
	Full_Adder FA3442 (S[3192], S[3193], S[3194], S[3503], Cout[3503]);
	Full_Adder FA3443 (Cout[3192], Cout[3193], Cout[3194], S[3504], Cout[3504]);
	Full_Adder FA3444 (S[3195], S[3196], S[3197], S[3505], Cout[3505]);
	Full_Adder FA3445 (Cout[3195], Cout[3196], Cout[3197], S[3506], Cout[3506]);
	Full_Adder FA3446 (S[3198], S[3199], S[3200], S[3507], Cout[3507]);
	Full_Adder FA3447 (Cout[3198], Cout[3199], Cout[3200], S[3508], Cout[3508]);
	Full_Adder FA3448 (S[3201], S[3202], S[3203], S[3509], Cout[3509]);
	Full_Adder FA3449 (Cout[3201], Cout[3202], Cout[3203], S[3510], Cout[3510]);
	Full_Adder FA3450 (S[3204], S[3205], S[3206], S[3511], Cout[3511]);
	Full_Adder FA3451 (Cout[3204], Cout[3205], Cout[3206], S[3512], Cout[3512]);
	Full_Adder FA3452 (S[3207], S[3208], S[3209], S[3513], Cout[3513]);
	Full_Adder FA3453 (Cout[3207], Cout[3208], Cout[3209], S[3514], Cout[3514]);
	Full_Adder FA3454 (S[3210], S[3211], S[3212], S[3515], Cout[3515]);
	Full_Adder FA3455 (Cout[3210], Cout[3211], Cout[3212], S[3516], Cout[3516]);
	Full_Adder FA3456 (S[3213], S[3214], S[3215], S[3517], Cout[3517]);
	Full_Adder FA3457 (Cout[3213], Cout[3214], Cout[3215], S[3518], Cout[3518]);
	Full_Adder FA3458 (S[3216], S[3217], S[3218], S[3519], Cout[3519]);
	Full_Adder FA3459 (Cout[3216], Cout[3217], Cout[3218], S[3520], Cout[3520]);
	Full_Adder FA3460 (S[3219], S[3220], S[3221], S[3521], Cout[3521]);
	Full_Adder FA3461 (Cout[3219], Cout[3220], Cout[3221], S[3522], Cout[3522]);
	Full_Adder FA3462 (S[3222], S[3223], S[3224], S[3523], Cout[3523]);
	Full_Adder FA3463 (Cout[3222], Cout[3223], Cout[3224], S[3524], Cout[3524]);
	Full_Adder FA3464 (S[3225], S[3226], S[3227], S[3525], Cout[3525]);
	Full_Adder FA3465 (Cout[3225], Cout[3226], Cout[3227], S[3526], Cout[3526]);
	Full_Adder FA3466 (S[3228], S[3229], S[3230], S[3527], Cout[3527]);
	Full_Adder FA3467 (Cout[3228], Cout[3229], Cout[3230], S[3528], Cout[3528]);
	Full_Adder FA3468 (S[3231], S[3232], S[3233], S[3529], Cout[3529]);
	Full_Adder FA3469 (Cout[3231], Cout[3232], Cout[3233], S[3530], Cout[3530]);
	Full_Adder FA3470 (S[3234], S[3235], S[3236], S[3531], Cout[3531]);
	Full_Adder FA3471 (Cout[3234], Cout[3235], Cout[3236], S[3532], Cout[3532]);
	Full_Adder FA3472 (S[3237], S[3238], S[3239], S[3533], Cout[3533]);
	Full_Adder FA3473 (Cout[3237], Cout[3238], Cout[3239], S[3534], Cout[3534]);
	Full_Adder FA3474 (S[3240], S[3241], S[3242], S[3535], Cout[3535]);
	Full_Adder FA3475 (Cout[3240], Cout[3241], Cout[3242], S[3536], Cout[3536]);
	Full_Adder FA3476 (S[3243], S[3244], S[3245], S[3537], Cout[3537]);
	Full_Adder FA3477 (Cout[3243], Cout[3244], Cout[3245], S[3538], Cout[3538]);
	Full_Adder FA3478 (S[3246], S[3247], S[3248], S[3539], Cout[3539]);
	Full_Adder FA3479 (Cout[3246], Cout[3247], Cout[3248], S[3540], Cout[3540]);
	Full_Adder FA3480 (S[3249], S[3250], S[3251], S[3541], Cout[3541]);
	Full_Adder FA3481 (Cout[3249], Cout[3250], Cout[3251], S[3542], Cout[3542]);
	Full_Adder FA3482 (S[3252], S[3253], S[3254], S[3543], Cout[3543]);
	Full_Adder FA3483 (Cout[3252], Cout[3253], Cout[3254], S[3544], Cout[3544]);
	Full_Adder FA3484 (S[3255], S[3256], S[3257], S[3545], Cout[3545]);
	Full_Adder FA3485 (Cout[3255], Cout[3256], Cout[3257], S[3546], Cout[3546]);
	Full_Adder FA3486 (S[3258], S[3259], S[3260], S[3547], Cout[3547]);
	Full_Adder FA3487 (Cout[3258], Cout[3259], Cout[3260], S[3548], Cout[3548]);
	Full_Adder FA3488 (S[3261], S[3262], S[3263], S[3549], Cout[3549]);
	Full_Adder FA3489 (Cout[3261], Cout[3262], Cout[3263], S[3550], Cout[3550]);
	Full_Adder FA3490 (S[3264], S[3265], S[3266], S[3551], Cout[3551]);
	Full_Adder FA3491 (Cout[3264], Cout[3265], Cout[3266], S[3552], Cout[3552]);
	Full_Adder FA3492 (S[3267], S[3268], S[3269], S[3553], Cout[3553]);
	Full_Adder FA3493 (Cout[3267], Cout[3268], Cout[3269], S[3554], Cout[3554]);
	Full_Adder FA3494 (S[3270], S[3271], S[3272], S[3555], Cout[3555]);
	Full_Adder FA3495 (Cout[3270], Cout[3271], Cout[3272], S[3556], Cout[3556]);
	Full_Adder FA3496 (S[3273], S[3274], S[3275], S[3557], Cout[3557]);
	Full_Adder FA3497 (Cout[3273], Cout[3274], Cout[3275], S[3558], Cout[3558]);
	Full_Adder FA3498 (S[3276], S[3277], S[3278], S[3559], Cout[3559]);
	Full_Adder FA3499 (Cout[3276], Cout[3277], Cout[3278], S[3560], Cout[3560]);
	Full_Adder FA3500 (S[3279], S[3280], S[3281], S[3561], Cout[3561]);
	Full_Adder FA3501 (Cout[3279], Cout[3280], Cout[3281], S[3562], Cout[3562]);
	Full_Adder FA3502 (S[3282], S[3283], S[3284], S[3563], Cout[3563]);
	Full_Adder FA3503 (Cout[3282], Cout[3283], Cout[3284], S[3564], Cout[3564]);
	Full_Adder FA3504 (S[3285], S[3286], S[3287], S[3565], Cout[3565]);
	Full_Adder FA3505 (Cout[3285], Cout[3286], Cout[3287], S[3566], Cout[3566]);
	Full_Adder FA3506 (S[3288], S[3289], S[3290], S[3567], Cout[3567]);
	Full_Adder FA3507 (Cout[3288], Cout[3289], Cout[3290], S[3568], Cout[3568]);
	Full_Adder FA3508 (S[3291], S[3292], S[3293], S[3569], Cout[3569]);
	Full_Adder FA3509 (Cout[3291], Cout[3292], Cout[3293], S[3570], Cout[3570]);
	Full_Adder FA3510 (S[3294], S[3295], S[3296], S[3571], Cout[3571]);
	Full_Adder FA3511 (Cout[3294], Cout[3295], Cout[3296], S[3572], Cout[3572]);
	Full_Adder FA3512 (S[3297], S[3298], S[3299], S[3573], Cout[3573]);
	Full_Adder FA3513 (Cout[3297], Cout[3298], Cout[3299], S[3574], Cout[3574]);
	Full_Adder FA3514 (S[3300], S[3301], S[3302], S[3575], Cout[3575]);
	Full_Adder FA3515 (Cout[3300], Cout[3301], Cout[3302], S[3576], Cout[3576]);
	Full_Adder FA3516 (S[3303], S[3304], S[3305], S[3577], Cout[3577]);
	Full_Adder FA3517 (Cout[3303], Cout[3304], Cout[3305], S[3578], Cout[3578]);
	Full_Adder FA3518 (S[3306], S[3307], S[3308], S[3579], Cout[3579]);
	Full_Adder FA3519 (Cout[3306], Cout[3307], Cout[3308], S[3580], Cout[3580]);
	Full_Adder FA3520 (S[3309], S[3310], S[3311], S[3581], Cout[3581]);
	Full_Adder FA3521 (Cout[3309], Cout[3310], Cout[3311], S[3582], Cout[3582]);
	Full_Adder FA3522 (S[3312], S[3313], S[3314], S[3583], Cout[3583]);
	Full_Adder FA3523 (Cout[3312], Cout[3313], Cout[3314], S[3584], Cout[3584]);
	Full_Adder FA3524 (S[3315], S[3316], S[3317], S[3585], Cout[3585]);
	Full_Adder FA3525 (Cout[3315], Cout[3316], Cout[3317], S[3586], Cout[3586]);
	Full_Adder FA3526 (S[3318], S[3319], S[3320], S[3587], Cout[3587]);
	Full_Adder FA3527 (Cout[3318], Cout[3319], Cout[3320], S[3588], Cout[3588]);
	Full_Adder FA3528 (S[3321], S[3322], S[3323], S[3589], Cout[3589]);
	Full_Adder FA3529 (Cout[3321], Cout[3322], Cout[3323], S[3590], Cout[3590]);
	Full_Adder FA3530 (S[3324], S[3325], S[3326], S[3591], Cout[3591]);
	Full_Adder FA3531 (Cout[3324], Cout[3325], Cout[3326], S[3592], Cout[3592]);
	Full_Adder FA3532 (S[3327], S[3328], S[3329], S[3593], Cout[3593]);
	Full_Adder FA3533 (Cout[3327], Cout[3328], Cout[3329], S[3594], Cout[3594]);
	Full_Adder FA3534 (S[3330], S[3331], S[3332], S[3595], Cout[3595]);
	Full_Adder FA3535 (Cout[3330], Cout[3331], Cout[3332], S[3596], Cout[3596]);
	Full_Adder FA3536 (S[3333], S[3334], S[3335], S[3597], Cout[3597]);
	Full_Adder FA3537 (Cout[3333], Cout[3334], Cout[3335], S[3598], Cout[3598]);
	Full_Adder FA3538 (S[3336], S[3337], S[3338], S[3599], Cout[3599]);
	Full_Adder FA3539 (Cout[3336], Cout[3337], Cout[3338], S[3600], Cout[3600]);
	Full_Adder FA3540 (S[3339], S[3340], S[3341], S[3601], Cout[3601]);
	Full_Adder FA3541 (Cout[3339], Cout[3340], Cout[3341], S[3602], Cout[3602]);
	Full_Adder FA3542 (S[3342], S[3343], S[3344], S[3603], Cout[3603]);
	Full_Adder FA3543 (Cout[3342], Cout[3343], Cout[3344], S[3604], Cout[3604]);
	Full_Adder FA3544 (S[3345], S[3346], S[3347], S[3605], Cout[3605]);
	Full_Adder FA3545 (Cout[3345], Cout[3346], Cout[3347], S[3606], Cout[3606]);
	Full_Adder FA3546 (S[3348], S[3349], S[3350], S[3607], Cout[3607]);
	Full_Adder FA3547 (Cout[3348], Cout[3349], Cout[3350], S[3608], Cout[3608]);
	Full_Adder FA3548 (S[3351], S[3352], S[3353], S[3609], Cout[3609]);
	Full_Adder FA3549 (Cout[3351], Cout[3352], Cout[3353], S[3610], Cout[3610]);
	Full_Adder FA3550 (S[3354], S[3355], S[3356], S[3611], Cout[3611]);
	Full_Adder FA3551 (Cout[3354], Cout[3355], Cout[3356], S[3612], Cout[3612]);
	Full_Adder FA3552 (S[3357], S[3358], S[3359], S[3613], Cout[3613]);
	Full_Adder FA3553 (Cout[3357], Cout[3358], Cout[3359], S[3614], Cout[3614]);
	Full_Adder FA3554 (S[3360], S[3361], S[3362], S[3615], Cout[3615]);
	Full_Adder FA3555 (Cout[3360], Cout[3361], Cout[3362], S[3616], Cout[3616]);
	Full_Adder FA3556 (S[3363], S[3364], S[3365], S[3617], Cout[3617]);
	Full_Adder FA3557 (Cout[3363], Cout[3364], Cout[3365], S[3618], Cout[3618]);
	Full_Adder FA3558 (S[3366], S[3367], S[3368], S[3619], Cout[3619]);
	Full_Adder FA3559 (Cout[3366], Cout[3367], Cout[3368], S[3620], Cout[3620]);
	Full_Adder FA3560 (S[3369], S[3370], S[3371], S[3621], Cout[3621]);
	Full_Adder FA3561 (Cout[3369], Cout[3370], Cout[3371], S[3622], Cout[3622]);
	Full_Adder FA3562 (S[3372], S[3373], S[3374], S[3623], Cout[3623]);
	Full_Adder FA3563 (Cout[3372], Cout[3373], Cout[3374], S[3624], Cout[3624]);
	Full_Adder FA3564 (S[3375], S[3376], S[3377], S[3625], Cout[3625]);
	Full_Adder FA3565 (Cout[3375], Cout[3376], Cout[3377], S[3626], Cout[3626]);
	Full_Adder FA3566 (S[3378], S[3379], S[3380], S[3627], Cout[3627]);
	Full_Adder FA3567 (Cout[3378], Cout[3379], Cout[3380], S[3628], Cout[3628]);
	Full_Adder FA3568 (S[3381], S[3382], S[3383], S[3629], Cout[3629]);
	Full_Adder FA3569 (Cout[3381], Cout[3382], Cout[3383], S[3630], Cout[3630]);
	Full_Adder FA3570 (S[3384], S[3385], S[3386], S[3631], Cout[3631]);
	Full_Adder FA3571 (Cout[3384], Cout[3385], Cout[3386], S[3632], Cout[3632]);
	Full_Adder FA3572 (S[3387], S[3388], S[3389], S[3633], Cout[3633]);
	Full_Adder FA3573 (Cout[3387], Cout[3388], Cout[3389], S[3634], Cout[3634]);
	Full_Adder FA3574 (S[3390], S[3391], S[3392], S[3635], Cout[3635]);
	Full_Adder FA3575 (Cout[3390], Cout[3391], Cout[3392], S[3636], Cout[3636]);
	Full_Adder FA3576 (S[3393], S[3394], S[3395], S[3637], Cout[3637]);
	Full_Adder FA3577 (Cout[3393], Cout[3394], Cout[3395], S[3638], Cout[3638]);
	Full_Adder FA3578 (S[3396], S[3397], S[3398], S[3639], Cout[3639]);
	Full_Adder FA3579 (Cout[3396], Cout[3397], Cout[3398], S[3640], Cout[3640]);
	Full_Adder FA3580 (S[3399], S[3400], S[3401], S[3641], Cout[3641]);
	Full_Adder FA3581 (Cout[3399], Cout[3400], Cout[3401], S[3642], Cout[3642]);
	Full_Adder FA3582 (S[3402], S[3403], S[3404], S[3643], Cout[3643]);
	Full_Adder FA3583 (Cout[3402], Cout[3403], Cout[3404], S[3644], Cout[3644]);
	Full_Adder FA3584 (S[3405], S[3406], S[3407], S[3645], Cout[3645]);
	Full_Adder FA3585 (Cout[3405], Cout[3406], Cout[3407], S[3646], Cout[3646]);
	Full_Adder FA3586 (S[3408], S[3409], S[3410], S[3647], Cout[3647]);
	Full_Adder FA3587 (Cout[3408], Cout[3409], Cout[3410], S[3648], Cout[3648]);
	Full_Adder FA3588 (S[3411], S[3412], S[3413], S[3649], Cout[3649]);
	Full_Adder FA3589 (Cout[3411], Cout[3412], Cout[3413], S[3650], Cout[3650]);
	Full_Adder FA3590 (S[3414], S[3415], S[3416], S[3651], Cout[3651]);
	Full_Adder FA3591 (Cout[3414], Cout[3415], Cout[3416], S[3652], Cout[3652]);
	Full_Adder FA3592 (S[3417], S[3418], S[3419], S[3653], Cout[3653]);
	Full_Adder FA3593 (pp63[57], Cout[3417], Cout[3418], S[3654], Cout[3654]);
	Full_Adder FA3594 (Cout[3419], S[3420], S[3421], S[3655], Cout[3655]);
	Full_Adder FA3595 (pp61[60], pp62[59], pp63[58], S[3656], Cout[3656]);
	Full_Adder FA3596 (Cout[3420], Cout[3421], S[3422], S[3657], Cout[3657]);
	Full_Adder FA3597 (pp59[63], pp60[62], pp61[61], S[3658], Cout[3658]);
	Full_Adder FA3598 (pp62[60], pp63[59], Cout[3422], S[3659], Cout[3659]);
	Full_Adder FA3599 (pp60[63], pp61[62], pp62[61], S[3660], Cout[3660]);
	Half_Adder HA62 (pp0[3], pp1[2], S[3661], Cout[3661]);
	Full_Adder FA3600 (pp2[2], pp3[1], pp4[0], S[3662], Cout[3662]);
	Full_Adder FA3601 (pp5[0], Cout[3423], S[3424], S[3663], Cout[3663]);
	Full_Adder FA3602 (Cout[3424], Cout[3425], S[3426], S[3664], Cout[3664]);
	Full_Adder FA3603 (Cout[3426], Cout[3427], S[3428], S[3665], Cout[3665]);
	Full_Adder FA3604 (Cout[3428], Cout[3429], S[3430], S[3666], Cout[3666]);
	Full_Adder FA3605 (Cout[3430], Cout[3431], S[3432], S[3667], Cout[3667]);
	Full_Adder FA3606 (Cout[3432], Cout[3433], S[3434], S[3668], Cout[3668]);
	Full_Adder FA3607 (Cout[3434], Cout[3435], S[3436], S[3669], Cout[3669]);
	Full_Adder FA3608 (Cout[3436], Cout[3437], S[3438], S[3670], Cout[3670]);
	Full_Adder FA3609 (Cout[3438], Cout[3439], S[3440], S[3671], Cout[3671]);
	Full_Adder FA3610 (Cout[3440], Cout[3441], S[3442], S[3672], Cout[3672]);
	Full_Adder FA3611 (Cout[3442], Cout[3443], S[3444], S[3673], Cout[3673]);
	Full_Adder FA3612 (Cout[3444], Cout[3445], S[3446], S[3674], Cout[3674]);
	Full_Adder FA3613 (Cout[3446], Cout[3447], S[3448], S[3675], Cout[3675]);
	Full_Adder FA3614 (Cout[3448], Cout[3449], S[3450], S[3676], Cout[3676]);
	Full_Adder FA3615 (Cout[3450], Cout[3451], S[3452], S[3677], Cout[3677]);
	Full_Adder FA3616 (Cout[3452], Cout[3453], S[3454], S[3678], Cout[3678]);
	Full_Adder FA3617 (Cout[3454], Cout[3455], S[3456], S[3679], Cout[3679]);
	Full_Adder FA3618 (Cout[3456], Cout[3457], S[3458], S[3680], Cout[3680]);
	Full_Adder FA3619 (Cout[3458], Cout[3459], S[3460], S[3681], Cout[3681]);
	Full_Adder FA3620 (Cout[3460], Cout[3461], S[3462], S[3682], Cout[3682]);
	Full_Adder FA3621 (Cout[3462], Cout[3463], S[3464], S[3683], Cout[3683]);
	Full_Adder FA3622 (Cout[3464], Cout[3465], S[3466], S[3684], Cout[3684]);
	Full_Adder FA3623 (Cout[3466], Cout[3467], S[3468], S[3685], Cout[3685]);
	Full_Adder FA3624 (Cout[3468], Cout[3469], S[3470], S[3686], Cout[3686]);
	Full_Adder FA3625 (Cout[3470], Cout[3471], S[3472], S[3687], Cout[3687]);
	Full_Adder FA3626 (Cout[3472], Cout[3473], S[3474], S[3688], Cout[3688]);
	Full_Adder FA3627 (Cout[3474], Cout[3475], S[3476], S[3689], Cout[3689]);
	Full_Adder FA3628 (Cout[3476], Cout[3477], S[3478], S[3690], Cout[3690]);
	Full_Adder FA3629 (Cout[3478], Cout[3479], S[3480], S[3691], Cout[3691]);
	Full_Adder FA3630 (Cout[3480], Cout[3481], S[3482], S[3692], Cout[3692]);
	Full_Adder FA3631 (Cout[3482], Cout[3483], S[3484], S[3693], Cout[3693]);
	Full_Adder FA3632 (Cout[3484], Cout[3485], S[3486], S[3694], Cout[3694]);
	Full_Adder FA3633 (Cout[3486], Cout[3487], S[3488], S[3695], Cout[3695]);
	Full_Adder FA3634 (Cout[3488], Cout[3489], S[3490], S[3696], Cout[3696]);
	Full_Adder FA3635 (Cout[3490], Cout[3491], S[3492], S[3697], Cout[3697]);
	Full_Adder FA3636 (Cout[3492], Cout[3493], S[3494], S[3698], Cout[3698]);
	Full_Adder FA3637 (Cout[3494], Cout[3495], S[3496], S[3699], Cout[3699]);
	Full_Adder FA3638 (Cout[3496], Cout[3497], S[3498], S[3700], Cout[3700]);
	Full_Adder FA3639 (Cout[3498], Cout[3499], S[3500], S[3701], Cout[3701]);
	Full_Adder FA3640 (Cout[3500], Cout[3501], S[3502], S[3702], Cout[3702]);
	Full_Adder FA3641 (Cout[3502], Cout[3503], S[3504], S[3703], Cout[3703]);
	Full_Adder FA3642 (Cout[3504], Cout[3505], S[3506], S[3704], Cout[3704]);
	Full_Adder FA3643 (Cout[3506], Cout[3507], S[3508], S[3705], Cout[3705]);
	Full_Adder FA3644 (Cout[3508], Cout[3509], S[3510], S[3706], Cout[3706]);
	Full_Adder FA3645 (Cout[3510], Cout[3511], S[3512], S[3707], Cout[3707]);
	Full_Adder FA3646 (Cout[3512], Cout[3513], S[3514], S[3708], Cout[3708]);
	Full_Adder FA3647 (Cout[3514], Cout[3515], S[3516], S[3709], Cout[3709]);
	Full_Adder FA3648 (Cout[3516], Cout[3517], S[3518], S[3710], Cout[3710]);
	Full_Adder FA3649 (Cout[3518], Cout[3519], S[3520], S[3711], Cout[3711]);
	Full_Adder FA3650 (Cout[3520], Cout[3521], S[3522], S[3712], Cout[3712]);
	Full_Adder FA3651 (Cout[3522], Cout[3523], S[3524], S[3713], Cout[3713]);
	Full_Adder FA3652 (Cout[3524], Cout[3525], S[3526], S[3714], Cout[3714]);
	Full_Adder FA3653 (Cout[3526], Cout[3527], S[3528], S[3715], Cout[3715]);
	Full_Adder FA3654 (Cout[3528], Cout[3529], S[3530], S[3716], Cout[3716]);
	Full_Adder FA3655 (Cout[3530], Cout[3531], S[3532], S[3717], Cout[3717]);
	Full_Adder FA3656 (Cout[3532], Cout[3533], S[3534], S[3718], Cout[3718]);
	Full_Adder FA3657 (Cout[3534], Cout[3535], S[3536], S[3719], Cout[3719]);
	Full_Adder FA3658 (Cout[3536], Cout[3537], S[3538], S[3720], Cout[3720]);
	Full_Adder FA3659 (Cout[3538], Cout[3539], S[3540], S[3721], Cout[3721]);
	Full_Adder FA3660 (Cout[3540], Cout[3541], S[3542], S[3722], Cout[3722]);
	Full_Adder FA3661 (Cout[3542], Cout[3543], S[3544], S[3723], Cout[3723]);
	Full_Adder FA3662 (Cout[3544], Cout[3545], S[3546], S[3724], Cout[3724]);
	Full_Adder FA3663 (Cout[3546], Cout[3547], S[3548], S[3725], Cout[3725]);
	Full_Adder FA3664 (Cout[3548], Cout[3549], S[3550], S[3726], Cout[3726]);
	Full_Adder FA3665 (Cout[3550], Cout[3551], S[3552], S[3727], Cout[3727]);
	Full_Adder FA3666 (Cout[3552], Cout[3553], S[3554], S[3728], Cout[3728]);
	Full_Adder FA3667 (Cout[3554], Cout[3555], S[3556], S[3729], Cout[3729]);
	Full_Adder FA3668 (Cout[3556], Cout[3557], S[3558], S[3730], Cout[3730]);
	Full_Adder FA3669 (Cout[3558], Cout[3559], S[3560], S[3731], Cout[3731]);
	Full_Adder FA3670 (Cout[3560], Cout[3561], S[3562], S[3732], Cout[3732]);
	Full_Adder FA3671 (Cout[3562], Cout[3563], S[3564], S[3733], Cout[3733]);
	Full_Adder FA3672 (Cout[3564], Cout[3565], S[3566], S[3734], Cout[3734]);
	Full_Adder FA3673 (Cout[3566], Cout[3567], S[3568], S[3735], Cout[3735]);
	Full_Adder FA3674 (Cout[3568], Cout[3569], S[3570], S[3736], Cout[3736]);
	Full_Adder FA3675 (Cout[3570], Cout[3571], S[3572], S[3737], Cout[3737]);
	Full_Adder FA3676 (Cout[3572], Cout[3573], S[3574], S[3738], Cout[3738]);
	Full_Adder FA3677 (Cout[3574], Cout[3575], S[3576], S[3739], Cout[3739]);
	Full_Adder FA3678 (Cout[3576], Cout[3577], S[3578], S[3740], Cout[3740]);
	Full_Adder FA3679 (Cout[3578], Cout[3579], S[3580], S[3741], Cout[3741]);
	Full_Adder FA3680 (Cout[3580], Cout[3581], S[3582], S[3742], Cout[3742]);
	Full_Adder FA3681 (Cout[3582], Cout[3583], S[3584], S[3743], Cout[3743]);
	Full_Adder FA3682 (Cout[3584], Cout[3585], S[3586], S[3744], Cout[3744]);
	Full_Adder FA3683 (Cout[3586], Cout[3587], S[3588], S[3745], Cout[3745]);
	Full_Adder FA3684 (Cout[3588], Cout[3589], S[3590], S[3746], Cout[3746]);
	Full_Adder FA3685 (Cout[3590], Cout[3591], S[3592], S[3747], Cout[3747]);
	Full_Adder FA3686 (Cout[3592], Cout[3593], S[3594], S[3748], Cout[3748]);
	Full_Adder FA3687 (Cout[3594], Cout[3595], S[3596], S[3749], Cout[3749]);
	Full_Adder FA3688 (Cout[3596], Cout[3597], S[3598], S[3750], Cout[3750]);
	Full_Adder FA3689 (Cout[3598], Cout[3599], S[3600], S[3751], Cout[3751]);
	Full_Adder FA3690 (Cout[3600], Cout[3601], S[3602], S[3752], Cout[3752]);
	Full_Adder FA3691 (Cout[3602], Cout[3603], S[3604], S[3753], Cout[3753]);
	Full_Adder FA3692 (Cout[3604], Cout[3605], S[3606], S[3754], Cout[3754]);
	Full_Adder FA3693 (Cout[3606], Cout[3607], S[3608], S[3755], Cout[3755]);
	Full_Adder FA3694 (Cout[3608], Cout[3609], S[3610], S[3756], Cout[3756]);
	Full_Adder FA3695 (Cout[3610], Cout[3611], S[3612], S[3757], Cout[3757]);
	Full_Adder FA3696 (Cout[3612], Cout[3613], S[3614], S[3758], Cout[3758]);
	Full_Adder FA3697 (Cout[3614], Cout[3615], S[3616], S[3759], Cout[3759]);
	Full_Adder FA3698 (Cout[3616], Cout[3617], S[3618], S[3760], Cout[3760]);
	Full_Adder FA3699 (Cout[3618], Cout[3619], S[3620], S[3761], Cout[3761]);
	Full_Adder FA3700 (Cout[3620], Cout[3621], S[3622], S[3762], Cout[3762]);
	Full_Adder FA3701 (Cout[3622], Cout[3623], S[3624], S[3763], Cout[3763]);
	Full_Adder FA3702 (Cout[3624], Cout[3625], S[3626], S[3764], Cout[3764]);
	Full_Adder FA3703 (Cout[3626], Cout[3627], S[3628], S[3765], Cout[3765]);
	Full_Adder FA3704 (Cout[3628], Cout[3629], S[3630], S[3766], Cout[3766]);
	Full_Adder FA3705 (Cout[3630], Cout[3631], S[3632], S[3767], Cout[3767]);
	Full_Adder FA3706 (Cout[3632], Cout[3633], S[3634], S[3768], Cout[3768]);
	Full_Adder FA3707 (Cout[3634], Cout[3635], S[3636], S[3769], Cout[3769]);
	Full_Adder FA3708 (Cout[3636], Cout[3637], S[3638], S[3770], Cout[3770]);
	Full_Adder FA3709 (Cout[3638], Cout[3639], S[3640], S[3771], Cout[3771]);
	Full_Adder FA3710 (Cout[3640], Cout[3641], S[3642], S[3772], Cout[3772]);
	Full_Adder FA3711 (Cout[3642], Cout[3643], S[3644], S[3773], Cout[3773]);
	Full_Adder FA3712 (Cout[3644], Cout[3645], S[3646], S[3774], Cout[3774]);
	Full_Adder FA3713 (Cout[3646], Cout[3647], S[3648], S[3775], Cout[3775]);
	Full_Adder FA3714 (Cout[3648], Cout[3649], S[3650], S[3776], Cout[3776]);
	Full_Adder FA3715 (Cout[3650], Cout[3651], S[3652], S[3777], Cout[3777]);
	Full_Adder FA3716 (Cout[3652], Cout[3653], S[3654], S[3778], Cout[3778]);
	Full_Adder FA3717 (Cout[3654], Cout[3655], S[3656], S[3779], Cout[3779]);
	Full_Adder FA3718 (Cout[3656], Cout[3657], S[3658], S[3780], Cout[3780]);
	Full_Adder FA3719 (pp63[60], Cout[3658], Cout[3659], S[3781], Cout[3781]);
	Full_Adder FA3720 (pp61[63], pp62[62], pp63[61], S[3782], Cout[3782]);
	Half_Adder HA63 (pp0[2], pp1[1], S[3783], Cout[3783]);
	Full_Adder FA3721 (pp2[1], pp3[0], S[3661], S[3784], Cout[3784]);
	Full_Adder FA3722 (S[3423], Cout[3661], S[3662], S[3785], Cout[3785]);
	Full_Adder FA3723 (S[3425], Cout[3662], S[3663], S[3786], Cout[3786]);
	Full_Adder FA3724 (S[3427], Cout[3663], S[3664], S[3787], Cout[3787]);
	Full_Adder FA3725 (S[3429], Cout[3664], S[3665], S[3788], Cout[3788]);
	Full_Adder FA3726 (S[3431], Cout[3665], S[3666], S[3789], Cout[3789]);
	Full_Adder FA3727 (S[3433], Cout[3666], S[3667], S[3790], Cout[3790]);
	Full_Adder FA3728 (S[3435], Cout[3667], S[3668], S[3791], Cout[3791]);
	Full_Adder FA3729 (S[3437], Cout[3668], S[3669], S[3792], Cout[3792]);
	Full_Adder FA3730 (S[3439], Cout[3669], S[3670], S[3793], Cout[3793]);
	Full_Adder FA3731 (S[3441], Cout[3670], S[3671], S[3794], Cout[3794]);
	Full_Adder FA3732 (S[3443], Cout[3671], S[3672], S[3795], Cout[3795]);
	Full_Adder FA3733 (S[3445], Cout[3672], S[3673], S[3796], Cout[3796]);
	Full_Adder FA3734 (S[3447], Cout[3673], S[3674], S[3797], Cout[3797]);
	Full_Adder FA3735 (S[3449], Cout[3674], S[3675], S[3798], Cout[3798]);
	Full_Adder FA3736 (S[3451], Cout[3675], S[3676], S[3799], Cout[3799]);
	Full_Adder FA3737 (S[3453], Cout[3676], S[3677], S[3800], Cout[3800]);
	Full_Adder FA3738 (S[3455], Cout[3677], S[3678], S[3801], Cout[3801]);
	Full_Adder FA3739 (S[3457], Cout[3678], S[3679], S[3802], Cout[3802]);
	Full_Adder FA3740 (S[3459], Cout[3679], S[3680], S[3803], Cout[3803]);
	Full_Adder FA3741 (S[3461], Cout[3680], S[3681], S[3804], Cout[3804]);
	Full_Adder FA3742 (S[3463], Cout[3681], S[3682], S[3805], Cout[3805]);
	Full_Adder FA3743 (S[3465], Cout[3682], S[3683], S[3806], Cout[3806]);
	Full_Adder FA3744 (S[3467], Cout[3683], S[3684], S[3807], Cout[3807]);
	Full_Adder FA3745 (S[3469], Cout[3684], S[3685], S[3808], Cout[3808]);
	Full_Adder FA3746 (S[3471], Cout[3685], S[3686], S[3809], Cout[3809]);
	Full_Adder FA3747 (S[3473], Cout[3686], S[3687], S[3810], Cout[3810]);
	Full_Adder FA3748 (S[3475], Cout[3687], S[3688], S[3811], Cout[3811]);
	Full_Adder FA3749 (S[3477], Cout[3688], S[3689], S[3812], Cout[3812]);
	Full_Adder FA3750 (S[3479], Cout[3689], S[3690], S[3813], Cout[3813]);
	Full_Adder FA3751 (S[3481], Cout[3690], S[3691], S[3814], Cout[3814]);
	Full_Adder FA3752 (S[3483], Cout[3691], S[3692], S[3815], Cout[3815]);
	Full_Adder FA3753 (S[3485], Cout[3692], S[3693], S[3816], Cout[3816]);
	Full_Adder FA3754 (S[3487], Cout[3693], S[3694], S[3817], Cout[3817]);
	Full_Adder FA3755 (S[3489], Cout[3694], S[3695], S[3818], Cout[3818]);
	Full_Adder FA3756 (S[3491], Cout[3695], S[3696], S[3819], Cout[3819]);
	Full_Adder FA3757 (S[3493], Cout[3696], S[3697], S[3820], Cout[3820]);
	Full_Adder FA3758 (S[3495], Cout[3697], S[3698], S[3821], Cout[3821]);
	Full_Adder FA3759 (S[3497], Cout[3698], S[3699], S[3822], Cout[3822]);
	Full_Adder FA3760 (S[3499], Cout[3699], S[3700], S[3823], Cout[3823]);
	Full_Adder FA3761 (S[3501], Cout[3700], S[3701], S[3824], Cout[3824]);
	Full_Adder FA3762 (S[3503], Cout[3701], S[3702], S[3825], Cout[3825]);
	Full_Adder FA3763 (S[3505], Cout[3702], S[3703], S[3826], Cout[3826]);
	Full_Adder FA3764 (S[3507], Cout[3703], S[3704], S[3827], Cout[3827]);
	Full_Adder FA3765 (S[3509], Cout[3704], S[3705], S[3828], Cout[3828]);
	Full_Adder FA3766 (S[3511], Cout[3705], S[3706], S[3829], Cout[3829]);
	Full_Adder FA3767 (S[3513], Cout[3706], S[3707], S[3830], Cout[3830]);
	Full_Adder FA3768 (S[3515], Cout[3707], S[3708], S[3831], Cout[3831]);
	Full_Adder FA3769 (S[3517], Cout[3708], S[3709], S[3832], Cout[3832]);
	Full_Adder FA3770 (S[3519], Cout[3709], S[3710], S[3833], Cout[3833]);
	Full_Adder FA3771 (S[3521], Cout[3710], S[3711], S[3834], Cout[3834]);
	Full_Adder FA3772 (S[3523], Cout[3711], S[3712], S[3835], Cout[3835]);
	Full_Adder FA3773 (S[3525], Cout[3712], S[3713], S[3836], Cout[3836]);
	Full_Adder FA3774 (S[3527], Cout[3713], S[3714], S[3837], Cout[3837]);
	Full_Adder FA3775 (S[3529], Cout[3714], S[3715], S[3838], Cout[3838]);
	Full_Adder FA3776 (S[3531], Cout[3715], S[3716], S[3839], Cout[3839]);
	Full_Adder FA3777 (S[3533], Cout[3716], S[3717], S[3840], Cout[3840]);
	Full_Adder FA3778 (S[3535], Cout[3717], S[3718], S[3841], Cout[3841]);
	Full_Adder FA3779 (S[3537], Cout[3718], S[3719], S[3842], Cout[3842]);
	Full_Adder FA3780 (S[3539], Cout[3719], S[3720], S[3843], Cout[3843]);
	Full_Adder FA3781 (S[3541], Cout[3720], S[3721], S[3844], Cout[3844]);
	Full_Adder FA3782 (S[3543], Cout[3721], S[3722], S[3845], Cout[3845]);
	Full_Adder FA3783 (S[3545], Cout[3722], S[3723], S[3846], Cout[3846]);
	Full_Adder FA3784 (S[3547], Cout[3723], S[3724], S[3847], Cout[3847]);
	Full_Adder FA3785 (S[3549], Cout[3724], S[3725], S[3848], Cout[3848]);
	Full_Adder FA3786 (S[3551], Cout[3725], S[3726], S[3849], Cout[3849]);
	Full_Adder FA3787 (S[3553], Cout[3726], S[3727], S[3850], Cout[3850]);
	Full_Adder FA3788 (S[3555], Cout[3727], S[3728], S[3851], Cout[3851]);
	Full_Adder FA3789 (S[3557], Cout[3728], S[3729], S[3852], Cout[3852]);
	Full_Adder FA3790 (S[3559], Cout[3729], S[3730], S[3853], Cout[3853]);
	Full_Adder FA3791 (S[3561], Cout[3730], S[3731], S[3854], Cout[3854]);
	Full_Adder FA3792 (S[3563], Cout[3731], S[3732], S[3855], Cout[3855]);
	Full_Adder FA3793 (S[3565], Cout[3732], S[3733], S[3856], Cout[3856]);
	Full_Adder FA3794 (S[3567], Cout[3733], S[3734], S[3857], Cout[3857]);
	Full_Adder FA3795 (S[3569], Cout[3734], S[3735], S[3858], Cout[3858]);
	Full_Adder FA3796 (S[3571], Cout[3735], S[3736], S[3859], Cout[3859]);
	Full_Adder FA3797 (S[3573], Cout[3736], S[3737], S[3860], Cout[3860]);
	Full_Adder FA3798 (S[3575], Cout[3737], S[3738], S[3861], Cout[3861]);
	Full_Adder FA3799 (S[3577], Cout[3738], S[3739], S[3862], Cout[3862]);
	Full_Adder FA3800 (S[3579], Cout[3739], S[3740], S[3863], Cout[3863]);
	Full_Adder FA3801 (S[3581], Cout[3740], S[3741], S[3864], Cout[3864]);
	Full_Adder FA3802 (S[3583], Cout[3741], S[3742], S[3865], Cout[3865]);
	Full_Adder FA3803 (S[3585], Cout[3742], S[3743], S[3866], Cout[3866]);
	Full_Adder FA3804 (S[3587], Cout[3743], S[3744], S[3867], Cout[3867]);
	Full_Adder FA3805 (S[3589], Cout[3744], S[3745], S[3868], Cout[3868]);
	Full_Adder FA3806 (S[3591], Cout[3745], S[3746], S[3869], Cout[3869]);
	Full_Adder FA3807 (S[3593], Cout[3746], S[3747], S[3870], Cout[3870]);
	Full_Adder FA3808 (S[3595], Cout[3747], S[3748], S[3871], Cout[3871]);
	Full_Adder FA3809 (S[3597], Cout[3748], S[3749], S[3872], Cout[3872]);
	Full_Adder FA3810 (S[3599], Cout[3749], S[3750], S[3873], Cout[3873]);
	Full_Adder FA3811 (S[3601], Cout[3750], S[3751], S[3874], Cout[3874]);
	Full_Adder FA3812 (S[3603], Cout[3751], S[3752], S[3875], Cout[3875]);
	Full_Adder FA3813 (S[3605], Cout[3752], S[3753], S[3876], Cout[3876]);
	Full_Adder FA3814 (S[3607], Cout[3753], S[3754], S[3877], Cout[3877]);
	Full_Adder FA3815 (S[3609], Cout[3754], S[3755], S[3878], Cout[3878]);
	Full_Adder FA3816 (S[3611], Cout[3755], S[3756], S[3879], Cout[3879]);
	Full_Adder FA3817 (S[3613], Cout[3756], S[3757], S[3880], Cout[3880]);
	Full_Adder FA3818 (S[3615], Cout[3757], S[3758], S[3881], Cout[3881]);
	Full_Adder FA3819 (S[3617], Cout[3758], S[3759], S[3882], Cout[3882]);
	Full_Adder FA3820 (S[3619], Cout[3759], S[3760], S[3883], Cout[3883]);
	Full_Adder FA3821 (S[3621], Cout[3760], S[3761], S[3884], Cout[3884]);
	Full_Adder FA3822 (S[3623], Cout[3761], S[3762], S[3885], Cout[3885]);
	Full_Adder FA3823 (S[3625], Cout[3762], S[3763], S[3886], Cout[3886]);
	Full_Adder FA3824 (S[3627], Cout[3763], S[3764], S[3887], Cout[3887]);
	Full_Adder FA3825 (S[3629], Cout[3764], S[3765], S[3888], Cout[3888]);
	Full_Adder FA3826 (S[3631], Cout[3765], S[3766], S[3889], Cout[3889]);
	Full_Adder FA3827 (S[3633], Cout[3766], S[3767], S[3890], Cout[3890]);
	Full_Adder FA3828 (S[3635], Cout[3767], S[3768], S[3891], Cout[3891]);
	Full_Adder FA3829 (S[3637], Cout[3768], S[3769], S[3892], Cout[3892]);
	Full_Adder FA3830 (S[3639], Cout[3769], S[3770], S[3893], Cout[3893]);
	Full_Adder FA3831 (S[3641], Cout[3770], S[3771], S[3894], Cout[3894]);
	Full_Adder FA3832 (S[3643], Cout[3771], S[3772], S[3895], Cout[3895]);
	Full_Adder FA3833 (S[3645], Cout[3772], S[3773], S[3896], Cout[3896]);
	Full_Adder FA3834 (S[3647], Cout[3773], S[3774], S[3897], Cout[3897]);
	Full_Adder FA3835 (S[3649], Cout[3774], S[3775], S[3898], Cout[3898]);
	Full_Adder FA3836 (S[3651], Cout[3775], S[3776], S[3899], Cout[3899]);
	Full_Adder FA3837 (S[3653], Cout[3776], S[3777], S[3900], Cout[3900]);
	Full_Adder FA3838 (S[3655], Cout[3777], S[3778], S[3901], Cout[3901]);
	Full_Adder FA3839 (S[3657], Cout[3778], S[3779], S[3902], Cout[3902]);
	Full_Adder FA3840 (S[3659], Cout[3779], S[3780], S[3903], Cout[3903]);
	Full_Adder FA3841 (S[3660], Cout[3780], S[3781], S[3904], Cout[3904]);
	Full_Adder FA3842 (Cout[3660], Cout[3781], S[3782], S[3905], Cout[3905]);
	Full_Adder FA3843 (pp62[63], pp63[62], Cout[3782], S[3906], Cout[3906]);
	Half_Adder HA64 (pp0[1], pp1[0], S[0], Cout[0]);
	Full_Adder FA3844 (pp2[0], S[3783], Cout[0], S[3907], Cout[3907]);
	Full_Adder FA3845 (Cout[3783], S[3784], Cout[3907], S[3908], Cout[3908]);
	Full_Adder FA3846 (Cout[3784], S[3785], Cout[3908], S[3909], Cout[3909]);
	Full_Adder FA3847 (Cout[3785], S[3786], Cout[3909], S[3910], Cout[3910]);
	Full_Adder FA3848 (Cout[3786], S[3787], Cout[3910], S[3911], Cout[3911]);
	Full_Adder FA3849 (Cout[3787], S[3788], Cout[3911], S[3912], Cout[3912]);
	Full_Adder FA3850 (Cout[3788], S[3789], Cout[3912], S[3913], Cout[3913]);
	Full_Adder FA3851 (Cout[3789], S[3790], Cout[3913], S[3914], Cout[3914]);
	Full_Adder FA3852 (Cout[3790], S[3791], Cout[3914], S[3915], Cout[3915]);
	Full_Adder FA3853 (Cout[3791], S[3792], Cout[3915], S[3916], Cout[3916]);
	Full_Adder FA3854 (Cout[3792], S[3793], Cout[3916], S[3917], Cout[3917]);
	Full_Adder FA3855 (Cout[3793], S[3794], Cout[3917], S[3918], Cout[3918]);
	Full_Adder FA3856 (Cout[3794], S[3795], Cout[3918], S[3919], Cout[3919]);
	Full_Adder FA3857 (Cout[3795], S[3796], Cout[3919], S[3920], Cout[3920]);
	Full_Adder FA3858 (Cout[3796], S[3797], Cout[3920], S[3921], Cout[3921]);
	Full_Adder FA3859 (Cout[3797], S[3798], Cout[3921], S[3922], Cout[3922]);
	Full_Adder FA3860 (Cout[3798], S[3799], Cout[3922], S[3923], Cout[3923]);
	Full_Adder FA3861 (Cout[3799], S[3800], Cout[3923], S[3924], Cout[3924]);
	Full_Adder FA3862 (Cout[3800], S[3801], Cout[3924], S[3925], Cout[3925]);
	Full_Adder FA3863 (Cout[3801], S[3802], Cout[3925], S[3926], Cout[3926]);
	Full_Adder FA3864 (Cout[3802], S[3803], Cout[3926], S[3927], Cout[3927]);
	Full_Adder FA3865 (Cout[3803], S[3804], Cout[3927], S[3928], Cout[3928]);
	Full_Adder FA3866 (Cout[3804], S[3805], Cout[3928], S[3929], Cout[3929]);
	Full_Adder FA3867 (Cout[3805], S[3806], Cout[3929], S[3930], Cout[3930]);
	Full_Adder FA3868 (Cout[3806], S[3807], Cout[3930], S[3931], Cout[3931]);
	Full_Adder FA3869 (Cout[3807], S[3808], Cout[3931], S[3932], Cout[3932]);
	Full_Adder FA3870 (Cout[3808], S[3809], Cout[3932], S[3933], Cout[3933]);
	Full_Adder FA3871 (Cout[3809], S[3810], Cout[3933], S[3934], Cout[3934]);
	Full_Adder FA3872 (Cout[3810], S[3811], Cout[3934], S[3935], Cout[3935]);
	Full_Adder FA3873 (Cout[3811], S[3812], Cout[3935], S[3936], Cout[3936]);
	Full_Adder FA3874 (Cout[3812], S[3813], Cout[3936], S[3937], Cout[3937]);
	Full_Adder FA3875 (Cout[3813], S[3814], Cout[3937], S[3938], Cout[3938]);
	Full_Adder FA3876 (Cout[3814], S[3815], Cout[3938], S[3939], Cout[3939]);
	Full_Adder FA3877 (Cout[3815], S[3816], Cout[3939], S[3940], Cout[3940]);
	Full_Adder FA3878 (Cout[3816], S[3817], Cout[3940], S[3941], Cout[3941]);
	Full_Adder FA3879 (Cout[3817], S[3818], Cout[3941], S[3942], Cout[3942]);
	Full_Adder FA3880 (Cout[3818], S[3819], Cout[3942], S[3943], Cout[3943]);
	Full_Adder FA3881 (Cout[3819], S[3820], Cout[3943], S[3944], Cout[3944]);
	Full_Adder FA3882 (Cout[3820], S[3821], Cout[3944], S[3945], Cout[3945]);
	Full_Adder FA3883 (Cout[3821], S[3822], Cout[3945], S[3946], Cout[3946]);
	Full_Adder FA3884 (Cout[3822], S[3823], Cout[3946], S[3947], Cout[3947]);
	Full_Adder FA3885 (Cout[3823], S[3824], Cout[3947], S[3948], Cout[3948]);
	Full_Adder FA3886 (Cout[3824], S[3825], Cout[3948], S[3949], Cout[3949]);
	Full_Adder FA3887 (Cout[3825], S[3826], Cout[3949], S[3950], Cout[3950]);
	Full_Adder FA3888 (Cout[3826], S[3827], Cout[3950], S[3951], Cout[3951]);
	Full_Adder FA3889 (Cout[3827], S[3828], Cout[3951], S[3952], Cout[3952]);
	Full_Adder FA3890 (Cout[3828], S[3829], Cout[3952], S[3953], Cout[3953]);
	Full_Adder FA3891 (Cout[3829], S[3830], Cout[3953], S[3954], Cout[3954]);
	Full_Adder FA3892 (Cout[3830], S[3831], Cout[3954], S[3955], Cout[3955]);
	Full_Adder FA3893 (Cout[3831], S[3832], Cout[3955], S[3956], Cout[3956]);
	Full_Adder FA3894 (Cout[3832], S[3833], Cout[3956], S[3957], Cout[3957]);
	Full_Adder FA3895 (Cout[3833], S[3834], Cout[3957], S[3958], Cout[3958]);
	Full_Adder FA3896 (Cout[3834], S[3835], Cout[3958], S[3959], Cout[3959]);
	Full_Adder FA3897 (Cout[3835], S[3836], Cout[3959], S[3960], Cout[3960]);
	Full_Adder FA3898 (Cout[3836], S[3837], Cout[3960], S[3961], Cout[3961]);
	Full_Adder FA3899 (Cout[3837], S[3838], Cout[3961], S[3962], Cout[3962]);
	Full_Adder FA3900 (Cout[3838], S[3839], Cout[3962], S[3963], Cout[3963]);
	Full_Adder FA3901 (Cout[3839], S[3840], Cout[3963], S[3964], Cout[3964]);
	Full_Adder FA3902 (Cout[3840], S[3841], Cout[3964], S[3965], Cout[3965]);
	Full_Adder FA3903 (Cout[3841], S[3842], Cout[3965], S[3966], Cout[3966]);
	Full_Adder FA3904 (Cout[3842], S[3843], Cout[3966], S[3967], Cout[3967]);
	Full_Adder FA3905 (Cout[3843], S[3844], Cout[3967], S[3968], Cout[3968]);
	Full_Adder FA3906 (Cout[3844], S[3845], Cout[3968], S[3969], Cout[3969]);
	Full_Adder FA3907 (Cout[3845], S[3846], Cout[3969], S[3970], Cout[3970]);
	Full_Adder FA3908 (Cout[3846], S[3847], Cout[3970], S[3971], Cout[3971]);
	Full_Adder FA3909 (Cout[3847], S[3848], Cout[3971], S[3972], Cout[3972]);
	Full_Adder FA3910 (Cout[3848], S[3849], Cout[3972], S[3973], Cout[3973]);
	Full_Adder FA3911 (Cout[3849], S[3850], Cout[3973], S[3974], Cout[3974]);
	Full_Adder FA3912 (Cout[3850], S[3851], Cout[3974], S[3975], Cout[3975]);
	Full_Adder FA3913 (Cout[3851], S[3852], Cout[3975], S[3976], Cout[3976]);
	Full_Adder FA3914 (Cout[3852], S[3853], Cout[3976], S[3977], Cout[3977]);
	Full_Adder FA3915 (Cout[3853], S[3854], Cout[3977], S[3978], Cout[3978]);
	Full_Adder FA3916 (Cout[3854], S[3855], Cout[3978], S[3979], Cout[3979]);
	Full_Adder FA3917 (Cout[3855], S[3856], Cout[3979], S[3980], Cout[3980]);
	Full_Adder FA3918 (Cout[3856], S[3857], Cout[3980], S[3981], Cout[3981]);
	Full_Adder FA3919 (Cout[3857], S[3858], Cout[3981], S[3982], Cout[3982]);
	Full_Adder FA3920 (Cout[3858], S[3859], Cout[3982], S[3983], Cout[3983]);
	Full_Adder FA3921 (Cout[3859], S[3860], Cout[3983], S[3984], Cout[3984]);
	Full_Adder FA3922 (Cout[3860], S[3861], Cout[3984], S[3985], Cout[3985]);
	Full_Adder FA3923 (Cout[3861], S[3862], Cout[3985], S[3986], Cout[3986]);
	Full_Adder FA3924 (Cout[3862], S[3863], Cout[3986], S[3987], Cout[3987]);
	Full_Adder FA3925 (Cout[3863], S[3864], Cout[3987], S[3988], Cout[3988]);
	Full_Adder FA3926 (Cout[3864], S[3865], Cout[3988], S[3989], Cout[3989]);
	Full_Adder FA3927 (Cout[3865], S[3866], Cout[3989], S[3990], Cout[3990]);
	Full_Adder FA3928 (Cout[3866], S[3867], Cout[3990], S[3991], Cout[3991]);
	Full_Adder FA3929 (Cout[3867], S[3868], Cout[3991], S[3992], Cout[3992]);
	Full_Adder FA3930 (Cout[3868], S[3869], Cout[3992], S[3993], Cout[3993]);
	Full_Adder FA3931 (Cout[3869], S[3870], Cout[3993], S[3994], Cout[3994]);
	Full_Adder FA3932 (Cout[3870], S[3871], Cout[3994], S[3995], Cout[3995]);
	Full_Adder FA3933 (Cout[3871], S[3872], Cout[3995], S[3996], Cout[3996]);
	Full_Adder FA3934 (Cout[3872], S[3873], Cout[3996], S[3997], Cout[3997]);
	Full_Adder FA3935 (Cout[3873], S[3874], Cout[3997], S[3998], Cout[3998]);
	Full_Adder FA3936 (Cout[3874], S[3875], Cout[3998], S[3999], Cout[3999]);
	Full_Adder FA3937 (Cout[3875], S[3876], Cout[3999], S[4000], Cout[4000]);
	Full_Adder FA3938 (Cout[3876], S[3877], Cout[4000], S[4001], Cout[4001]);
	Full_Adder FA3939 (Cout[3877], S[3878], Cout[4001], S[4002], Cout[4002]);
	Full_Adder FA3940 (Cout[3878], S[3879], Cout[4002], S[4003], Cout[4003]);
	Full_Adder FA3941 (Cout[3879], S[3880], Cout[4003], S[4004], Cout[4004]);
	Full_Adder FA3942 (Cout[3880], S[3881], Cout[4004], S[4005], Cout[4005]);
	Full_Adder FA3943 (Cout[3881], S[3882], Cout[4005], S[4006], Cout[4006]);
	Full_Adder FA3944 (Cout[3882], S[3883], Cout[4006], S[4007], Cout[4007]);
	Full_Adder FA3945 (Cout[3883], S[3884], Cout[4007], S[4008], Cout[4008]);
	Full_Adder FA3946 (Cout[3884], S[3885], Cout[4008], S[4009], Cout[4009]);
	Full_Adder FA3947 (Cout[3885], S[3886], Cout[4009], S[4010], Cout[4010]);
	Full_Adder FA3948 (Cout[3886], S[3887], Cout[4010], S[4011], Cout[4011]);
	Full_Adder FA3949 (Cout[3887], S[3888], Cout[4011], S[4012], Cout[4012]);
	Full_Adder FA3950 (Cout[3888], S[3889], Cout[4012], S[4013], Cout[4013]);
	Full_Adder FA3951 (Cout[3889], S[3890], Cout[4013], S[4014], Cout[4014]);
	Full_Adder FA3952 (Cout[3890], S[3891], Cout[4014], S[4015], Cout[4015]);
	Full_Adder FA3953 (Cout[3891], S[3892], Cout[4015], S[4016], Cout[4016]);
	Full_Adder FA3954 (Cout[3892], S[3893], Cout[4016], S[4017], Cout[4017]);
	Full_Adder FA3955 (Cout[3893], S[3894], Cout[4017], S[4018], Cout[4018]);
	Full_Adder FA3956 (Cout[3894], S[3895], Cout[4018], S[4019], Cout[4019]);
	Full_Adder FA3957 (Cout[3895], S[3896], Cout[4019], S[4020], Cout[4020]);
	Full_Adder FA3958 (Cout[3896], S[3897], Cout[4020], S[4021], Cout[4021]);
	Full_Adder FA3959 (Cout[3897], S[3898], Cout[4021], S[4022], Cout[4022]);
	Full_Adder FA3960 (Cout[3898], S[3899], Cout[4022], S[4023], Cout[4023]);
	Full_Adder FA3961 (Cout[3899], S[3900], Cout[4023], S[4024], Cout[4024]);
	Full_Adder FA3962 (Cout[3900], S[3901], Cout[4024], S[4025], Cout[4025]);
	Full_Adder FA3963 (Cout[3901], S[3902], Cout[4025], S[4026], Cout[4026]);
	Full_Adder FA3964 (Cout[3902], S[3903], Cout[4026], S[4027], Cout[4027]);
	Full_Adder FA3965 (Cout[3903], S[3904], Cout[4027], S[4028], Cout[4028]);
	Full_Adder FA3966 (Cout[3904], S[3905], Cout[4028], S[4029], Cout[4029]);
	Full_Adder FA3967 (Cout[3905], S[3906], Cout[4029], S[4030], Cout[4030]);
	Full_Adder FA3968 (pp63[63], Cout[3906], Cout[4030], S[4031], Cout[4031]);

        wire[124:0] sum, in_1, in_2;
        wire c;
        assign in_1 = {pp2[0], Cout[3783], Cout[3784], Cout[3785], Cout[3786], Cout[3787], Cout[3788], Cout[3789], Cout[3790], Cout[3791], Cout[3792], Cout[3793], Cout[3794], Cout[3795], Cout[3796], Cout[3797], Cout[3798], Cout[3799], Cout[3800], Cout[3801], Cout[3802], Cout[3803], Cout[3804], Cout[3805], Cout[3806], Cout[3807], Cout[3808], Cout[3809], Cout[3810], Cout[3811], Cout[3812], Cout[3813], Cout[3814], Cout[3815], Cout[3816], Cout[3817], Cout[3818], Cout[3819], Cout[3820], Cout[3821], Cout[3822], Cout[3823], Cout[3824], Cout[3825], Cout[3826], Cout[3827], Cout[3828], Cout[3829], Cout[3830], Cout[3831], Cout[3832], Cout[3833], Cout[3834], Cout[3835], Cout[3836], Cout[3837], Cout[3838], Cout[3839], Cout[3840], Cout[3841], Cout[3842], Cout[3843], Cout[3844], Cout[3845], Cout[3846], Cout[3847], Cout[3848], Cout[3849], Cout[3850], Cout[3851], Cout[3852], Cout[3853], Cout[3854], Cout[3855], Cout[3856], Cout[3857], Cout[3858], Cout[3859], Cout[3860], Cout[3861], Cout[3862], Cout[3863], Cout[3864], Cout[3865], Cout[3866], Cout[3867], Cout[3868], Cout[3869], Cout[3870], Cout[3871], Cout[3872], Cout[3873], Cout[3874], Cout[3875], Cout[3876], Cout[3877], Cout[3878], Cout[3879], Cout[3880], Cout[3881], Cout[3882], Cout[3883], Cout[3884], Cout[3885], Cout[3886], Cout[3887], Cout[3888], Cout[3889], Cout[3890], Cout[3891], Cout[3892], Cout[3893], Cout[3894], Cout[3895], Cout[3896], Cout[3897], Cout[3898], Cout[3899], Cout[3900], Cout[3901], Cout[3902], Cout[3903], Cout[3904], Cout[3905], pp63[63]};
        assign in_1 = {S[3783], S[3784], S[3785], S[3786], S[3787], S[3788], S[3789], S[3790], S[3791], S[3792], S[3793], S[3794], S[3795], S[3796], S[3797], S[3798], S[3799], S[3800], S[3801], S[3802], S[3803], S[3804], S[3805], S[3806], S[3807], S[3808], S[3809], S[3810], S[3811], S[3812], S[3813], S[3814], S[3815], S[3816], S[3817], S[3818], S[3819], S[3820], S[3821], S[3822], S[3823], S[3824], S[3825], S[3826], S[3827], S[3828], S[3829], S[3830], S[3831], S[3832], S[3833], S[3834], S[3835], S[3836], S[3837], S[3838], S[3839], S[3840], S[3841], S[3842], S[3843], S[3844], S[3845], S[3846], S[3847], S[3848], S[3849], S[3850], S[3851], S[3852], S[3853], S[3854], S[3855], S[3856], S[3857], S[3858], S[3859], S[3860], S[3861], S[3862], S[3863], S[3864], S[3865], S[3866], S[3867], S[3868], S[3869], S[3870], S[3871], S[3872], S[3873], S[3874], S[3875], S[3876], S[3877], S[3878], S[3879], S[3880], S[3881], S[3882], S[3883], S[3884], S[3885], S[3886], S[3887], S[3888], S[3889], S[3890], S[3891], S[3892], S[3893], S[3894], S[3895], S[3896], S[3897], S[3898], S[3899], S[3900], S[3901], S[3902], S[3903], S[3904], S[3905], S[3906], Cout[3906]};
        CLA_125 CLA(sum, c, in_1, in_2);

	assign product[127] = c;
	assign product[126] = s[124];
	assign product[125] = s[123];
	assign product[124] = s[122];
	assign product[123] = s[121];
	assign product[122] = s[120];
	assign product[121] = s[119];
	assign product[120] = s[118];
	assign product[119] = s[117];
	assign product[118] = s[116];
	assign product[117] = s[115];
	assign product[116] = s[114];
	assign product[115] = s[113];
	assign product[114] = s[112];
	assign product[113] = s[111];
	assign product[112] = s[110];
	assign product[111] = s[109];
	assign product[110] = s[108];
	assign product[109] = s[107];
	assign product[108] = s[106];
	assign product[107] = s[105];
	assign product[106] = s[104];
	assign product[105] = s[103];
	assign product[104] = s[102];
	assign product[103] = s[101];
	assign product[102] = s[100];
	assign product[101] = s[99];
	assign product[100] = s[98];
	assign product[99]  = s[97];
	assign product[98]  = s[96];
	assign product[97]  = s[95];
	assign product[96]  = s[94];
	assign product[95]  = s[93];
	assign product[94]  = s[92];
	assign product[93]  = s[91];
	assign product[92]  = s[90];
	assign product[91]  = s[89];
	assign product[90]  = s[88];
	assign product[89]  = s[87];
	assign product[88]  = s[86];
	assign product[87]  = s[85];
	assign product[86]  = s[84];
	assign product[85]  = s[83];
	assign product[84]  = s[82];
	assign product[83]  = s[81];
	assign product[82]  = s[80];
	assign product[81]  = s[79];
	assign product[80]  = s[78];
	assign product[79]  = s[77];
	assign product[78]  = s[76];
	assign product[77]  = s[75];
	assign product[76]  = s[74];
	assign product[75]  = s[73];
	assign product[74]  = s[72];
	assign product[73]  = s[71];
	assign product[72]  = s[70];
	assign product[71]  = s[69];
	assign product[70]  = s[68];
	assign product[69]  = s[67];
	assign product[68]  = s[66];
	assign product[67]  = s[65];
	assign product[66]  = s[64];
	assign product[65]  = s[63];
	assign product[64]  = s[62];
	assign product[63]  = s[61];
	assign product[62]  = s[60];
	assign product[61]  = s[59];
	assign product[60]  = s[58];
	assign product[59]  = s[57];
	assign product[58]  = s[56];
	assign product[57]  = s[55];
	assign product[56]  = s[54];
	assign product[55]  = s[53];
	assign product[54]  = s[52];
	assign product[53]  = s[51];
	assign product[52]  = s[50];
	assign product[51]  = s[49];
	assign product[50]  = s[48];
	assign product[49]  = s[47];
	assign product[48]  = s[46];
	assign product[47]  = s[45];
	assign product[46]  = s[44];
	assign product[45]  = s[43];
	assign product[44]  = s[42];
	assign product[43]  = s[41];
	assign product[42]  = s[40];
	assign product[41]  = s[39];
	assign product[40]  = s[38];
	assign product[39]  = s[37];
	assign product[38]  = s[36];
	assign product[37]  = s[35];
	assign product[36]  = s[34];
	assign product[35]  = s[33];
	assign product[34]  = s[32];
	assign product[33]  = s[31];
	assign product[32]  = s[30;
	assign product[31]  = s[29];
	assign product[30]  = s[28];
	assign product[29]  = s[27];
	assign product[28]  = s[26];
	assign product[27]  = s[25];
	assign product[26]  = s[24];
	assign product[25]  = s[23];
	assign product[24]  = s[22];
	assign product[23]  = s[21];
	assign product[22]  = s[20];
	assign product[21]  = s[19];
	assign product[20]  = s[18];
	assign product[19]  = s[17];
	assign product[18]  = s[16];
	assign product[17]  = s[15];
	assign product[16]  = s[14];
	assign product[15]  = s[13];
	assign product[14]  = s[12];
	assign product[13]  = s[11];
	assign product[12]  = s[10];
	assign product[11]  = s[9];
	assign product[10]  = s[8];
	assign product[9]   = s[7];
	assign product[8]   = s[6];
	assign product[7]   = s[5];
	assign product[6]   = s[4];
	assign product[5]   = s[3];
	assign product[4]   = s[2];
	assign product[3]   = s[1];
	assign product[2]   = s[0];
	assign product[1]   = S[0];
	assign product[0]   = pp0[0];

endmodule

module CLA_128(output [127:0] sum, output cout, input [127:0] in1, input [127:0] in2);

    wire[127:0] G;
    wire[127:0] C;
    wire[127:0] P;

    assign G[0] = in1[127] & in2[127];
    assign P[0] = in1[127] ^ in2[127];
    assign G[1] = in1[126] & in2[126];
    assign P[1] = in1[126] ^ in2[126];
    assign G[2] = in1[125] & in2[125];
    assign P[2] = in1[125] ^ in2[125];
    assign G[3] = in1[124] & in2[124];
    assign P[3] = in1[124] ^ in2[124];
    assign G[4] = in1[123] & in2[123];
    assign P[4] = in1[123] ^ in2[123];
    assign G[5] = in1[122] & in2[122];
    assign P[5] = in1[122] ^ in2[122];
    assign G[6] = in1[121] & in2[121];
    assign P[6] = in1[121] ^ in2[121];
    assign G[7] = in1[120] & in2[120];
    assign P[7] = in1[120] ^ in2[120];
    assign G[8] = in1[119] & in2[119];
    assign P[8] = in1[119] ^ in2[119];
    assign G[9] = in1[118] & in2[118];
    assign P[9] = in1[118] ^ in2[118];
    assign G[10] = in1[117] & in2[117];
    assign P[10] = in1[117] ^ in2[117];
    assign G[11] = in1[116] & in2[116];
    assign P[11] = in1[116] ^ in2[116];
    assign G[12] = in1[115] & in2[115];
    assign P[12] = in1[115] ^ in2[115];
    assign G[13] = in1[114] & in2[114];
    assign P[13] = in1[114] ^ in2[114];
    assign G[14] = in1[113] & in2[113];
    assign P[14] = in1[113] ^ in2[113];
    assign G[15] = in1[112] & in2[112];
    assign P[15] = in1[112] ^ in2[112];
    assign G[16] = in1[111] & in2[111];
    assign P[16] = in1[111] ^ in2[111];
    assign G[17] = in1[110] & in2[110];
    assign P[17] = in1[110] ^ in2[110];
    assign G[18] = in1[109] & in2[109];
    assign P[18] = in1[109] ^ in2[109];
    assign G[19] = in1[108] & in2[108];
    assign P[19] = in1[108] ^ in2[108];
    assign G[20] = in1[107] & in2[107];
    assign P[20] = in1[107] ^ in2[107];
    assign G[21] = in1[106] & in2[106];
    assign P[21] = in1[106] ^ in2[106];
    assign G[22] = in1[105] & in2[105];
    assign P[22] = in1[105] ^ in2[105];
    assign G[23] = in1[104] & in2[104];
    assign P[23] = in1[104] ^ in2[104];
    assign G[24] = in1[103] & in2[103];
    assign P[24] = in1[103] ^ in2[103];
    assign G[25] = in1[102] & in2[102];
    assign P[25] = in1[102] ^ in2[102];
    assign G[26] = in1[101] & in2[101];
    assign P[26] = in1[101] ^ in2[101];
    assign G[27] = in1[100] & in2[100];
    assign P[27] = in1[100] ^ in2[100];
    assign G[28] = in1[99] & in2[99];
    assign P[28] = in1[99] ^ in2[99];
    assign G[29] = in1[98] & in2[98];
    assign P[29] = in1[98] ^ in2[98];
    assign G[30] = in1[97] & in2[97];
    assign P[30] = in1[97] ^ in2[97];
    assign G[31] = in1[96] & in2[96];
    assign P[31] = in1[96] ^ in2[96];
    assign G[32] = in1[95] & in2[95];
    assign P[32] = in1[95] ^ in2[95];
    assign G[33] = in1[94] & in2[94];
    assign P[33] = in1[94] ^ in2[94];
    assign G[34] = in1[93] & in2[93];
    assign P[34] = in1[93] ^ in2[93];
    assign G[35] = in1[92] & in2[92];
    assign P[35] = in1[92] ^ in2[92];
    assign G[36] = in1[91] & in2[91];
    assign P[36] = in1[91] ^ in2[91];
    assign G[37] = in1[90] & in2[90];
    assign P[37] = in1[90] ^ in2[90];
    assign G[38] = in1[89] & in2[89];
    assign P[38] = in1[89] ^ in2[89];
    assign G[39] = in1[88] & in2[88];
    assign P[39] = in1[88] ^ in2[88];
    assign G[40] = in1[87] & in2[87];
    assign P[40] = in1[87] ^ in2[87];
    assign G[41] = in1[86] & in2[86];
    assign P[41] = in1[86] ^ in2[86];
    assign G[42] = in1[85] & in2[85];
    assign P[42] = in1[85] ^ in2[85];
    assign G[43] = in1[84] & in2[84];
    assign P[43] = in1[84] ^ in2[84];
    assign G[44] = in1[83] & in2[83];
    assign P[44] = in1[83] ^ in2[83];
    assign G[45] = in1[82] & in2[82];
    assign P[45] = in1[82] ^ in2[82];
    assign G[46] = in1[81] & in2[81];
    assign P[46] = in1[81] ^ in2[81];
    assign G[47] = in1[80] & in2[80];
    assign P[47] = in1[80] ^ in2[80];
    assign G[48] = in1[79] & in2[79];
    assign P[48] = in1[79] ^ in2[79];
    assign G[49] = in1[78] & in2[78];
    assign P[49] = in1[78] ^ in2[78];
    assign G[50] = in1[77] & in2[77];
    assign P[50] = in1[77] ^ in2[77];
    assign G[51] = in1[76] & in2[76];
    assign P[51] = in1[76] ^ in2[76];
    assign G[52] = in1[75] & in2[75];
    assign P[52] = in1[75] ^ in2[75];
    assign G[53] = in1[74] & in2[74];
    assign P[53] = in1[74] ^ in2[74];
    assign G[54] = in1[73] & in2[73];
    assign P[54] = in1[73] ^ in2[73];
    assign G[55] = in1[72] & in2[72];
    assign P[55] = in1[72] ^ in2[72];
    assign G[56] = in1[71] & in2[71];
    assign P[56] = in1[71] ^ in2[71];
    assign G[57] = in1[70] & in2[70];
    assign P[57] = in1[70] ^ in2[70];
    assign G[58] = in1[69] & in2[69];
    assign P[58] = in1[69] ^ in2[69];
    assign G[59] = in1[68] & in2[68];
    assign P[59] = in1[68] ^ in2[68];
    assign G[60] = in1[67] & in2[67];
    assign P[60] = in1[67] ^ in2[67];
    assign G[61] = in1[66] & in2[66];
    assign P[61] = in1[66] ^ in2[66];
    assign G[62] = in1[65] & in2[65];
    assign P[62] = in1[65] ^ in2[65];
    assign G[63] = in1[64] & in2[64];
    assign P[63] = in1[64] ^ in2[64];
    assign G[64] = in1[63] & in2[63];
    assign P[64] = in1[63] ^ in2[63];
    assign G[65] = in1[62] & in2[62];
    assign P[65] = in1[62] ^ in2[62];
    assign G[66] = in1[61] & in2[61];
    assign P[66] = in1[61] ^ in2[61];
    assign G[67] = in1[60] & in2[60];
    assign P[67] = in1[60] ^ in2[60];
    assign G[68] = in1[59] & in2[59];
    assign P[68] = in1[59] ^ in2[59];
    assign G[69] = in1[58] & in2[58];
    assign P[69] = in1[58] ^ in2[58];
    assign G[70] = in1[57] & in2[57];
    assign P[70] = in1[57] ^ in2[57];
    assign G[71] = in1[56] & in2[56];
    assign P[71] = in1[56] ^ in2[56];
    assign G[72] = in1[55] & in2[55];
    assign P[72] = in1[55] ^ in2[55];
    assign G[73] = in1[54] & in2[54];
    assign P[73] = in1[54] ^ in2[54];
    assign G[74] = in1[53] & in2[53];
    assign P[74] = in1[53] ^ in2[53];
    assign G[75] = in1[52] & in2[52];
    assign P[75] = in1[52] ^ in2[52];
    assign G[76] = in1[51] & in2[51];
    assign P[76] = in1[51] ^ in2[51];
    assign G[77] = in1[50] & in2[50];
    assign P[77] = in1[50] ^ in2[50];
    assign G[78] = in1[49] & in2[49];
    assign P[78] = in1[49] ^ in2[49];
    assign G[79] = in1[48] & in2[48];
    assign P[79] = in1[48] ^ in2[48];
    assign G[80] = in1[47] & in2[47];
    assign P[80] = in1[47] ^ in2[47];
    assign G[81] = in1[46] & in2[46];
    assign P[81] = in1[46] ^ in2[46];
    assign G[82] = in1[45] & in2[45];
    assign P[82] = in1[45] ^ in2[45];
    assign G[83] = in1[44] & in2[44];
    assign P[83] = in1[44] ^ in2[44];
    assign G[84] = in1[43] & in2[43];
    assign P[84] = in1[43] ^ in2[43];
    assign G[85] = in1[42] & in2[42];
    assign P[85] = in1[42] ^ in2[42];
    assign G[86] = in1[41] & in2[41];
    assign P[86] = in1[41] ^ in2[41];
    assign G[87] = in1[40] & in2[40];
    assign P[87] = in1[40] ^ in2[40];
    assign G[88] = in1[39] & in2[39];
    assign P[88] = in1[39] ^ in2[39];
    assign G[89] = in1[38] & in2[38];
    assign P[89] = in1[38] ^ in2[38];
    assign G[90] = in1[37] & in2[37];
    assign P[90] = in1[37] ^ in2[37];
    assign G[91] = in1[36] & in2[36];
    assign P[91] = in1[36] ^ in2[36];
    assign G[92] = in1[35] & in2[35];
    assign P[92] = in1[35] ^ in2[35];
    assign G[93] = in1[34] & in2[34];
    assign P[93] = in1[34] ^ in2[34];
    assign G[94] = in1[33] & in2[33];
    assign P[94] = in1[33] ^ in2[33];
    assign G[95] = in1[32] & in2[32];
    assign P[95] = in1[32] ^ in2[32];
    assign G[96] = in1[31] & in2[31];
    assign P[96] = in1[31] ^ in2[31];
    assign G[97] = in1[30] & in2[30];
    assign P[97] = in1[30] ^ in2[30];
    assign G[98] = in1[29] & in2[29];
    assign P[98] = in1[29] ^ in2[29];
    assign G[99] = in1[28] & in2[28];
    assign P[99] = in1[28] ^ in2[28];
    assign G[100] = in1[27] & in2[27];
    assign P[100] = in1[27] ^ in2[27];
    assign G[101] = in1[26] & in2[26];
    assign P[101] = in1[26] ^ in2[26];
    assign G[102] = in1[25] & in2[25];
    assign P[102] = in1[25] ^ in2[25];
    assign G[103] = in1[24] & in2[24];
    assign P[103] = in1[24] ^ in2[24];
    assign G[104] = in1[23] & in2[23];
    assign P[104] = in1[23] ^ in2[23];
    assign G[105] = in1[22] & in2[22];
    assign P[105] = in1[22] ^ in2[22];
    assign G[106] = in1[21] & in2[21];
    assign P[106] = in1[21] ^ in2[21];
    assign G[107] = in1[20] & in2[20];
    assign P[107] = in1[20] ^ in2[20];
    assign G[108] = in1[19] & in2[19];
    assign P[108] = in1[19] ^ in2[19];
    assign G[109] = in1[18] & in2[18];
    assign P[109] = in1[18] ^ in2[18];
    assign G[110] = in1[17] & in2[17];
    assign P[110] = in1[17] ^ in2[17];
    assign G[111] = in1[16] & in2[16];
    assign P[111] = in1[16] ^ in2[16];
    assign G[112] = in1[15] & in2[15];
    assign P[112] = in1[15] ^ in2[15];
    assign G[113] = in1[14] & in2[14];
    assign P[113] = in1[14] ^ in2[14];
    assign G[114] = in1[13] & in2[13];
    assign P[114] = in1[13] ^ in2[13];
    assign G[115] = in1[12] & in2[12];
    assign P[115] = in1[12] ^ in2[12];
    assign G[116] = in1[11] & in2[11];
    assign P[116] = in1[11] ^ in2[11];
    assign G[117] = in1[10] & in2[10];
    assign P[117] = in1[10] ^ in2[10];
    assign G[118] = in1[9] & in2[9];
    assign P[118] = in1[9] ^ in2[9];
    assign G[119] = in1[8] & in2[8];
    assign P[119] = in1[8] ^ in2[8];
    assign G[120] = in1[7] & in2[7];
    assign P[120] = in1[7] ^ in2[7];
    assign G[121] = in1[6] & in2[6];
    assign P[121] = in1[6] ^ in2[6];
    assign G[122] = in1[5] & in2[5];
    assign P[122] = in1[5] ^ in2[5];
    assign G[123] = in1[4] & in2[4];
    assign P[123] = in1[4] ^ in2[4];
    assign G[124] = in1[3] & in2[3];
    assign P[124] = in1[3] ^ in2[3];
    assign G[125] = in1[2] & in2[2];
    assign P[125] = in1[2] ^ in2[2];
    assign G[126] = in1[1] & in2[1];
    assign P[126] = in1[1] ^ in2[1];
    assign G[127] = in1[0] & in2[0];
    assign P[127] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign cout = G[127] | (P[127] & C[127]);
    assign sum = P ^ C;
endmodule

module CLA_127(output [126:0] sum, output cout, input [126:0] in1, input [126:0] in2);

    wire[126:0] G;
    wire[126:0] C;
    wire[126:0] P;

    assign G[0] = in1[126] & in2[126];
    assign P[0] = in1[126] ^ in2[126];
    assign G[1] = in1[125] & in2[125];
    assign P[1] = in1[125] ^ in2[125];
    assign G[2] = in1[124] & in2[124];
    assign P[2] = in1[124] ^ in2[124];
    assign G[3] = in1[123] & in2[123];
    assign P[3] = in1[123] ^ in2[123];
    assign G[4] = in1[122] & in2[122];
    assign P[4] = in1[122] ^ in2[122];
    assign G[5] = in1[121] & in2[121];
    assign P[5] = in1[121] ^ in2[121];
    assign G[6] = in1[120] & in2[120];
    assign P[6] = in1[120] ^ in2[120];
    assign G[7] = in1[119] & in2[119];
    assign P[7] = in1[119] ^ in2[119];
    assign G[8] = in1[118] & in2[118];
    assign P[8] = in1[118] ^ in2[118];
    assign G[9] = in1[117] & in2[117];
    assign P[9] = in1[117] ^ in2[117];
    assign G[10] = in1[116] & in2[116];
    assign P[10] = in1[116] ^ in2[116];
    assign G[11] = in1[115] & in2[115];
    assign P[11] = in1[115] ^ in2[115];
    assign G[12] = in1[114] & in2[114];
    assign P[12] = in1[114] ^ in2[114];
    assign G[13] = in1[113] & in2[113];
    assign P[13] = in1[113] ^ in2[113];
    assign G[14] = in1[112] & in2[112];
    assign P[14] = in1[112] ^ in2[112];
    assign G[15] = in1[111] & in2[111];
    assign P[15] = in1[111] ^ in2[111];
    assign G[16] = in1[110] & in2[110];
    assign P[16] = in1[110] ^ in2[110];
    assign G[17] = in1[109] & in2[109];
    assign P[17] = in1[109] ^ in2[109];
    assign G[18] = in1[108] & in2[108];
    assign P[18] = in1[108] ^ in2[108];
    assign G[19] = in1[107] & in2[107];
    assign P[19] = in1[107] ^ in2[107];
    assign G[20] = in1[106] & in2[106];
    assign P[20] = in1[106] ^ in2[106];
    assign G[21] = in1[105] & in2[105];
    assign P[21] = in1[105] ^ in2[105];
    assign G[22] = in1[104] & in2[104];
    assign P[22] = in1[104] ^ in2[104];
    assign G[23] = in1[103] & in2[103];
    assign P[23] = in1[103] ^ in2[103];
    assign G[24] = in1[102] & in2[102];
    assign P[24] = in1[102] ^ in2[102];
    assign G[25] = in1[101] & in2[101];
    assign P[25] = in1[101] ^ in2[101];
    assign G[26] = in1[100] & in2[100];
    assign P[26] = in1[100] ^ in2[100];
    assign G[27] = in1[99] & in2[99];
    assign P[27] = in1[99] ^ in2[99];
    assign G[28] = in1[98] & in2[98];
    assign P[28] = in1[98] ^ in2[98];
    assign G[29] = in1[97] & in2[97];
    assign P[29] = in1[97] ^ in2[97];
    assign G[30] = in1[96] & in2[96];
    assign P[30] = in1[96] ^ in2[96];
    assign G[31] = in1[95] & in2[95];
    assign P[31] = in1[95] ^ in2[95];
    assign G[32] = in1[94] & in2[94];
    assign P[32] = in1[94] ^ in2[94];
    assign G[33] = in1[93] & in2[93];
    assign P[33] = in1[93] ^ in2[93];
    assign G[34] = in1[92] & in2[92];
    assign P[34] = in1[92] ^ in2[92];
    assign G[35] = in1[91] & in2[91];
    assign P[35] = in1[91] ^ in2[91];
    assign G[36] = in1[90] & in2[90];
    assign P[36] = in1[90] ^ in2[90];
    assign G[37] = in1[89] & in2[89];
    assign P[37] = in1[89] ^ in2[89];
    assign G[38] = in1[88] & in2[88];
    assign P[38] = in1[88] ^ in2[88];
    assign G[39] = in1[87] & in2[87];
    assign P[39] = in1[87] ^ in2[87];
    assign G[40] = in1[86] & in2[86];
    assign P[40] = in1[86] ^ in2[86];
    assign G[41] = in1[85] & in2[85];
    assign P[41] = in1[85] ^ in2[85];
    assign G[42] = in1[84] & in2[84];
    assign P[42] = in1[84] ^ in2[84];
    assign G[43] = in1[83] & in2[83];
    assign P[43] = in1[83] ^ in2[83];
    assign G[44] = in1[82] & in2[82];
    assign P[44] = in1[82] ^ in2[82];
    assign G[45] = in1[81] & in2[81];
    assign P[45] = in1[81] ^ in2[81];
    assign G[46] = in1[80] & in2[80];
    assign P[46] = in1[80] ^ in2[80];
    assign G[47] = in1[79] & in2[79];
    assign P[47] = in1[79] ^ in2[79];
    assign G[48] = in1[78] & in2[78];
    assign P[48] = in1[78] ^ in2[78];
    assign G[49] = in1[77] & in2[77];
    assign P[49] = in1[77] ^ in2[77];
    assign G[50] = in1[76] & in2[76];
    assign P[50] = in1[76] ^ in2[76];
    assign G[51] = in1[75] & in2[75];
    assign P[51] = in1[75] ^ in2[75];
    assign G[52] = in1[74] & in2[74];
    assign P[52] = in1[74] ^ in2[74];
    assign G[53] = in1[73] & in2[73];
    assign P[53] = in1[73] ^ in2[73];
    assign G[54] = in1[72] & in2[72];
    assign P[54] = in1[72] ^ in2[72];
    assign G[55] = in1[71] & in2[71];
    assign P[55] = in1[71] ^ in2[71];
    assign G[56] = in1[70] & in2[70];
    assign P[56] = in1[70] ^ in2[70];
    assign G[57] = in1[69] & in2[69];
    assign P[57] = in1[69] ^ in2[69];
    assign G[58] = in1[68] & in2[68];
    assign P[58] = in1[68] ^ in2[68];
    assign G[59] = in1[67] & in2[67];
    assign P[59] = in1[67] ^ in2[67];
    assign G[60] = in1[66] & in2[66];
    assign P[60] = in1[66] ^ in2[66];
    assign G[61] = in1[65] & in2[65];
    assign P[61] = in1[65] ^ in2[65];
    assign G[62] = in1[64] & in2[64];
    assign P[62] = in1[64] ^ in2[64];
    assign G[63] = in1[63] & in2[63];
    assign P[63] = in1[63] ^ in2[63];
    assign G[64] = in1[62] & in2[62];
    assign P[64] = in1[62] ^ in2[62];
    assign G[65] = in1[61] & in2[61];
    assign P[65] = in1[61] ^ in2[61];
    assign G[66] = in1[60] & in2[60];
    assign P[66] = in1[60] ^ in2[60];
    assign G[67] = in1[59] & in2[59];
    assign P[67] = in1[59] ^ in2[59];
    assign G[68] = in1[58] & in2[58];
    assign P[68] = in1[58] ^ in2[58];
    assign G[69] = in1[57] & in2[57];
    assign P[69] = in1[57] ^ in2[57];
    assign G[70] = in1[56] & in2[56];
    assign P[70] = in1[56] ^ in2[56];
    assign G[71] = in1[55] & in2[55];
    assign P[71] = in1[55] ^ in2[55];
    assign G[72] = in1[54] & in2[54];
    assign P[72] = in1[54] ^ in2[54];
    assign G[73] = in1[53] & in2[53];
    assign P[73] = in1[53] ^ in2[53];
    assign G[74] = in1[52] & in2[52];
    assign P[74] = in1[52] ^ in2[52];
    assign G[75] = in1[51] & in2[51];
    assign P[75] = in1[51] ^ in2[51];
    assign G[76] = in1[50] & in2[50];
    assign P[76] = in1[50] ^ in2[50];
    assign G[77] = in1[49] & in2[49];
    assign P[77] = in1[49] ^ in2[49];
    assign G[78] = in1[48] & in2[48];
    assign P[78] = in1[48] ^ in2[48];
    assign G[79] = in1[47] & in2[47];
    assign P[79] = in1[47] ^ in2[47];
    assign G[80] = in1[46] & in2[46];
    assign P[80] = in1[46] ^ in2[46];
    assign G[81] = in1[45] & in2[45];
    assign P[81] = in1[45] ^ in2[45];
    assign G[82] = in1[44] & in2[44];
    assign P[82] = in1[44] ^ in2[44];
    assign G[83] = in1[43] & in2[43];
    assign P[83] = in1[43] ^ in2[43];
    assign G[84] = in1[42] & in2[42];
    assign P[84] = in1[42] ^ in2[42];
    assign G[85] = in1[41] & in2[41];
    assign P[85] = in1[41] ^ in2[41];
    assign G[86] = in1[40] & in2[40];
    assign P[86] = in1[40] ^ in2[40];
    assign G[87] = in1[39] & in2[39];
    assign P[87] = in1[39] ^ in2[39];
    assign G[88] = in1[38] & in2[38];
    assign P[88] = in1[38] ^ in2[38];
    assign G[89] = in1[37] & in2[37];
    assign P[89] = in1[37] ^ in2[37];
    assign G[90] = in1[36] & in2[36];
    assign P[90] = in1[36] ^ in2[36];
    assign G[91] = in1[35] & in2[35];
    assign P[91] = in1[35] ^ in2[35];
    assign G[92] = in1[34] & in2[34];
    assign P[92] = in1[34] ^ in2[34];
    assign G[93] = in1[33] & in2[33];
    assign P[93] = in1[33] ^ in2[33];
    assign G[94] = in1[32] & in2[32];
    assign P[94] = in1[32] ^ in2[32];
    assign G[95] = in1[31] & in2[31];
    assign P[95] = in1[31] ^ in2[31];
    assign G[96] = in1[30] & in2[30];
    assign P[96] = in1[30] ^ in2[30];
    assign G[97] = in1[29] & in2[29];
    assign P[97] = in1[29] ^ in2[29];
    assign G[98] = in1[28] & in2[28];
    assign P[98] = in1[28] ^ in2[28];
    assign G[99] = in1[27] & in2[27];
    assign P[99] = in1[27] ^ in2[27];
    assign G[100] = in1[26] & in2[26];
    assign P[100] = in1[26] ^ in2[26];
    assign G[101] = in1[25] & in2[25];
    assign P[101] = in1[25] ^ in2[25];
    assign G[102] = in1[24] & in2[24];
    assign P[102] = in1[24] ^ in2[24];
    assign G[103] = in1[23] & in2[23];
    assign P[103] = in1[23] ^ in2[23];
    assign G[104] = in1[22] & in2[22];
    assign P[104] = in1[22] ^ in2[22];
    assign G[105] = in1[21] & in2[21];
    assign P[105] = in1[21] ^ in2[21];
    assign G[106] = in1[20] & in2[20];
    assign P[106] = in1[20] ^ in2[20];
    assign G[107] = in1[19] & in2[19];
    assign P[107] = in1[19] ^ in2[19];
    assign G[108] = in1[18] & in2[18];
    assign P[108] = in1[18] ^ in2[18];
    assign G[109] = in1[17] & in2[17];
    assign P[109] = in1[17] ^ in2[17];
    assign G[110] = in1[16] & in2[16];
    assign P[110] = in1[16] ^ in2[16];
    assign G[111] = in1[15] & in2[15];
    assign P[111] = in1[15] ^ in2[15];
    assign G[112] = in1[14] & in2[14];
    assign P[112] = in1[14] ^ in2[14];
    assign G[113] = in1[13] & in2[13];
    assign P[113] = in1[13] ^ in2[13];
    assign G[114] = in1[12] & in2[12];
    assign P[114] = in1[12] ^ in2[12];
    assign G[115] = in1[11] & in2[11];
    assign P[115] = in1[11] ^ in2[11];
    assign G[116] = in1[10] & in2[10];
    assign P[116] = in1[10] ^ in2[10];
    assign G[117] = in1[9] & in2[9];
    assign P[117] = in1[9] ^ in2[9];
    assign G[118] = in1[8] & in2[8];
    assign P[118] = in1[8] ^ in2[8];
    assign G[119] = in1[7] & in2[7];
    assign P[119] = in1[7] ^ in2[7];
    assign G[120] = in1[6] & in2[6];
    assign P[120] = in1[6] ^ in2[6];
    assign G[121] = in1[5] & in2[5];
    assign P[121] = in1[5] ^ in2[5];
    assign G[122] = in1[4] & in2[4];
    assign P[122] = in1[4] ^ in2[4];
    assign G[123] = in1[3] & in2[3];
    assign P[123] = in1[3] ^ in2[3];
    assign G[124] = in1[2] & in2[2];
    assign P[124] = in1[2] ^ in2[2];
    assign G[125] = in1[1] & in2[1];
    assign P[125] = in1[1] ^ in2[1];
    assign G[126] = in1[0] & in2[0];
    assign P[126] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign cout = G[126] | (P[126] & C[126]);
    assign sum = P ^ C;
endmodule

module CLA_126(output [125:0] sum, output cout, input [125:0] in1, input [125:0] in2);

    wire[125:0] G;
    wire[125:0] C;
    wire[125:0] P;

    assign G[0] = in1[125] & in2[125];
    assign P[0] = in1[125] ^ in2[125];
    assign G[1] = in1[124] & in2[124];
    assign P[1] = in1[124] ^ in2[124];
    assign G[2] = in1[123] & in2[123];
    assign P[2] = in1[123] ^ in2[123];
    assign G[3] = in1[122] & in2[122];
    assign P[3] = in1[122] ^ in2[122];
    assign G[4] = in1[121] & in2[121];
    assign P[4] = in1[121] ^ in2[121];
    assign G[5] = in1[120] & in2[120];
    assign P[5] = in1[120] ^ in2[120];
    assign G[6] = in1[119] & in2[119];
    assign P[6] = in1[119] ^ in2[119];
    assign G[7] = in1[118] & in2[118];
    assign P[7] = in1[118] ^ in2[118];
    assign G[8] = in1[117] & in2[117];
    assign P[8] = in1[117] ^ in2[117];
    assign G[9] = in1[116] & in2[116];
    assign P[9] = in1[116] ^ in2[116];
    assign G[10] = in1[115] & in2[115];
    assign P[10] = in1[115] ^ in2[115];
    assign G[11] = in1[114] & in2[114];
    assign P[11] = in1[114] ^ in2[114];
    assign G[12] = in1[113] & in2[113];
    assign P[12] = in1[113] ^ in2[113];
    assign G[13] = in1[112] & in2[112];
    assign P[13] = in1[112] ^ in2[112];
    assign G[14] = in1[111] & in2[111];
    assign P[14] = in1[111] ^ in2[111];
    assign G[15] = in1[110] & in2[110];
    assign P[15] = in1[110] ^ in2[110];
    assign G[16] = in1[109] & in2[109];
    assign P[16] = in1[109] ^ in2[109];
    assign G[17] = in1[108] & in2[108];
    assign P[17] = in1[108] ^ in2[108];
    assign G[18] = in1[107] & in2[107];
    assign P[18] = in1[107] ^ in2[107];
    assign G[19] = in1[106] & in2[106];
    assign P[19] = in1[106] ^ in2[106];
    assign G[20] = in1[105] & in2[105];
    assign P[20] = in1[105] ^ in2[105];
    assign G[21] = in1[104] & in2[104];
    assign P[21] = in1[104] ^ in2[104];
    assign G[22] = in1[103] & in2[103];
    assign P[22] = in1[103] ^ in2[103];
    assign G[23] = in1[102] & in2[102];
    assign P[23] = in1[102] ^ in2[102];
    assign G[24] = in1[101] & in2[101];
    assign P[24] = in1[101] ^ in2[101];
    assign G[25] = in1[100] & in2[100];
    assign P[25] = in1[100] ^ in2[100];
    assign G[26] = in1[99] & in2[99];
    assign P[26] = in1[99] ^ in2[99];
    assign G[27] = in1[98] & in2[98];
    assign P[27] = in1[98] ^ in2[98];
    assign G[28] = in1[97] & in2[97];
    assign P[28] = in1[97] ^ in2[97];
    assign G[29] = in1[96] & in2[96];
    assign P[29] = in1[96] ^ in2[96];
    assign G[30] = in1[95] & in2[95];
    assign P[30] = in1[95] ^ in2[95];
    assign G[31] = in1[94] & in2[94];
    assign P[31] = in1[94] ^ in2[94];
    assign G[32] = in1[93] & in2[93];
    assign P[32] = in1[93] ^ in2[93];
    assign G[33] = in1[92] & in2[92];
    assign P[33] = in1[92] ^ in2[92];
    assign G[34] = in1[91] & in2[91];
    assign P[34] = in1[91] ^ in2[91];
    assign G[35] = in1[90] & in2[90];
    assign P[35] = in1[90] ^ in2[90];
    assign G[36] = in1[89] & in2[89];
    assign P[36] = in1[89] ^ in2[89];
    assign G[37] = in1[88] & in2[88];
    assign P[37] = in1[88] ^ in2[88];
    assign G[38] = in1[87] & in2[87];
    assign P[38] = in1[87] ^ in2[87];
    assign G[39] = in1[86] & in2[86];
    assign P[39] = in1[86] ^ in2[86];
    assign G[40] = in1[85] & in2[85];
    assign P[40] = in1[85] ^ in2[85];
    assign G[41] = in1[84] & in2[84];
    assign P[41] = in1[84] ^ in2[84];
    assign G[42] = in1[83] & in2[83];
    assign P[42] = in1[83] ^ in2[83];
    assign G[43] = in1[82] & in2[82];
    assign P[43] = in1[82] ^ in2[82];
    assign G[44] = in1[81] & in2[81];
    assign P[44] = in1[81] ^ in2[81];
    assign G[45] = in1[80] & in2[80];
    assign P[45] = in1[80] ^ in2[80];
    assign G[46] = in1[79] & in2[79];
    assign P[46] = in1[79] ^ in2[79];
    assign G[47] = in1[78] & in2[78];
    assign P[47] = in1[78] ^ in2[78];
    assign G[48] = in1[77] & in2[77];
    assign P[48] = in1[77] ^ in2[77];
    assign G[49] = in1[76] & in2[76];
    assign P[49] = in1[76] ^ in2[76];
    assign G[50] = in1[75] & in2[75];
    assign P[50] = in1[75] ^ in2[75];
    assign G[51] = in1[74] & in2[74];
    assign P[51] = in1[74] ^ in2[74];
    assign G[52] = in1[73] & in2[73];
    assign P[52] = in1[73] ^ in2[73];
    assign G[53] = in1[72] & in2[72];
    assign P[53] = in1[72] ^ in2[72];
    assign G[54] = in1[71] & in2[71];
    assign P[54] = in1[71] ^ in2[71];
    assign G[55] = in1[70] & in2[70];
    assign P[55] = in1[70] ^ in2[70];
    assign G[56] = in1[69] & in2[69];
    assign P[56] = in1[69] ^ in2[69];
    assign G[57] = in1[68] & in2[68];
    assign P[57] = in1[68] ^ in2[68];
    assign G[58] = in1[67] & in2[67];
    assign P[58] = in1[67] ^ in2[67];
    assign G[59] = in1[66] & in2[66];
    assign P[59] = in1[66] ^ in2[66];
    assign G[60] = in1[65] & in2[65];
    assign P[60] = in1[65] ^ in2[65];
    assign G[61] = in1[64] & in2[64];
    assign P[61] = in1[64] ^ in2[64];
    assign G[62] = in1[63] & in2[63];
    assign P[62] = in1[63] ^ in2[63];
    assign G[63] = in1[62] & in2[62];
    assign P[63] = in1[62] ^ in2[62];
    assign G[64] = in1[61] & in2[61];
    assign P[64] = in1[61] ^ in2[61];
    assign G[65] = in1[60] & in2[60];
    assign P[65] = in1[60] ^ in2[60];
    assign G[66] = in1[59] & in2[59];
    assign P[66] = in1[59] ^ in2[59];
    assign G[67] = in1[58] & in2[58];
    assign P[67] = in1[58] ^ in2[58];
    assign G[68] = in1[57] & in2[57];
    assign P[68] = in1[57] ^ in2[57];
    assign G[69] = in1[56] & in2[56];
    assign P[69] = in1[56] ^ in2[56];
    assign G[70] = in1[55] & in2[55];
    assign P[70] = in1[55] ^ in2[55];
    assign G[71] = in1[54] & in2[54];
    assign P[71] = in1[54] ^ in2[54];
    assign G[72] = in1[53] & in2[53];
    assign P[72] = in1[53] ^ in2[53];
    assign G[73] = in1[52] & in2[52];
    assign P[73] = in1[52] ^ in2[52];
    assign G[74] = in1[51] & in2[51];
    assign P[74] = in1[51] ^ in2[51];
    assign G[75] = in1[50] & in2[50];
    assign P[75] = in1[50] ^ in2[50];
    assign G[76] = in1[49] & in2[49];
    assign P[76] = in1[49] ^ in2[49];
    assign G[77] = in1[48] & in2[48];
    assign P[77] = in1[48] ^ in2[48];
    assign G[78] = in1[47] & in2[47];
    assign P[78] = in1[47] ^ in2[47];
    assign G[79] = in1[46] & in2[46];
    assign P[79] = in1[46] ^ in2[46];
    assign G[80] = in1[45] & in2[45];
    assign P[80] = in1[45] ^ in2[45];
    assign G[81] = in1[44] & in2[44];
    assign P[81] = in1[44] ^ in2[44];
    assign G[82] = in1[43] & in2[43];
    assign P[82] = in1[43] ^ in2[43];
    assign G[83] = in1[42] & in2[42];
    assign P[83] = in1[42] ^ in2[42];
    assign G[84] = in1[41] & in2[41];
    assign P[84] = in1[41] ^ in2[41];
    assign G[85] = in1[40] & in2[40];
    assign P[85] = in1[40] ^ in2[40];
    assign G[86] = in1[39] & in2[39];
    assign P[86] = in1[39] ^ in2[39];
    assign G[87] = in1[38] & in2[38];
    assign P[87] = in1[38] ^ in2[38];
    assign G[88] = in1[37] & in2[37];
    assign P[88] = in1[37] ^ in2[37];
    assign G[89] = in1[36] & in2[36];
    assign P[89] = in1[36] ^ in2[36];
    assign G[90] = in1[35] & in2[35];
    assign P[90] = in1[35] ^ in2[35];
    assign G[91] = in1[34] & in2[34];
    assign P[91] = in1[34] ^ in2[34];
    assign G[92] = in1[33] & in2[33];
    assign P[92] = in1[33] ^ in2[33];
    assign G[93] = in1[32] & in2[32];
    assign P[93] = in1[32] ^ in2[32];
    assign G[94] = in1[31] & in2[31];
    assign P[94] = in1[31] ^ in2[31];
    assign G[95] = in1[30] & in2[30];
    assign P[95] = in1[30] ^ in2[30];
    assign G[96] = in1[29] & in2[29];
    assign P[96] = in1[29] ^ in2[29];
    assign G[97] = in1[28] & in2[28];
    assign P[97] = in1[28] ^ in2[28];
    assign G[98] = in1[27] & in2[27];
    assign P[98] = in1[27] ^ in2[27];
    assign G[99] = in1[26] & in2[26];
    assign P[99] = in1[26] ^ in2[26];
    assign G[100] = in1[25] & in2[25];
    assign P[100] = in1[25] ^ in2[25];
    assign G[101] = in1[24] & in2[24];
    assign P[101] = in1[24] ^ in2[24];
    assign G[102] = in1[23] & in2[23];
    assign P[102] = in1[23] ^ in2[23];
    assign G[103] = in1[22] & in2[22];
    assign P[103] = in1[22] ^ in2[22];
    assign G[104] = in1[21] & in2[21];
    assign P[104] = in1[21] ^ in2[21];
    assign G[105] = in1[20] & in2[20];
    assign P[105] = in1[20] ^ in2[20];
    assign G[106] = in1[19] & in2[19];
    assign P[106] = in1[19] ^ in2[19];
    assign G[107] = in1[18] & in2[18];
    assign P[107] = in1[18] ^ in2[18];
    assign G[108] = in1[17] & in2[17];
    assign P[108] = in1[17] ^ in2[17];
    assign G[109] = in1[16] & in2[16];
    assign P[109] = in1[16] ^ in2[16];
    assign G[110] = in1[15] & in2[15];
    assign P[110] = in1[15] ^ in2[15];
    assign G[111] = in1[14] & in2[14];
    assign P[111] = in1[14] ^ in2[14];
    assign G[112] = in1[13] & in2[13];
    assign P[112] = in1[13] ^ in2[13];
    assign G[113] = in1[12] & in2[12];
    assign P[113] = in1[12] ^ in2[12];
    assign G[114] = in1[11] & in2[11];
    assign P[114] = in1[11] ^ in2[11];
    assign G[115] = in1[10] & in2[10];
    assign P[115] = in1[10] ^ in2[10];
    assign G[116] = in1[9] & in2[9];
    assign P[116] = in1[9] ^ in2[9];
    assign G[117] = in1[8] & in2[8];
    assign P[117] = in1[8] ^ in2[8];
    assign G[118] = in1[7] & in2[7];
    assign P[118] = in1[7] ^ in2[7];
    assign G[119] = in1[6] & in2[6];
    assign P[119] = in1[6] ^ in2[6];
    assign G[120] = in1[5] & in2[5];
    assign P[120] = in1[5] ^ in2[5];
    assign G[121] = in1[4] & in2[4];
    assign P[121] = in1[4] ^ in2[4];
    assign G[122] = in1[3] & in2[3];
    assign P[122] = in1[3] ^ in2[3];
    assign G[123] = in1[2] & in2[2];
    assign P[123] = in1[2] ^ in2[2];
    assign G[124] = in1[1] & in2[1];
    assign P[124] = in1[1] ^ in2[1];
    assign G[125] = in1[0] & in2[0];
    assign P[125] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign cout = G[125] | (P[125] & C[125]);
    assign sum = P ^ C;
endmodule

module CLA_125(output [124:0] sum, output cout, input [124:0] in1, input [124:0] in2);

    wire[124:0] G;
    wire[124:0] C;
    wire[124:0] P;

    assign G[0] = in1[124] & in2[124];
    assign P[0] = in1[124] ^ in2[124];
    assign G[1] = in1[123] & in2[123];
    assign P[1] = in1[123] ^ in2[123];
    assign G[2] = in1[122] & in2[122];
    assign P[2] = in1[122] ^ in2[122];
    assign G[3] = in1[121] & in2[121];
    assign P[3] = in1[121] ^ in2[121];
    assign G[4] = in1[120] & in2[120];
    assign P[4] = in1[120] ^ in2[120];
    assign G[5] = in1[119] & in2[119];
    assign P[5] = in1[119] ^ in2[119];
    assign G[6] = in1[118] & in2[118];
    assign P[6] = in1[118] ^ in2[118];
    assign G[7] = in1[117] & in2[117];
    assign P[7] = in1[117] ^ in2[117];
    assign G[8] = in1[116] & in2[116];
    assign P[8] = in1[116] ^ in2[116];
    assign G[9] = in1[115] & in2[115];
    assign P[9] = in1[115] ^ in2[115];
    assign G[10] = in1[114] & in2[114];
    assign P[10] = in1[114] ^ in2[114];
    assign G[11] = in1[113] & in2[113];
    assign P[11] = in1[113] ^ in2[113];
    assign G[12] = in1[112] & in2[112];
    assign P[12] = in1[112] ^ in2[112];
    assign G[13] = in1[111] & in2[111];
    assign P[13] = in1[111] ^ in2[111];
    assign G[14] = in1[110] & in2[110];
    assign P[14] = in1[110] ^ in2[110];
    assign G[15] = in1[109] & in2[109];
    assign P[15] = in1[109] ^ in2[109];
    assign G[16] = in1[108] & in2[108];
    assign P[16] = in1[108] ^ in2[108];
    assign G[17] = in1[107] & in2[107];
    assign P[17] = in1[107] ^ in2[107];
    assign G[18] = in1[106] & in2[106];
    assign P[18] = in1[106] ^ in2[106];
    assign G[19] = in1[105] & in2[105];
    assign P[19] = in1[105] ^ in2[105];
    assign G[20] = in1[104] & in2[104];
    assign P[20] = in1[104] ^ in2[104];
    assign G[21] = in1[103] & in2[103];
    assign P[21] = in1[103] ^ in2[103];
    assign G[22] = in1[102] & in2[102];
    assign P[22] = in1[102] ^ in2[102];
    assign G[23] = in1[101] & in2[101];
    assign P[23] = in1[101] ^ in2[101];
    assign G[24] = in1[100] & in2[100];
    assign P[24] = in1[100] ^ in2[100];
    assign G[25] = in1[99] & in2[99];
    assign P[25] = in1[99] ^ in2[99];
    assign G[26] = in1[98] & in2[98];
    assign P[26] = in1[98] ^ in2[98];
    assign G[27] = in1[97] & in2[97];
    assign P[27] = in1[97] ^ in2[97];
    assign G[28] = in1[96] & in2[96];
    assign P[28] = in1[96] ^ in2[96];
    assign G[29] = in1[95] & in2[95];
    assign P[29] = in1[95] ^ in2[95];
    assign G[30] = in1[94] & in2[94];
    assign P[30] = in1[94] ^ in2[94];
    assign G[31] = in1[93] & in2[93];
    assign P[31] = in1[93] ^ in2[93];
    assign G[32] = in1[92] & in2[92];
    assign P[32] = in1[92] ^ in2[92];
    assign G[33] = in1[91] & in2[91];
    assign P[33] = in1[91] ^ in2[91];
    assign G[34] = in1[90] & in2[90];
    assign P[34] = in1[90] ^ in2[90];
    assign G[35] = in1[89] & in2[89];
    assign P[35] = in1[89] ^ in2[89];
    assign G[36] = in1[88] & in2[88];
    assign P[36] = in1[88] ^ in2[88];
    assign G[37] = in1[87] & in2[87];
    assign P[37] = in1[87] ^ in2[87];
    assign G[38] = in1[86] & in2[86];
    assign P[38] = in1[86] ^ in2[86];
    assign G[39] = in1[85] & in2[85];
    assign P[39] = in1[85] ^ in2[85];
    assign G[40] = in1[84] & in2[84];
    assign P[40] = in1[84] ^ in2[84];
    assign G[41] = in1[83] & in2[83];
    assign P[41] = in1[83] ^ in2[83];
    assign G[42] = in1[82] & in2[82];
    assign P[42] = in1[82] ^ in2[82];
    assign G[43] = in1[81] & in2[81];
    assign P[43] = in1[81] ^ in2[81];
    assign G[44] = in1[80] & in2[80];
    assign P[44] = in1[80] ^ in2[80];
    assign G[45] = in1[79] & in2[79];
    assign P[45] = in1[79] ^ in2[79];
    assign G[46] = in1[78] & in2[78];
    assign P[46] = in1[78] ^ in2[78];
    assign G[47] = in1[77] & in2[77];
    assign P[47] = in1[77] ^ in2[77];
    assign G[48] = in1[76] & in2[76];
    assign P[48] = in1[76] ^ in2[76];
    assign G[49] = in1[75] & in2[75];
    assign P[49] = in1[75] ^ in2[75];
    assign G[50] = in1[74] & in2[74];
    assign P[50] = in1[74] ^ in2[74];
    assign G[51] = in1[73] & in2[73];
    assign P[51] = in1[73] ^ in2[73];
    assign G[52] = in1[72] & in2[72];
    assign P[52] = in1[72] ^ in2[72];
    assign G[53] = in1[71] & in2[71];
    assign P[53] = in1[71] ^ in2[71];
    assign G[54] = in1[70] & in2[70];
    assign P[54] = in1[70] ^ in2[70];
    assign G[55] = in1[69] & in2[69];
    assign P[55] = in1[69] ^ in2[69];
    assign G[56] = in1[68] & in2[68];
    assign P[56] = in1[68] ^ in2[68];
    assign G[57] = in1[67] & in2[67];
    assign P[57] = in1[67] ^ in2[67];
    assign G[58] = in1[66] & in2[66];
    assign P[58] = in1[66] ^ in2[66];
    assign G[59] = in1[65] & in2[65];
    assign P[59] = in1[65] ^ in2[65];
    assign G[60] = in1[64] & in2[64];
    assign P[60] = in1[64] ^ in2[64];
    assign G[61] = in1[63] & in2[63];
    assign P[61] = in1[63] ^ in2[63];
    assign G[62] = in1[62] & in2[62];
    assign P[62] = in1[62] ^ in2[62];
    assign G[63] = in1[61] & in2[61];
    assign P[63] = in1[61] ^ in2[61];
    assign G[64] = in1[60] & in2[60];
    assign P[64] = in1[60] ^ in2[60];
    assign G[65] = in1[59] & in2[59];
    assign P[65] = in1[59] ^ in2[59];
    assign G[66] = in1[58] & in2[58];
    assign P[66] = in1[58] ^ in2[58];
    assign G[67] = in1[57] & in2[57];
    assign P[67] = in1[57] ^ in2[57];
    assign G[68] = in1[56] & in2[56];
    assign P[68] = in1[56] ^ in2[56];
    assign G[69] = in1[55] & in2[55];
    assign P[69] = in1[55] ^ in2[55];
    assign G[70] = in1[54] & in2[54];
    assign P[70] = in1[54] ^ in2[54];
    assign G[71] = in1[53] & in2[53];
    assign P[71] = in1[53] ^ in2[53];
    assign G[72] = in1[52] & in2[52];
    assign P[72] = in1[52] ^ in2[52];
    assign G[73] = in1[51] & in2[51];
    assign P[73] = in1[51] ^ in2[51];
    assign G[74] = in1[50] & in2[50];
    assign P[74] = in1[50] ^ in2[50];
    assign G[75] = in1[49] & in2[49];
    assign P[75] = in1[49] ^ in2[49];
    assign G[76] = in1[48] & in2[48];
    assign P[76] = in1[48] ^ in2[48];
    assign G[77] = in1[47] & in2[47];
    assign P[77] = in1[47] ^ in2[47];
    assign G[78] = in1[46] & in2[46];
    assign P[78] = in1[46] ^ in2[46];
    assign G[79] = in1[45] & in2[45];
    assign P[79] = in1[45] ^ in2[45];
    assign G[80] = in1[44] & in2[44];
    assign P[80] = in1[44] ^ in2[44];
    assign G[81] = in1[43] & in2[43];
    assign P[81] = in1[43] ^ in2[43];
    assign G[82] = in1[42] & in2[42];
    assign P[82] = in1[42] ^ in2[42];
    assign G[83] = in1[41] & in2[41];
    assign P[83] = in1[41] ^ in2[41];
    assign G[84] = in1[40] & in2[40];
    assign P[84] = in1[40] ^ in2[40];
    assign G[85] = in1[39] & in2[39];
    assign P[85] = in1[39] ^ in2[39];
    assign G[86] = in1[38] & in2[38];
    assign P[86] = in1[38] ^ in2[38];
    assign G[87] = in1[37] & in2[37];
    assign P[87] = in1[37] ^ in2[37];
    assign G[88] = in1[36] & in2[36];
    assign P[88] = in1[36] ^ in2[36];
    assign G[89] = in1[35] & in2[35];
    assign P[89] = in1[35] ^ in2[35];
    assign G[90] = in1[34] & in2[34];
    assign P[90] = in1[34] ^ in2[34];
    assign G[91] = in1[33] & in2[33];
    assign P[91] = in1[33] ^ in2[33];
    assign G[92] = in1[32] & in2[32];
    assign P[92] = in1[32] ^ in2[32];
    assign G[93] = in1[31] & in2[31];
    assign P[93] = in1[31] ^ in2[31];
    assign G[94] = in1[30] & in2[30];
    assign P[94] = in1[30] ^ in2[30];
    assign G[95] = in1[29] & in2[29];
    assign P[95] = in1[29] ^ in2[29];
    assign G[96] = in1[28] & in2[28];
    assign P[96] = in1[28] ^ in2[28];
    assign G[97] = in1[27] & in2[27];
    assign P[97] = in1[27] ^ in2[27];
    assign G[98] = in1[26] & in2[26];
    assign P[98] = in1[26] ^ in2[26];
    assign G[99] = in1[25] & in2[25];
    assign P[99] = in1[25] ^ in2[25];
    assign G[100] = in1[24] & in2[24];
    assign P[100] = in1[24] ^ in2[24];
    assign G[101] = in1[23] & in2[23];
    assign P[101] = in1[23] ^ in2[23];
    assign G[102] = in1[22] & in2[22];
    assign P[102] = in1[22] ^ in2[22];
    assign G[103] = in1[21] & in2[21];
    assign P[103] = in1[21] ^ in2[21];
    assign G[104] = in1[20] & in2[20];
    assign P[104] = in1[20] ^ in2[20];
    assign G[105] = in1[19] & in2[19];
    assign P[105] = in1[19] ^ in2[19];
    assign G[106] = in1[18] & in2[18];
    assign P[106] = in1[18] ^ in2[18];
    assign G[107] = in1[17] & in2[17];
    assign P[107] = in1[17] ^ in2[17];
    assign G[108] = in1[16] & in2[16];
    assign P[108] = in1[16] ^ in2[16];
    assign G[109] = in1[15] & in2[15];
    assign P[109] = in1[15] ^ in2[15];
    assign G[110] = in1[14] & in2[14];
    assign P[110] = in1[14] ^ in2[14];
    assign G[111] = in1[13] & in2[13];
    assign P[111] = in1[13] ^ in2[13];
    assign G[112] = in1[12] & in2[12];
    assign P[112] = in1[12] ^ in2[12];
    assign G[113] = in1[11] & in2[11];
    assign P[113] = in1[11] ^ in2[11];
    assign G[114] = in1[10] & in2[10];
    assign P[114] = in1[10] ^ in2[10];
    assign G[115] = in1[9] & in2[9];
    assign P[115] = in1[9] ^ in2[9];
    assign G[116] = in1[8] & in2[8];
    assign P[116] = in1[8] ^ in2[8];
    assign G[117] = in1[7] & in2[7];
    assign P[117] = in1[7] ^ in2[7];
    assign G[118] = in1[6] & in2[6];
    assign P[118] = in1[6] ^ in2[6];
    assign G[119] = in1[5] & in2[5];
    assign P[119] = in1[5] ^ in2[5];
    assign G[120] = in1[4] & in2[4];
    assign P[120] = in1[4] ^ in2[4];
    assign G[121] = in1[3] & in2[3];
    assign P[121] = in1[3] ^ in2[3];
    assign G[122] = in1[2] & in2[2];
    assign P[122] = in1[2] ^ in2[2];
    assign G[123] = in1[1] & in2[1];
    assign P[123] = in1[1] ^ in2[1];
    assign G[124] = in1[0] & in2[0];
    assign P[124] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign cout = G[124] | (P[124] & C[124]);
    assign sum = P ^ C;
endmodule

module CLA_124(output [123:0] sum, output cout, input [123:0] in1, input [123:0] in2);

    wire[123:0] G;
    wire[123:0] C;
    wire[123:0] P;

    assign G[0] = in1[123] & in2[123];
    assign P[0] = in1[123] ^ in2[123];
    assign G[1] = in1[122] & in2[122];
    assign P[1] = in1[122] ^ in2[122];
    assign G[2] = in1[121] & in2[121];
    assign P[2] = in1[121] ^ in2[121];
    assign G[3] = in1[120] & in2[120];
    assign P[3] = in1[120] ^ in2[120];
    assign G[4] = in1[119] & in2[119];
    assign P[4] = in1[119] ^ in2[119];
    assign G[5] = in1[118] & in2[118];
    assign P[5] = in1[118] ^ in2[118];
    assign G[6] = in1[117] & in2[117];
    assign P[6] = in1[117] ^ in2[117];
    assign G[7] = in1[116] & in2[116];
    assign P[7] = in1[116] ^ in2[116];
    assign G[8] = in1[115] & in2[115];
    assign P[8] = in1[115] ^ in2[115];
    assign G[9] = in1[114] & in2[114];
    assign P[9] = in1[114] ^ in2[114];
    assign G[10] = in1[113] & in2[113];
    assign P[10] = in1[113] ^ in2[113];
    assign G[11] = in1[112] & in2[112];
    assign P[11] = in1[112] ^ in2[112];
    assign G[12] = in1[111] & in2[111];
    assign P[12] = in1[111] ^ in2[111];
    assign G[13] = in1[110] & in2[110];
    assign P[13] = in1[110] ^ in2[110];
    assign G[14] = in1[109] & in2[109];
    assign P[14] = in1[109] ^ in2[109];
    assign G[15] = in1[108] & in2[108];
    assign P[15] = in1[108] ^ in2[108];
    assign G[16] = in1[107] & in2[107];
    assign P[16] = in1[107] ^ in2[107];
    assign G[17] = in1[106] & in2[106];
    assign P[17] = in1[106] ^ in2[106];
    assign G[18] = in1[105] & in2[105];
    assign P[18] = in1[105] ^ in2[105];
    assign G[19] = in1[104] & in2[104];
    assign P[19] = in1[104] ^ in2[104];
    assign G[20] = in1[103] & in2[103];
    assign P[20] = in1[103] ^ in2[103];
    assign G[21] = in1[102] & in2[102];
    assign P[21] = in1[102] ^ in2[102];
    assign G[22] = in1[101] & in2[101];
    assign P[22] = in1[101] ^ in2[101];
    assign G[23] = in1[100] & in2[100];
    assign P[23] = in1[100] ^ in2[100];
    assign G[24] = in1[99] & in2[99];
    assign P[24] = in1[99] ^ in2[99];
    assign G[25] = in1[98] & in2[98];
    assign P[25] = in1[98] ^ in2[98];
    assign G[26] = in1[97] & in2[97];
    assign P[26] = in1[97] ^ in2[97];
    assign G[27] = in1[96] & in2[96];
    assign P[27] = in1[96] ^ in2[96];
    assign G[28] = in1[95] & in2[95];
    assign P[28] = in1[95] ^ in2[95];
    assign G[29] = in1[94] & in2[94];
    assign P[29] = in1[94] ^ in2[94];
    assign G[30] = in1[93] & in2[93];
    assign P[30] = in1[93] ^ in2[93];
    assign G[31] = in1[92] & in2[92];
    assign P[31] = in1[92] ^ in2[92];
    assign G[32] = in1[91] & in2[91];
    assign P[32] = in1[91] ^ in2[91];
    assign G[33] = in1[90] & in2[90];
    assign P[33] = in1[90] ^ in2[90];
    assign G[34] = in1[89] & in2[89];
    assign P[34] = in1[89] ^ in2[89];
    assign G[35] = in1[88] & in2[88];
    assign P[35] = in1[88] ^ in2[88];
    assign G[36] = in1[87] & in2[87];
    assign P[36] = in1[87] ^ in2[87];
    assign G[37] = in1[86] & in2[86];
    assign P[37] = in1[86] ^ in2[86];
    assign G[38] = in1[85] & in2[85];
    assign P[38] = in1[85] ^ in2[85];
    assign G[39] = in1[84] & in2[84];
    assign P[39] = in1[84] ^ in2[84];
    assign G[40] = in1[83] & in2[83];
    assign P[40] = in1[83] ^ in2[83];
    assign G[41] = in1[82] & in2[82];
    assign P[41] = in1[82] ^ in2[82];
    assign G[42] = in1[81] & in2[81];
    assign P[42] = in1[81] ^ in2[81];
    assign G[43] = in1[80] & in2[80];
    assign P[43] = in1[80] ^ in2[80];
    assign G[44] = in1[79] & in2[79];
    assign P[44] = in1[79] ^ in2[79];
    assign G[45] = in1[78] & in2[78];
    assign P[45] = in1[78] ^ in2[78];
    assign G[46] = in1[77] & in2[77];
    assign P[46] = in1[77] ^ in2[77];
    assign G[47] = in1[76] & in2[76];
    assign P[47] = in1[76] ^ in2[76];
    assign G[48] = in1[75] & in2[75];
    assign P[48] = in1[75] ^ in2[75];
    assign G[49] = in1[74] & in2[74];
    assign P[49] = in1[74] ^ in2[74];
    assign G[50] = in1[73] & in2[73];
    assign P[50] = in1[73] ^ in2[73];
    assign G[51] = in1[72] & in2[72];
    assign P[51] = in1[72] ^ in2[72];
    assign G[52] = in1[71] & in2[71];
    assign P[52] = in1[71] ^ in2[71];
    assign G[53] = in1[70] & in2[70];
    assign P[53] = in1[70] ^ in2[70];
    assign G[54] = in1[69] & in2[69];
    assign P[54] = in1[69] ^ in2[69];
    assign G[55] = in1[68] & in2[68];
    assign P[55] = in1[68] ^ in2[68];
    assign G[56] = in1[67] & in2[67];
    assign P[56] = in1[67] ^ in2[67];
    assign G[57] = in1[66] & in2[66];
    assign P[57] = in1[66] ^ in2[66];
    assign G[58] = in1[65] & in2[65];
    assign P[58] = in1[65] ^ in2[65];
    assign G[59] = in1[64] & in2[64];
    assign P[59] = in1[64] ^ in2[64];
    assign G[60] = in1[63] & in2[63];
    assign P[60] = in1[63] ^ in2[63];
    assign G[61] = in1[62] & in2[62];
    assign P[61] = in1[62] ^ in2[62];
    assign G[62] = in1[61] & in2[61];
    assign P[62] = in1[61] ^ in2[61];
    assign G[63] = in1[60] & in2[60];
    assign P[63] = in1[60] ^ in2[60];
    assign G[64] = in1[59] & in2[59];
    assign P[64] = in1[59] ^ in2[59];
    assign G[65] = in1[58] & in2[58];
    assign P[65] = in1[58] ^ in2[58];
    assign G[66] = in1[57] & in2[57];
    assign P[66] = in1[57] ^ in2[57];
    assign G[67] = in1[56] & in2[56];
    assign P[67] = in1[56] ^ in2[56];
    assign G[68] = in1[55] & in2[55];
    assign P[68] = in1[55] ^ in2[55];
    assign G[69] = in1[54] & in2[54];
    assign P[69] = in1[54] ^ in2[54];
    assign G[70] = in1[53] & in2[53];
    assign P[70] = in1[53] ^ in2[53];
    assign G[71] = in1[52] & in2[52];
    assign P[71] = in1[52] ^ in2[52];
    assign G[72] = in1[51] & in2[51];
    assign P[72] = in1[51] ^ in2[51];
    assign G[73] = in1[50] & in2[50];
    assign P[73] = in1[50] ^ in2[50];
    assign G[74] = in1[49] & in2[49];
    assign P[74] = in1[49] ^ in2[49];
    assign G[75] = in1[48] & in2[48];
    assign P[75] = in1[48] ^ in2[48];
    assign G[76] = in1[47] & in2[47];
    assign P[76] = in1[47] ^ in2[47];
    assign G[77] = in1[46] & in2[46];
    assign P[77] = in1[46] ^ in2[46];
    assign G[78] = in1[45] & in2[45];
    assign P[78] = in1[45] ^ in2[45];
    assign G[79] = in1[44] & in2[44];
    assign P[79] = in1[44] ^ in2[44];
    assign G[80] = in1[43] & in2[43];
    assign P[80] = in1[43] ^ in2[43];
    assign G[81] = in1[42] & in2[42];
    assign P[81] = in1[42] ^ in2[42];
    assign G[82] = in1[41] & in2[41];
    assign P[82] = in1[41] ^ in2[41];
    assign G[83] = in1[40] & in2[40];
    assign P[83] = in1[40] ^ in2[40];
    assign G[84] = in1[39] & in2[39];
    assign P[84] = in1[39] ^ in2[39];
    assign G[85] = in1[38] & in2[38];
    assign P[85] = in1[38] ^ in2[38];
    assign G[86] = in1[37] & in2[37];
    assign P[86] = in1[37] ^ in2[37];
    assign G[87] = in1[36] & in2[36];
    assign P[87] = in1[36] ^ in2[36];
    assign G[88] = in1[35] & in2[35];
    assign P[88] = in1[35] ^ in2[35];
    assign G[89] = in1[34] & in2[34];
    assign P[89] = in1[34] ^ in2[34];
    assign G[90] = in1[33] & in2[33];
    assign P[90] = in1[33] ^ in2[33];
    assign G[91] = in1[32] & in2[32];
    assign P[91] = in1[32] ^ in2[32];
    assign G[92] = in1[31] & in2[31];
    assign P[92] = in1[31] ^ in2[31];
    assign G[93] = in1[30] & in2[30];
    assign P[93] = in1[30] ^ in2[30];
    assign G[94] = in1[29] & in2[29];
    assign P[94] = in1[29] ^ in2[29];
    assign G[95] = in1[28] & in2[28];
    assign P[95] = in1[28] ^ in2[28];
    assign G[96] = in1[27] & in2[27];
    assign P[96] = in1[27] ^ in2[27];
    assign G[97] = in1[26] & in2[26];
    assign P[97] = in1[26] ^ in2[26];
    assign G[98] = in1[25] & in2[25];
    assign P[98] = in1[25] ^ in2[25];
    assign G[99] = in1[24] & in2[24];
    assign P[99] = in1[24] ^ in2[24];
    assign G[100] = in1[23] & in2[23];
    assign P[100] = in1[23] ^ in2[23];
    assign G[101] = in1[22] & in2[22];
    assign P[101] = in1[22] ^ in2[22];
    assign G[102] = in1[21] & in2[21];
    assign P[102] = in1[21] ^ in2[21];
    assign G[103] = in1[20] & in2[20];
    assign P[103] = in1[20] ^ in2[20];
    assign G[104] = in1[19] & in2[19];
    assign P[104] = in1[19] ^ in2[19];
    assign G[105] = in1[18] & in2[18];
    assign P[105] = in1[18] ^ in2[18];
    assign G[106] = in1[17] & in2[17];
    assign P[106] = in1[17] ^ in2[17];
    assign G[107] = in1[16] & in2[16];
    assign P[107] = in1[16] ^ in2[16];
    assign G[108] = in1[15] & in2[15];
    assign P[108] = in1[15] ^ in2[15];
    assign G[109] = in1[14] & in2[14];
    assign P[109] = in1[14] ^ in2[14];
    assign G[110] = in1[13] & in2[13];
    assign P[110] = in1[13] ^ in2[13];
    assign G[111] = in1[12] & in2[12];
    assign P[111] = in1[12] ^ in2[12];
    assign G[112] = in1[11] & in2[11];
    assign P[112] = in1[11] ^ in2[11];
    assign G[113] = in1[10] & in2[10];
    assign P[113] = in1[10] ^ in2[10];
    assign G[114] = in1[9] & in2[9];
    assign P[114] = in1[9] ^ in2[9];
    assign G[115] = in1[8] & in2[8];
    assign P[115] = in1[8] ^ in2[8];
    assign G[116] = in1[7] & in2[7];
    assign P[116] = in1[7] ^ in2[7];
    assign G[117] = in1[6] & in2[6];
    assign P[117] = in1[6] ^ in2[6];
    assign G[118] = in1[5] & in2[5];
    assign P[118] = in1[5] ^ in2[5];
    assign G[119] = in1[4] & in2[4];
    assign P[119] = in1[4] ^ in2[4];
    assign G[120] = in1[3] & in2[3];
    assign P[120] = in1[3] ^ in2[3];
    assign G[121] = in1[2] & in2[2];
    assign P[121] = in1[2] ^ in2[2];
    assign G[122] = in1[1] & in2[1];
    assign P[122] = in1[1] ^ in2[1];
    assign G[123] = in1[0] & in2[0];
    assign P[123] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign cout = G[123] | (P[123] & C[123]);
    assign sum = P ^ C;
endmodule

module CLA_123(output [122:0] sum, output cout, input [122:0] in1, input [122:0] in2);

    wire[122:0] G;
    wire[122:0] C;
    wire[122:0] P;

    assign G[0] = in1[122] & in2[122];
    assign P[0] = in1[122] ^ in2[122];
    assign G[1] = in1[121] & in2[121];
    assign P[1] = in1[121] ^ in2[121];
    assign G[2] = in1[120] & in2[120];
    assign P[2] = in1[120] ^ in2[120];
    assign G[3] = in1[119] & in2[119];
    assign P[3] = in1[119] ^ in2[119];
    assign G[4] = in1[118] & in2[118];
    assign P[4] = in1[118] ^ in2[118];
    assign G[5] = in1[117] & in2[117];
    assign P[5] = in1[117] ^ in2[117];
    assign G[6] = in1[116] & in2[116];
    assign P[6] = in1[116] ^ in2[116];
    assign G[7] = in1[115] & in2[115];
    assign P[7] = in1[115] ^ in2[115];
    assign G[8] = in1[114] & in2[114];
    assign P[8] = in1[114] ^ in2[114];
    assign G[9] = in1[113] & in2[113];
    assign P[9] = in1[113] ^ in2[113];
    assign G[10] = in1[112] & in2[112];
    assign P[10] = in1[112] ^ in2[112];
    assign G[11] = in1[111] & in2[111];
    assign P[11] = in1[111] ^ in2[111];
    assign G[12] = in1[110] & in2[110];
    assign P[12] = in1[110] ^ in2[110];
    assign G[13] = in1[109] & in2[109];
    assign P[13] = in1[109] ^ in2[109];
    assign G[14] = in1[108] & in2[108];
    assign P[14] = in1[108] ^ in2[108];
    assign G[15] = in1[107] & in2[107];
    assign P[15] = in1[107] ^ in2[107];
    assign G[16] = in1[106] & in2[106];
    assign P[16] = in1[106] ^ in2[106];
    assign G[17] = in1[105] & in2[105];
    assign P[17] = in1[105] ^ in2[105];
    assign G[18] = in1[104] & in2[104];
    assign P[18] = in1[104] ^ in2[104];
    assign G[19] = in1[103] & in2[103];
    assign P[19] = in1[103] ^ in2[103];
    assign G[20] = in1[102] & in2[102];
    assign P[20] = in1[102] ^ in2[102];
    assign G[21] = in1[101] & in2[101];
    assign P[21] = in1[101] ^ in2[101];
    assign G[22] = in1[100] & in2[100];
    assign P[22] = in1[100] ^ in2[100];
    assign G[23] = in1[99] & in2[99];
    assign P[23] = in1[99] ^ in2[99];
    assign G[24] = in1[98] & in2[98];
    assign P[24] = in1[98] ^ in2[98];
    assign G[25] = in1[97] & in2[97];
    assign P[25] = in1[97] ^ in2[97];
    assign G[26] = in1[96] & in2[96];
    assign P[26] = in1[96] ^ in2[96];
    assign G[27] = in1[95] & in2[95];
    assign P[27] = in1[95] ^ in2[95];
    assign G[28] = in1[94] & in2[94];
    assign P[28] = in1[94] ^ in2[94];
    assign G[29] = in1[93] & in2[93];
    assign P[29] = in1[93] ^ in2[93];
    assign G[30] = in1[92] & in2[92];
    assign P[30] = in1[92] ^ in2[92];
    assign G[31] = in1[91] & in2[91];
    assign P[31] = in1[91] ^ in2[91];
    assign G[32] = in1[90] & in2[90];
    assign P[32] = in1[90] ^ in2[90];
    assign G[33] = in1[89] & in2[89];
    assign P[33] = in1[89] ^ in2[89];
    assign G[34] = in1[88] & in2[88];
    assign P[34] = in1[88] ^ in2[88];
    assign G[35] = in1[87] & in2[87];
    assign P[35] = in1[87] ^ in2[87];
    assign G[36] = in1[86] & in2[86];
    assign P[36] = in1[86] ^ in2[86];
    assign G[37] = in1[85] & in2[85];
    assign P[37] = in1[85] ^ in2[85];
    assign G[38] = in1[84] & in2[84];
    assign P[38] = in1[84] ^ in2[84];
    assign G[39] = in1[83] & in2[83];
    assign P[39] = in1[83] ^ in2[83];
    assign G[40] = in1[82] & in2[82];
    assign P[40] = in1[82] ^ in2[82];
    assign G[41] = in1[81] & in2[81];
    assign P[41] = in1[81] ^ in2[81];
    assign G[42] = in1[80] & in2[80];
    assign P[42] = in1[80] ^ in2[80];
    assign G[43] = in1[79] & in2[79];
    assign P[43] = in1[79] ^ in2[79];
    assign G[44] = in1[78] & in2[78];
    assign P[44] = in1[78] ^ in2[78];
    assign G[45] = in1[77] & in2[77];
    assign P[45] = in1[77] ^ in2[77];
    assign G[46] = in1[76] & in2[76];
    assign P[46] = in1[76] ^ in2[76];
    assign G[47] = in1[75] & in2[75];
    assign P[47] = in1[75] ^ in2[75];
    assign G[48] = in1[74] & in2[74];
    assign P[48] = in1[74] ^ in2[74];
    assign G[49] = in1[73] & in2[73];
    assign P[49] = in1[73] ^ in2[73];
    assign G[50] = in1[72] & in2[72];
    assign P[50] = in1[72] ^ in2[72];
    assign G[51] = in1[71] & in2[71];
    assign P[51] = in1[71] ^ in2[71];
    assign G[52] = in1[70] & in2[70];
    assign P[52] = in1[70] ^ in2[70];
    assign G[53] = in1[69] & in2[69];
    assign P[53] = in1[69] ^ in2[69];
    assign G[54] = in1[68] & in2[68];
    assign P[54] = in1[68] ^ in2[68];
    assign G[55] = in1[67] & in2[67];
    assign P[55] = in1[67] ^ in2[67];
    assign G[56] = in1[66] & in2[66];
    assign P[56] = in1[66] ^ in2[66];
    assign G[57] = in1[65] & in2[65];
    assign P[57] = in1[65] ^ in2[65];
    assign G[58] = in1[64] & in2[64];
    assign P[58] = in1[64] ^ in2[64];
    assign G[59] = in1[63] & in2[63];
    assign P[59] = in1[63] ^ in2[63];
    assign G[60] = in1[62] & in2[62];
    assign P[60] = in1[62] ^ in2[62];
    assign G[61] = in1[61] & in2[61];
    assign P[61] = in1[61] ^ in2[61];
    assign G[62] = in1[60] & in2[60];
    assign P[62] = in1[60] ^ in2[60];
    assign G[63] = in1[59] & in2[59];
    assign P[63] = in1[59] ^ in2[59];
    assign G[64] = in1[58] & in2[58];
    assign P[64] = in1[58] ^ in2[58];
    assign G[65] = in1[57] & in2[57];
    assign P[65] = in1[57] ^ in2[57];
    assign G[66] = in1[56] & in2[56];
    assign P[66] = in1[56] ^ in2[56];
    assign G[67] = in1[55] & in2[55];
    assign P[67] = in1[55] ^ in2[55];
    assign G[68] = in1[54] & in2[54];
    assign P[68] = in1[54] ^ in2[54];
    assign G[69] = in1[53] & in2[53];
    assign P[69] = in1[53] ^ in2[53];
    assign G[70] = in1[52] & in2[52];
    assign P[70] = in1[52] ^ in2[52];
    assign G[71] = in1[51] & in2[51];
    assign P[71] = in1[51] ^ in2[51];
    assign G[72] = in1[50] & in2[50];
    assign P[72] = in1[50] ^ in2[50];
    assign G[73] = in1[49] & in2[49];
    assign P[73] = in1[49] ^ in2[49];
    assign G[74] = in1[48] & in2[48];
    assign P[74] = in1[48] ^ in2[48];
    assign G[75] = in1[47] & in2[47];
    assign P[75] = in1[47] ^ in2[47];
    assign G[76] = in1[46] & in2[46];
    assign P[76] = in1[46] ^ in2[46];
    assign G[77] = in1[45] & in2[45];
    assign P[77] = in1[45] ^ in2[45];
    assign G[78] = in1[44] & in2[44];
    assign P[78] = in1[44] ^ in2[44];
    assign G[79] = in1[43] & in2[43];
    assign P[79] = in1[43] ^ in2[43];
    assign G[80] = in1[42] & in2[42];
    assign P[80] = in1[42] ^ in2[42];
    assign G[81] = in1[41] & in2[41];
    assign P[81] = in1[41] ^ in2[41];
    assign G[82] = in1[40] & in2[40];
    assign P[82] = in1[40] ^ in2[40];
    assign G[83] = in1[39] & in2[39];
    assign P[83] = in1[39] ^ in2[39];
    assign G[84] = in1[38] & in2[38];
    assign P[84] = in1[38] ^ in2[38];
    assign G[85] = in1[37] & in2[37];
    assign P[85] = in1[37] ^ in2[37];
    assign G[86] = in1[36] & in2[36];
    assign P[86] = in1[36] ^ in2[36];
    assign G[87] = in1[35] & in2[35];
    assign P[87] = in1[35] ^ in2[35];
    assign G[88] = in1[34] & in2[34];
    assign P[88] = in1[34] ^ in2[34];
    assign G[89] = in1[33] & in2[33];
    assign P[89] = in1[33] ^ in2[33];
    assign G[90] = in1[32] & in2[32];
    assign P[90] = in1[32] ^ in2[32];
    assign G[91] = in1[31] & in2[31];
    assign P[91] = in1[31] ^ in2[31];
    assign G[92] = in1[30] & in2[30];
    assign P[92] = in1[30] ^ in2[30];
    assign G[93] = in1[29] & in2[29];
    assign P[93] = in1[29] ^ in2[29];
    assign G[94] = in1[28] & in2[28];
    assign P[94] = in1[28] ^ in2[28];
    assign G[95] = in1[27] & in2[27];
    assign P[95] = in1[27] ^ in2[27];
    assign G[96] = in1[26] & in2[26];
    assign P[96] = in1[26] ^ in2[26];
    assign G[97] = in1[25] & in2[25];
    assign P[97] = in1[25] ^ in2[25];
    assign G[98] = in1[24] & in2[24];
    assign P[98] = in1[24] ^ in2[24];
    assign G[99] = in1[23] & in2[23];
    assign P[99] = in1[23] ^ in2[23];
    assign G[100] = in1[22] & in2[22];
    assign P[100] = in1[22] ^ in2[22];
    assign G[101] = in1[21] & in2[21];
    assign P[101] = in1[21] ^ in2[21];
    assign G[102] = in1[20] & in2[20];
    assign P[102] = in1[20] ^ in2[20];
    assign G[103] = in1[19] & in2[19];
    assign P[103] = in1[19] ^ in2[19];
    assign G[104] = in1[18] & in2[18];
    assign P[104] = in1[18] ^ in2[18];
    assign G[105] = in1[17] & in2[17];
    assign P[105] = in1[17] ^ in2[17];
    assign G[106] = in1[16] & in2[16];
    assign P[106] = in1[16] ^ in2[16];
    assign G[107] = in1[15] & in2[15];
    assign P[107] = in1[15] ^ in2[15];
    assign G[108] = in1[14] & in2[14];
    assign P[108] = in1[14] ^ in2[14];
    assign G[109] = in1[13] & in2[13];
    assign P[109] = in1[13] ^ in2[13];
    assign G[110] = in1[12] & in2[12];
    assign P[110] = in1[12] ^ in2[12];
    assign G[111] = in1[11] & in2[11];
    assign P[111] = in1[11] ^ in2[11];
    assign G[112] = in1[10] & in2[10];
    assign P[112] = in1[10] ^ in2[10];
    assign G[113] = in1[9] & in2[9];
    assign P[113] = in1[9] ^ in2[9];
    assign G[114] = in1[8] & in2[8];
    assign P[114] = in1[8] ^ in2[8];
    assign G[115] = in1[7] & in2[7];
    assign P[115] = in1[7] ^ in2[7];
    assign G[116] = in1[6] & in2[6];
    assign P[116] = in1[6] ^ in2[6];
    assign G[117] = in1[5] & in2[5];
    assign P[117] = in1[5] ^ in2[5];
    assign G[118] = in1[4] & in2[4];
    assign P[118] = in1[4] ^ in2[4];
    assign G[119] = in1[3] & in2[3];
    assign P[119] = in1[3] ^ in2[3];
    assign G[120] = in1[2] & in2[2];
    assign P[120] = in1[2] ^ in2[2];
    assign G[121] = in1[1] & in2[1];
    assign P[121] = in1[1] ^ in2[1];
    assign G[122] = in1[0] & in2[0];
    assign P[122] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign cout = G[122] | (P[122] & C[122]);
    assign sum = P ^ C;
endmodule

module CLA_122(output [121:0] sum, output cout, input [121:0] in1, input [121:0] in2);

    wire[121:0] G;
    wire[121:0] C;
    wire[121:0] P;

    assign G[0] = in1[121] & in2[121];
    assign P[0] = in1[121] ^ in2[121];
    assign G[1] = in1[120] & in2[120];
    assign P[1] = in1[120] ^ in2[120];
    assign G[2] = in1[119] & in2[119];
    assign P[2] = in1[119] ^ in2[119];
    assign G[3] = in1[118] & in2[118];
    assign P[3] = in1[118] ^ in2[118];
    assign G[4] = in1[117] & in2[117];
    assign P[4] = in1[117] ^ in2[117];
    assign G[5] = in1[116] & in2[116];
    assign P[5] = in1[116] ^ in2[116];
    assign G[6] = in1[115] & in2[115];
    assign P[6] = in1[115] ^ in2[115];
    assign G[7] = in1[114] & in2[114];
    assign P[7] = in1[114] ^ in2[114];
    assign G[8] = in1[113] & in2[113];
    assign P[8] = in1[113] ^ in2[113];
    assign G[9] = in1[112] & in2[112];
    assign P[9] = in1[112] ^ in2[112];
    assign G[10] = in1[111] & in2[111];
    assign P[10] = in1[111] ^ in2[111];
    assign G[11] = in1[110] & in2[110];
    assign P[11] = in1[110] ^ in2[110];
    assign G[12] = in1[109] & in2[109];
    assign P[12] = in1[109] ^ in2[109];
    assign G[13] = in1[108] & in2[108];
    assign P[13] = in1[108] ^ in2[108];
    assign G[14] = in1[107] & in2[107];
    assign P[14] = in1[107] ^ in2[107];
    assign G[15] = in1[106] & in2[106];
    assign P[15] = in1[106] ^ in2[106];
    assign G[16] = in1[105] & in2[105];
    assign P[16] = in1[105] ^ in2[105];
    assign G[17] = in1[104] & in2[104];
    assign P[17] = in1[104] ^ in2[104];
    assign G[18] = in1[103] & in2[103];
    assign P[18] = in1[103] ^ in2[103];
    assign G[19] = in1[102] & in2[102];
    assign P[19] = in1[102] ^ in2[102];
    assign G[20] = in1[101] & in2[101];
    assign P[20] = in1[101] ^ in2[101];
    assign G[21] = in1[100] & in2[100];
    assign P[21] = in1[100] ^ in2[100];
    assign G[22] = in1[99] & in2[99];
    assign P[22] = in1[99] ^ in2[99];
    assign G[23] = in1[98] & in2[98];
    assign P[23] = in1[98] ^ in2[98];
    assign G[24] = in1[97] & in2[97];
    assign P[24] = in1[97] ^ in2[97];
    assign G[25] = in1[96] & in2[96];
    assign P[25] = in1[96] ^ in2[96];
    assign G[26] = in1[95] & in2[95];
    assign P[26] = in1[95] ^ in2[95];
    assign G[27] = in1[94] & in2[94];
    assign P[27] = in1[94] ^ in2[94];
    assign G[28] = in1[93] & in2[93];
    assign P[28] = in1[93] ^ in2[93];
    assign G[29] = in1[92] & in2[92];
    assign P[29] = in1[92] ^ in2[92];
    assign G[30] = in1[91] & in2[91];
    assign P[30] = in1[91] ^ in2[91];
    assign G[31] = in1[90] & in2[90];
    assign P[31] = in1[90] ^ in2[90];
    assign G[32] = in1[89] & in2[89];
    assign P[32] = in1[89] ^ in2[89];
    assign G[33] = in1[88] & in2[88];
    assign P[33] = in1[88] ^ in2[88];
    assign G[34] = in1[87] & in2[87];
    assign P[34] = in1[87] ^ in2[87];
    assign G[35] = in1[86] & in2[86];
    assign P[35] = in1[86] ^ in2[86];
    assign G[36] = in1[85] & in2[85];
    assign P[36] = in1[85] ^ in2[85];
    assign G[37] = in1[84] & in2[84];
    assign P[37] = in1[84] ^ in2[84];
    assign G[38] = in1[83] & in2[83];
    assign P[38] = in1[83] ^ in2[83];
    assign G[39] = in1[82] & in2[82];
    assign P[39] = in1[82] ^ in2[82];
    assign G[40] = in1[81] & in2[81];
    assign P[40] = in1[81] ^ in2[81];
    assign G[41] = in1[80] & in2[80];
    assign P[41] = in1[80] ^ in2[80];
    assign G[42] = in1[79] & in2[79];
    assign P[42] = in1[79] ^ in2[79];
    assign G[43] = in1[78] & in2[78];
    assign P[43] = in1[78] ^ in2[78];
    assign G[44] = in1[77] & in2[77];
    assign P[44] = in1[77] ^ in2[77];
    assign G[45] = in1[76] & in2[76];
    assign P[45] = in1[76] ^ in2[76];
    assign G[46] = in1[75] & in2[75];
    assign P[46] = in1[75] ^ in2[75];
    assign G[47] = in1[74] & in2[74];
    assign P[47] = in1[74] ^ in2[74];
    assign G[48] = in1[73] & in2[73];
    assign P[48] = in1[73] ^ in2[73];
    assign G[49] = in1[72] & in2[72];
    assign P[49] = in1[72] ^ in2[72];
    assign G[50] = in1[71] & in2[71];
    assign P[50] = in1[71] ^ in2[71];
    assign G[51] = in1[70] & in2[70];
    assign P[51] = in1[70] ^ in2[70];
    assign G[52] = in1[69] & in2[69];
    assign P[52] = in1[69] ^ in2[69];
    assign G[53] = in1[68] & in2[68];
    assign P[53] = in1[68] ^ in2[68];
    assign G[54] = in1[67] & in2[67];
    assign P[54] = in1[67] ^ in2[67];
    assign G[55] = in1[66] & in2[66];
    assign P[55] = in1[66] ^ in2[66];
    assign G[56] = in1[65] & in2[65];
    assign P[56] = in1[65] ^ in2[65];
    assign G[57] = in1[64] & in2[64];
    assign P[57] = in1[64] ^ in2[64];
    assign G[58] = in1[63] & in2[63];
    assign P[58] = in1[63] ^ in2[63];
    assign G[59] = in1[62] & in2[62];
    assign P[59] = in1[62] ^ in2[62];
    assign G[60] = in1[61] & in2[61];
    assign P[60] = in1[61] ^ in2[61];
    assign G[61] = in1[60] & in2[60];
    assign P[61] = in1[60] ^ in2[60];
    assign G[62] = in1[59] & in2[59];
    assign P[62] = in1[59] ^ in2[59];
    assign G[63] = in1[58] & in2[58];
    assign P[63] = in1[58] ^ in2[58];
    assign G[64] = in1[57] & in2[57];
    assign P[64] = in1[57] ^ in2[57];
    assign G[65] = in1[56] & in2[56];
    assign P[65] = in1[56] ^ in2[56];
    assign G[66] = in1[55] & in2[55];
    assign P[66] = in1[55] ^ in2[55];
    assign G[67] = in1[54] & in2[54];
    assign P[67] = in1[54] ^ in2[54];
    assign G[68] = in1[53] & in2[53];
    assign P[68] = in1[53] ^ in2[53];
    assign G[69] = in1[52] & in2[52];
    assign P[69] = in1[52] ^ in2[52];
    assign G[70] = in1[51] & in2[51];
    assign P[70] = in1[51] ^ in2[51];
    assign G[71] = in1[50] & in2[50];
    assign P[71] = in1[50] ^ in2[50];
    assign G[72] = in1[49] & in2[49];
    assign P[72] = in1[49] ^ in2[49];
    assign G[73] = in1[48] & in2[48];
    assign P[73] = in1[48] ^ in2[48];
    assign G[74] = in1[47] & in2[47];
    assign P[74] = in1[47] ^ in2[47];
    assign G[75] = in1[46] & in2[46];
    assign P[75] = in1[46] ^ in2[46];
    assign G[76] = in1[45] & in2[45];
    assign P[76] = in1[45] ^ in2[45];
    assign G[77] = in1[44] & in2[44];
    assign P[77] = in1[44] ^ in2[44];
    assign G[78] = in1[43] & in2[43];
    assign P[78] = in1[43] ^ in2[43];
    assign G[79] = in1[42] & in2[42];
    assign P[79] = in1[42] ^ in2[42];
    assign G[80] = in1[41] & in2[41];
    assign P[80] = in1[41] ^ in2[41];
    assign G[81] = in1[40] & in2[40];
    assign P[81] = in1[40] ^ in2[40];
    assign G[82] = in1[39] & in2[39];
    assign P[82] = in1[39] ^ in2[39];
    assign G[83] = in1[38] & in2[38];
    assign P[83] = in1[38] ^ in2[38];
    assign G[84] = in1[37] & in2[37];
    assign P[84] = in1[37] ^ in2[37];
    assign G[85] = in1[36] & in2[36];
    assign P[85] = in1[36] ^ in2[36];
    assign G[86] = in1[35] & in2[35];
    assign P[86] = in1[35] ^ in2[35];
    assign G[87] = in1[34] & in2[34];
    assign P[87] = in1[34] ^ in2[34];
    assign G[88] = in1[33] & in2[33];
    assign P[88] = in1[33] ^ in2[33];
    assign G[89] = in1[32] & in2[32];
    assign P[89] = in1[32] ^ in2[32];
    assign G[90] = in1[31] & in2[31];
    assign P[90] = in1[31] ^ in2[31];
    assign G[91] = in1[30] & in2[30];
    assign P[91] = in1[30] ^ in2[30];
    assign G[92] = in1[29] & in2[29];
    assign P[92] = in1[29] ^ in2[29];
    assign G[93] = in1[28] & in2[28];
    assign P[93] = in1[28] ^ in2[28];
    assign G[94] = in1[27] & in2[27];
    assign P[94] = in1[27] ^ in2[27];
    assign G[95] = in1[26] & in2[26];
    assign P[95] = in1[26] ^ in2[26];
    assign G[96] = in1[25] & in2[25];
    assign P[96] = in1[25] ^ in2[25];
    assign G[97] = in1[24] & in2[24];
    assign P[97] = in1[24] ^ in2[24];
    assign G[98] = in1[23] & in2[23];
    assign P[98] = in1[23] ^ in2[23];
    assign G[99] = in1[22] & in2[22];
    assign P[99] = in1[22] ^ in2[22];
    assign G[100] = in1[21] & in2[21];
    assign P[100] = in1[21] ^ in2[21];
    assign G[101] = in1[20] & in2[20];
    assign P[101] = in1[20] ^ in2[20];
    assign G[102] = in1[19] & in2[19];
    assign P[102] = in1[19] ^ in2[19];
    assign G[103] = in1[18] & in2[18];
    assign P[103] = in1[18] ^ in2[18];
    assign G[104] = in1[17] & in2[17];
    assign P[104] = in1[17] ^ in2[17];
    assign G[105] = in1[16] & in2[16];
    assign P[105] = in1[16] ^ in2[16];
    assign G[106] = in1[15] & in2[15];
    assign P[106] = in1[15] ^ in2[15];
    assign G[107] = in1[14] & in2[14];
    assign P[107] = in1[14] ^ in2[14];
    assign G[108] = in1[13] & in2[13];
    assign P[108] = in1[13] ^ in2[13];
    assign G[109] = in1[12] & in2[12];
    assign P[109] = in1[12] ^ in2[12];
    assign G[110] = in1[11] & in2[11];
    assign P[110] = in1[11] ^ in2[11];
    assign G[111] = in1[10] & in2[10];
    assign P[111] = in1[10] ^ in2[10];
    assign G[112] = in1[9] & in2[9];
    assign P[112] = in1[9] ^ in2[9];
    assign G[113] = in1[8] & in2[8];
    assign P[113] = in1[8] ^ in2[8];
    assign G[114] = in1[7] & in2[7];
    assign P[114] = in1[7] ^ in2[7];
    assign G[115] = in1[6] & in2[6];
    assign P[115] = in1[6] ^ in2[6];
    assign G[116] = in1[5] & in2[5];
    assign P[116] = in1[5] ^ in2[5];
    assign G[117] = in1[4] & in2[4];
    assign P[117] = in1[4] ^ in2[4];
    assign G[118] = in1[3] & in2[3];
    assign P[118] = in1[3] ^ in2[3];
    assign G[119] = in1[2] & in2[2];
    assign P[119] = in1[2] ^ in2[2];
    assign G[120] = in1[1] & in2[1];
    assign P[120] = in1[1] ^ in2[1];
    assign G[121] = in1[0] & in2[0];
    assign P[121] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign cout = G[121] | (P[121] & C[121]);
    assign sum = P ^ C;
endmodule

module CLA_121(output [120:0] sum, output cout, input [120:0] in1, input [120:0] in2);

    wire[120:0] G;
    wire[120:0] C;
    wire[120:0] P;

    assign G[0] = in1[120] & in2[120];
    assign P[0] = in1[120] ^ in2[120];
    assign G[1] = in1[119] & in2[119];
    assign P[1] = in1[119] ^ in2[119];
    assign G[2] = in1[118] & in2[118];
    assign P[2] = in1[118] ^ in2[118];
    assign G[3] = in1[117] & in2[117];
    assign P[3] = in1[117] ^ in2[117];
    assign G[4] = in1[116] & in2[116];
    assign P[4] = in1[116] ^ in2[116];
    assign G[5] = in1[115] & in2[115];
    assign P[5] = in1[115] ^ in2[115];
    assign G[6] = in1[114] & in2[114];
    assign P[6] = in1[114] ^ in2[114];
    assign G[7] = in1[113] & in2[113];
    assign P[7] = in1[113] ^ in2[113];
    assign G[8] = in1[112] & in2[112];
    assign P[8] = in1[112] ^ in2[112];
    assign G[9] = in1[111] & in2[111];
    assign P[9] = in1[111] ^ in2[111];
    assign G[10] = in1[110] & in2[110];
    assign P[10] = in1[110] ^ in2[110];
    assign G[11] = in1[109] & in2[109];
    assign P[11] = in1[109] ^ in2[109];
    assign G[12] = in1[108] & in2[108];
    assign P[12] = in1[108] ^ in2[108];
    assign G[13] = in1[107] & in2[107];
    assign P[13] = in1[107] ^ in2[107];
    assign G[14] = in1[106] & in2[106];
    assign P[14] = in1[106] ^ in2[106];
    assign G[15] = in1[105] & in2[105];
    assign P[15] = in1[105] ^ in2[105];
    assign G[16] = in1[104] & in2[104];
    assign P[16] = in1[104] ^ in2[104];
    assign G[17] = in1[103] & in2[103];
    assign P[17] = in1[103] ^ in2[103];
    assign G[18] = in1[102] & in2[102];
    assign P[18] = in1[102] ^ in2[102];
    assign G[19] = in1[101] & in2[101];
    assign P[19] = in1[101] ^ in2[101];
    assign G[20] = in1[100] & in2[100];
    assign P[20] = in1[100] ^ in2[100];
    assign G[21] = in1[99] & in2[99];
    assign P[21] = in1[99] ^ in2[99];
    assign G[22] = in1[98] & in2[98];
    assign P[22] = in1[98] ^ in2[98];
    assign G[23] = in1[97] & in2[97];
    assign P[23] = in1[97] ^ in2[97];
    assign G[24] = in1[96] & in2[96];
    assign P[24] = in1[96] ^ in2[96];
    assign G[25] = in1[95] & in2[95];
    assign P[25] = in1[95] ^ in2[95];
    assign G[26] = in1[94] & in2[94];
    assign P[26] = in1[94] ^ in2[94];
    assign G[27] = in1[93] & in2[93];
    assign P[27] = in1[93] ^ in2[93];
    assign G[28] = in1[92] & in2[92];
    assign P[28] = in1[92] ^ in2[92];
    assign G[29] = in1[91] & in2[91];
    assign P[29] = in1[91] ^ in2[91];
    assign G[30] = in1[90] & in2[90];
    assign P[30] = in1[90] ^ in2[90];
    assign G[31] = in1[89] & in2[89];
    assign P[31] = in1[89] ^ in2[89];
    assign G[32] = in1[88] & in2[88];
    assign P[32] = in1[88] ^ in2[88];
    assign G[33] = in1[87] & in2[87];
    assign P[33] = in1[87] ^ in2[87];
    assign G[34] = in1[86] & in2[86];
    assign P[34] = in1[86] ^ in2[86];
    assign G[35] = in1[85] & in2[85];
    assign P[35] = in1[85] ^ in2[85];
    assign G[36] = in1[84] & in2[84];
    assign P[36] = in1[84] ^ in2[84];
    assign G[37] = in1[83] & in2[83];
    assign P[37] = in1[83] ^ in2[83];
    assign G[38] = in1[82] & in2[82];
    assign P[38] = in1[82] ^ in2[82];
    assign G[39] = in1[81] & in2[81];
    assign P[39] = in1[81] ^ in2[81];
    assign G[40] = in1[80] & in2[80];
    assign P[40] = in1[80] ^ in2[80];
    assign G[41] = in1[79] & in2[79];
    assign P[41] = in1[79] ^ in2[79];
    assign G[42] = in1[78] & in2[78];
    assign P[42] = in1[78] ^ in2[78];
    assign G[43] = in1[77] & in2[77];
    assign P[43] = in1[77] ^ in2[77];
    assign G[44] = in1[76] & in2[76];
    assign P[44] = in1[76] ^ in2[76];
    assign G[45] = in1[75] & in2[75];
    assign P[45] = in1[75] ^ in2[75];
    assign G[46] = in1[74] & in2[74];
    assign P[46] = in1[74] ^ in2[74];
    assign G[47] = in1[73] & in2[73];
    assign P[47] = in1[73] ^ in2[73];
    assign G[48] = in1[72] & in2[72];
    assign P[48] = in1[72] ^ in2[72];
    assign G[49] = in1[71] & in2[71];
    assign P[49] = in1[71] ^ in2[71];
    assign G[50] = in1[70] & in2[70];
    assign P[50] = in1[70] ^ in2[70];
    assign G[51] = in1[69] & in2[69];
    assign P[51] = in1[69] ^ in2[69];
    assign G[52] = in1[68] & in2[68];
    assign P[52] = in1[68] ^ in2[68];
    assign G[53] = in1[67] & in2[67];
    assign P[53] = in1[67] ^ in2[67];
    assign G[54] = in1[66] & in2[66];
    assign P[54] = in1[66] ^ in2[66];
    assign G[55] = in1[65] & in2[65];
    assign P[55] = in1[65] ^ in2[65];
    assign G[56] = in1[64] & in2[64];
    assign P[56] = in1[64] ^ in2[64];
    assign G[57] = in1[63] & in2[63];
    assign P[57] = in1[63] ^ in2[63];
    assign G[58] = in1[62] & in2[62];
    assign P[58] = in1[62] ^ in2[62];
    assign G[59] = in1[61] & in2[61];
    assign P[59] = in1[61] ^ in2[61];
    assign G[60] = in1[60] & in2[60];
    assign P[60] = in1[60] ^ in2[60];
    assign G[61] = in1[59] & in2[59];
    assign P[61] = in1[59] ^ in2[59];
    assign G[62] = in1[58] & in2[58];
    assign P[62] = in1[58] ^ in2[58];
    assign G[63] = in1[57] & in2[57];
    assign P[63] = in1[57] ^ in2[57];
    assign G[64] = in1[56] & in2[56];
    assign P[64] = in1[56] ^ in2[56];
    assign G[65] = in1[55] & in2[55];
    assign P[65] = in1[55] ^ in2[55];
    assign G[66] = in1[54] & in2[54];
    assign P[66] = in1[54] ^ in2[54];
    assign G[67] = in1[53] & in2[53];
    assign P[67] = in1[53] ^ in2[53];
    assign G[68] = in1[52] & in2[52];
    assign P[68] = in1[52] ^ in2[52];
    assign G[69] = in1[51] & in2[51];
    assign P[69] = in1[51] ^ in2[51];
    assign G[70] = in1[50] & in2[50];
    assign P[70] = in1[50] ^ in2[50];
    assign G[71] = in1[49] & in2[49];
    assign P[71] = in1[49] ^ in2[49];
    assign G[72] = in1[48] & in2[48];
    assign P[72] = in1[48] ^ in2[48];
    assign G[73] = in1[47] & in2[47];
    assign P[73] = in1[47] ^ in2[47];
    assign G[74] = in1[46] & in2[46];
    assign P[74] = in1[46] ^ in2[46];
    assign G[75] = in1[45] & in2[45];
    assign P[75] = in1[45] ^ in2[45];
    assign G[76] = in1[44] & in2[44];
    assign P[76] = in1[44] ^ in2[44];
    assign G[77] = in1[43] & in2[43];
    assign P[77] = in1[43] ^ in2[43];
    assign G[78] = in1[42] & in2[42];
    assign P[78] = in1[42] ^ in2[42];
    assign G[79] = in1[41] & in2[41];
    assign P[79] = in1[41] ^ in2[41];
    assign G[80] = in1[40] & in2[40];
    assign P[80] = in1[40] ^ in2[40];
    assign G[81] = in1[39] & in2[39];
    assign P[81] = in1[39] ^ in2[39];
    assign G[82] = in1[38] & in2[38];
    assign P[82] = in1[38] ^ in2[38];
    assign G[83] = in1[37] & in2[37];
    assign P[83] = in1[37] ^ in2[37];
    assign G[84] = in1[36] & in2[36];
    assign P[84] = in1[36] ^ in2[36];
    assign G[85] = in1[35] & in2[35];
    assign P[85] = in1[35] ^ in2[35];
    assign G[86] = in1[34] & in2[34];
    assign P[86] = in1[34] ^ in2[34];
    assign G[87] = in1[33] & in2[33];
    assign P[87] = in1[33] ^ in2[33];
    assign G[88] = in1[32] & in2[32];
    assign P[88] = in1[32] ^ in2[32];
    assign G[89] = in1[31] & in2[31];
    assign P[89] = in1[31] ^ in2[31];
    assign G[90] = in1[30] & in2[30];
    assign P[90] = in1[30] ^ in2[30];
    assign G[91] = in1[29] & in2[29];
    assign P[91] = in1[29] ^ in2[29];
    assign G[92] = in1[28] & in2[28];
    assign P[92] = in1[28] ^ in2[28];
    assign G[93] = in1[27] & in2[27];
    assign P[93] = in1[27] ^ in2[27];
    assign G[94] = in1[26] & in2[26];
    assign P[94] = in1[26] ^ in2[26];
    assign G[95] = in1[25] & in2[25];
    assign P[95] = in1[25] ^ in2[25];
    assign G[96] = in1[24] & in2[24];
    assign P[96] = in1[24] ^ in2[24];
    assign G[97] = in1[23] & in2[23];
    assign P[97] = in1[23] ^ in2[23];
    assign G[98] = in1[22] & in2[22];
    assign P[98] = in1[22] ^ in2[22];
    assign G[99] = in1[21] & in2[21];
    assign P[99] = in1[21] ^ in2[21];
    assign G[100] = in1[20] & in2[20];
    assign P[100] = in1[20] ^ in2[20];
    assign G[101] = in1[19] & in2[19];
    assign P[101] = in1[19] ^ in2[19];
    assign G[102] = in1[18] & in2[18];
    assign P[102] = in1[18] ^ in2[18];
    assign G[103] = in1[17] & in2[17];
    assign P[103] = in1[17] ^ in2[17];
    assign G[104] = in1[16] & in2[16];
    assign P[104] = in1[16] ^ in2[16];
    assign G[105] = in1[15] & in2[15];
    assign P[105] = in1[15] ^ in2[15];
    assign G[106] = in1[14] & in2[14];
    assign P[106] = in1[14] ^ in2[14];
    assign G[107] = in1[13] & in2[13];
    assign P[107] = in1[13] ^ in2[13];
    assign G[108] = in1[12] & in2[12];
    assign P[108] = in1[12] ^ in2[12];
    assign G[109] = in1[11] & in2[11];
    assign P[109] = in1[11] ^ in2[11];
    assign G[110] = in1[10] & in2[10];
    assign P[110] = in1[10] ^ in2[10];
    assign G[111] = in1[9] & in2[9];
    assign P[111] = in1[9] ^ in2[9];
    assign G[112] = in1[8] & in2[8];
    assign P[112] = in1[8] ^ in2[8];
    assign G[113] = in1[7] & in2[7];
    assign P[113] = in1[7] ^ in2[7];
    assign G[114] = in1[6] & in2[6];
    assign P[114] = in1[6] ^ in2[6];
    assign G[115] = in1[5] & in2[5];
    assign P[115] = in1[5] ^ in2[5];
    assign G[116] = in1[4] & in2[4];
    assign P[116] = in1[4] ^ in2[4];
    assign G[117] = in1[3] & in2[3];
    assign P[117] = in1[3] ^ in2[3];
    assign G[118] = in1[2] & in2[2];
    assign P[118] = in1[2] ^ in2[2];
    assign G[119] = in1[1] & in2[1];
    assign P[119] = in1[1] ^ in2[1];
    assign G[120] = in1[0] & in2[0];
    assign P[120] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign cout = G[120] | (P[120] & C[120]);
    assign sum = P ^ C;
endmodule

module CLA_120(output [119:0] sum, output cout, input [119:0] in1, input [119:0] in2);

    wire[119:0] G;
    wire[119:0] C;
    wire[119:0] P;

    assign G[0] = in1[119] & in2[119];
    assign P[0] = in1[119] ^ in2[119];
    assign G[1] = in1[118] & in2[118];
    assign P[1] = in1[118] ^ in2[118];
    assign G[2] = in1[117] & in2[117];
    assign P[2] = in1[117] ^ in2[117];
    assign G[3] = in1[116] & in2[116];
    assign P[3] = in1[116] ^ in2[116];
    assign G[4] = in1[115] & in2[115];
    assign P[4] = in1[115] ^ in2[115];
    assign G[5] = in1[114] & in2[114];
    assign P[5] = in1[114] ^ in2[114];
    assign G[6] = in1[113] & in2[113];
    assign P[6] = in1[113] ^ in2[113];
    assign G[7] = in1[112] & in2[112];
    assign P[7] = in1[112] ^ in2[112];
    assign G[8] = in1[111] & in2[111];
    assign P[8] = in1[111] ^ in2[111];
    assign G[9] = in1[110] & in2[110];
    assign P[9] = in1[110] ^ in2[110];
    assign G[10] = in1[109] & in2[109];
    assign P[10] = in1[109] ^ in2[109];
    assign G[11] = in1[108] & in2[108];
    assign P[11] = in1[108] ^ in2[108];
    assign G[12] = in1[107] & in2[107];
    assign P[12] = in1[107] ^ in2[107];
    assign G[13] = in1[106] & in2[106];
    assign P[13] = in1[106] ^ in2[106];
    assign G[14] = in1[105] & in2[105];
    assign P[14] = in1[105] ^ in2[105];
    assign G[15] = in1[104] & in2[104];
    assign P[15] = in1[104] ^ in2[104];
    assign G[16] = in1[103] & in2[103];
    assign P[16] = in1[103] ^ in2[103];
    assign G[17] = in1[102] & in2[102];
    assign P[17] = in1[102] ^ in2[102];
    assign G[18] = in1[101] & in2[101];
    assign P[18] = in1[101] ^ in2[101];
    assign G[19] = in1[100] & in2[100];
    assign P[19] = in1[100] ^ in2[100];
    assign G[20] = in1[99] & in2[99];
    assign P[20] = in1[99] ^ in2[99];
    assign G[21] = in1[98] & in2[98];
    assign P[21] = in1[98] ^ in2[98];
    assign G[22] = in1[97] & in2[97];
    assign P[22] = in1[97] ^ in2[97];
    assign G[23] = in1[96] & in2[96];
    assign P[23] = in1[96] ^ in2[96];
    assign G[24] = in1[95] & in2[95];
    assign P[24] = in1[95] ^ in2[95];
    assign G[25] = in1[94] & in2[94];
    assign P[25] = in1[94] ^ in2[94];
    assign G[26] = in1[93] & in2[93];
    assign P[26] = in1[93] ^ in2[93];
    assign G[27] = in1[92] & in2[92];
    assign P[27] = in1[92] ^ in2[92];
    assign G[28] = in1[91] & in2[91];
    assign P[28] = in1[91] ^ in2[91];
    assign G[29] = in1[90] & in2[90];
    assign P[29] = in1[90] ^ in2[90];
    assign G[30] = in1[89] & in2[89];
    assign P[30] = in1[89] ^ in2[89];
    assign G[31] = in1[88] & in2[88];
    assign P[31] = in1[88] ^ in2[88];
    assign G[32] = in1[87] & in2[87];
    assign P[32] = in1[87] ^ in2[87];
    assign G[33] = in1[86] & in2[86];
    assign P[33] = in1[86] ^ in2[86];
    assign G[34] = in1[85] & in2[85];
    assign P[34] = in1[85] ^ in2[85];
    assign G[35] = in1[84] & in2[84];
    assign P[35] = in1[84] ^ in2[84];
    assign G[36] = in1[83] & in2[83];
    assign P[36] = in1[83] ^ in2[83];
    assign G[37] = in1[82] & in2[82];
    assign P[37] = in1[82] ^ in2[82];
    assign G[38] = in1[81] & in2[81];
    assign P[38] = in1[81] ^ in2[81];
    assign G[39] = in1[80] & in2[80];
    assign P[39] = in1[80] ^ in2[80];
    assign G[40] = in1[79] & in2[79];
    assign P[40] = in1[79] ^ in2[79];
    assign G[41] = in1[78] & in2[78];
    assign P[41] = in1[78] ^ in2[78];
    assign G[42] = in1[77] & in2[77];
    assign P[42] = in1[77] ^ in2[77];
    assign G[43] = in1[76] & in2[76];
    assign P[43] = in1[76] ^ in2[76];
    assign G[44] = in1[75] & in2[75];
    assign P[44] = in1[75] ^ in2[75];
    assign G[45] = in1[74] & in2[74];
    assign P[45] = in1[74] ^ in2[74];
    assign G[46] = in1[73] & in2[73];
    assign P[46] = in1[73] ^ in2[73];
    assign G[47] = in1[72] & in2[72];
    assign P[47] = in1[72] ^ in2[72];
    assign G[48] = in1[71] & in2[71];
    assign P[48] = in1[71] ^ in2[71];
    assign G[49] = in1[70] & in2[70];
    assign P[49] = in1[70] ^ in2[70];
    assign G[50] = in1[69] & in2[69];
    assign P[50] = in1[69] ^ in2[69];
    assign G[51] = in1[68] & in2[68];
    assign P[51] = in1[68] ^ in2[68];
    assign G[52] = in1[67] & in2[67];
    assign P[52] = in1[67] ^ in2[67];
    assign G[53] = in1[66] & in2[66];
    assign P[53] = in1[66] ^ in2[66];
    assign G[54] = in1[65] & in2[65];
    assign P[54] = in1[65] ^ in2[65];
    assign G[55] = in1[64] & in2[64];
    assign P[55] = in1[64] ^ in2[64];
    assign G[56] = in1[63] & in2[63];
    assign P[56] = in1[63] ^ in2[63];
    assign G[57] = in1[62] & in2[62];
    assign P[57] = in1[62] ^ in2[62];
    assign G[58] = in1[61] & in2[61];
    assign P[58] = in1[61] ^ in2[61];
    assign G[59] = in1[60] & in2[60];
    assign P[59] = in1[60] ^ in2[60];
    assign G[60] = in1[59] & in2[59];
    assign P[60] = in1[59] ^ in2[59];
    assign G[61] = in1[58] & in2[58];
    assign P[61] = in1[58] ^ in2[58];
    assign G[62] = in1[57] & in2[57];
    assign P[62] = in1[57] ^ in2[57];
    assign G[63] = in1[56] & in2[56];
    assign P[63] = in1[56] ^ in2[56];
    assign G[64] = in1[55] & in2[55];
    assign P[64] = in1[55] ^ in2[55];
    assign G[65] = in1[54] & in2[54];
    assign P[65] = in1[54] ^ in2[54];
    assign G[66] = in1[53] & in2[53];
    assign P[66] = in1[53] ^ in2[53];
    assign G[67] = in1[52] & in2[52];
    assign P[67] = in1[52] ^ in2[52];
    assign G[68] = in1[51] & in2[51];
    assign P[68] = in1[51] ^ in2[51];
    assign G[69] = in1[50] & in2[50];
    assign P[69] = in1[50] ^ in2[50];
    assign G[70] = in1[49] & in2[49];
    assign P[70] = in1[49] ^ in2[49];
    assign G[71] = in1[48] & in2[48];
    assign P[71] = in1[48] ^ in2[48];
    assign G[72] = in1[47] & in2[47];
    assign P[72] = in1[47] ^ in2[47];
    assign G[73] = in1[46] & in2[46];
    assign P[73] = in1[46] ^ in2[46];
    assign G[74] = in1[45] & in2[45];
    assign P[74] = in1[45] ^ in2[45];
    assign G[75] = in1[44] & in2[44];
    assign P[75] = in1[44] ^ in2[44];
    assign G[76] = in1[43] & in2[43];
    assign P[76] = in1[43] ^ in2[43];
    assign G[77] = in1[42] & in2[42];
    assign P[77] = in1[42] ^ in2[42];
    assign G[78] = in1[41] & in2[41];
    assign P[78] = in1[41] ^ in2[41];
    assign G[79] = in1[40] & in2[40];
    assign P[79] = in1[40] ^ in2[40];
    assign G[80] = in1[39] & in2[39];
    assign P[80] = in1[39] ^ in2[39];
    assign G[81] = in1[38] & in2[38];
    assign P[81] = in1[38] ^ in2[38];
    assign G[82] = in1[37] & in2[37];
    assign P[82] = in1[37] ^ in2[37];
    assign G[83] = in1[36] & in2[36];
    assign P[83] = in1[36] ^ in2[36];
    assign G[84] = in1[35] & in2[35];
    assign P[84] = in1[35] ^ in2[35];
    assign G[85] = in1[34] & in2[34];
    assign P[85] = in1[34] ^ in2[34];
    assign G[86] = in1[33] & in2[33];
    assign P[86] = in1[33] ^ in2[33];
    assign G[87] = in1[32] & in2[32];
    assign P[87] = in1[32] ^ in2[32];
    assign G[88] = in1[31] & in2[31];
    assign P[88] = in1[31] ^ in2[31];
    assign G[89] = in1[30] & in2[30];
    assign P[89] = in1[30] ^ in2[30];
    assign G[90] = in1[29] & in2[29];
    assign P[90] = in1[29] ^ in2[29];
    assign G[91] = in1[28] & in2[28];
    assign P[91] = in1[28] ^ in2[28];
    assign G[92] = in1[27] & in2[27];
    assign P[92] = in1[27] ^ in2[27];
    assign G[93] = in1[26] & in2[26];
    assign P[93] = in1[26] ^ in2[26];
    assign G[94] = in1[25] & in2[25];
    assign P[94] = in1[25] ^ in2[25];
    assign G[95] = in1[24] & in2[24];
    assign P[95] = in1[24] ^ in2[24];
    assign G[96] = in1[23] & in2[23];
    assign P[96] = in1[23] ^ in2[23];
    assign G[97] = in1[22] & in2[22];
    assign P[97] = in1[22] ^ in2[22];
    assign G[98] = in1[21] & in2[21];
    assign P[98] = in1[21] ^ in2[21];
    assign G[99] = in1[20] & in2[20];
    assign P[99] = in1[20] ^ in2[20];
    assign G[100] = in1[19] & in2[19];
    assign P[100] = in1[19] ^ in2[19];
    assign G[101] = in1[18] & in2[18];
    assign P[101] = in1[18] ^ in2[18];
    assign G[102] = in1[17] & in2[17];
    assign P[102] = in1[17] ^ in2[17];
    assign G[103] = in1[16] & in2[16];
    assign P[103] = in1[16] ^ in2[16];
    assign G[104] = in1[15] & in2[15];
    assign P[104] = in1[15] ^ in2[15];
    assign G[105] = in1[14] & in2[14];
    assign P[105] = in1[14] ^ in2[14];
    assign G[106] = in1[13] & in2[13];
    assign P[106] = in1[13] ^ in2[13];
    assign G[107] = in1[12] & in2[12];
    assign P[107] = in1[12] ^ in2[12];
    assign G[108] = in1[11] & in2[11];
    assign P[108] = in1[11] ^ in2[11];
    assign G[109] = in1[10] & in2[10];
    assign P[109] = in1[10] ^ in2[10];
    assign G[110] = in1[9] & in2[9];
    assign P[110] = in1[9] ^ in2[9];
    assign G[111] = in1[8] & in2[8];
    assign P[111] = in1[8] ^ in2[8];
    assign G[112] = in1[7] & in2[7];
    assign P[112] = in1[7] ^ in2[7];
    assign G[113] = in1[6] & in2[6];
    assign P[113] = in1[6] ^ in2[6];
    assign G[114] = in1[5] & in2[5];
    assign P[114] = in1[5] ^ in2[5];
    assign G[115] = in1[4] & in2[4];
    assign P[115] = in1[4] ^ in2[4];
    assign G[116] = in1[3] & in2[3];
    assign P[116] = in1[3] ^ in2[3];
    assign G[117] = in1[2] & in2[2];
    assign P[117] = in1[2] ^ in2[2];
    assign G[118] = in1[1] & in2[1];
    assign P[118] = in1[1] ^ in2[1];
    assign G[119] = in1[0] & in2[0];
    assign P[119] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign cout = G[119] | (P[119] & C[119]);
    assign sum = P ^ C;
endmodule

module CLA_119(output [118:0] sum, output cout, input [118:0] in1, input [118:0] in2);

    wire[118:0] G;
    wire[118:0] C;
    wire[118:0] P;

    assign G[0] = in1[118] & in2[118];
    assign P[0] = in1[118] ^ in2[118];
    assign G[1] = in1[117] & in2[117];
    assign P[1] = in1[117] ^ in2[117];
    assign G[2] = in1[116] & in2[116];
    assign P[2] = in1[116] ^ in2[116];
    assign G[3] = in1[115] & in2[115];
    assign P[3] = in1[115] ^ in2[115];
    assign G[4] = in1[114] & in2[114];
    assign P[4] = in1[114] ^ in2[114];
    assign G[5] = in1[113] & in2[113];
    assign P[5] = in1[113] ^ in2[113];
    assign G[6] = in1[112] & in2[112];
    assign P[6] = in1[112] ^ in2[112];
    assign G[7] = in1[111] & in2[111];
    assign P[7] = in1[111] ^ in2[111];
    assign G[8] = in1[110] & in2[110];
    assign P[8] = in1[110] ^ in2[110];
    assign G[9] = in1[109] & in2[109];
    assign P[9] = in1[109] ^ in2[109];
    assign G[10] = in1[108] & in2[108];
    assign P[10] = in1[108] ^ in2[108];
    assign G[11] = in1[107] & in2[107];
    assign P[11] = in1[107] ^ in2[107];
    assign G[12] = in1[106] & in2[106];
    assign P[12] = in1[106] ^ in2[106];
    assign G[13] = in1[105] & in2[105];
    assign P[13] = in1[105] ^ in2[105];
    assign G[14] = in1[104] & in2[104];
    assign P[14] = in1[104] ^ in2[104];
    assign G[15] = in1[103] & in2[103];
    assign P[15] = in1[103] ^ in2[103];
    assign G[16] = in1[102] & in2[102];
    assign P[16] = in1[102] ^ in2[102];
    assign G[17] = in1[101] & in2[101];
    assign P[17] = in1[101] ^ in2[101];
    assign G[18] = in1[100] & in2[100];
    assign P[18] = in1[100] ^ in2[100];
    assign G[19] = in1[99] & in2[99];
    assign P[19] = in1[99] ^ in2[99];
    assign G[20] = in1[98] & in2[98];
    assign P[20] = in1[98] ^ in2[98];
    assign G[21] = in1[97] & in2[97];
    assign P[21] = in1[97] ^ in2[97];
    assign G[22] = in1[96] & in2[96];
    assign P[22] = in1[96] ^ in2[96];
    assign G[23] = in1[95] & in2[95];
    assign P[23] = in1[95] ^ in2[95];
    assign G[24] = in1[94] & in2[94];
    assign P[24] = in1[94] ^ in2[94];
    assign G[25] = in1[93] & in2[93];
    assign P[25] = in1[93] ^ in2[93];
    assign G[26] = in1[92] & in2[92];
    assign P[26] = in1[92] ^ in2[92];
    assign G[27] = in1[91] & in2[91];
    assign P[27] = in1[91] ^ in2[91];
    assign G[28] = in1[90] & in2[90];
    assign P[28] = in1[90] ^ in2[90];
    assign G[29] = in1[89] & in2[89];
    assign P[29] = in1[89] ^ in2[89];
    assign G[30] = in1[88] & in2[88];
    assign P[30] = in1[88] ^ in2[88];
    assign G[31] = in1[87] & in2[87];
    assign P[31] = in1[87] ^ in2[87];
    assign G[32] = in1[86] & in2[86];
    assign P[32] = in1[86] ^ in2[86];
    assign G[33] = in1[85] & in2[85];
    assign P[33] = in1[85] ^ in2[85];
    assign G[34] = in1[84] & in2[84];
    assign P[34] = in1[84] ^ in2[84];
    assign G[35] = in1[83] & in2[83];
    assign P[35] = in1[83] ^ in2[83];
    assign G[36] = in1[82] & in2[82];
    assign P[36] = in1[82] ^ in2[82];
    assign G[37] = in1[81] & in2[81];
    assign P[37] = in1[81] ^ in2[81];
    assign G[38] = in1[80] & in2[80];
    assign P[38] = in1[80] ^ in2[80];
    assign G[39] = in1[79] & in2[79];
    assign P[39] = in1[79] ^ in2[79];
    assign G[40] = in1[78] & in2[78];
    assign P[40] = in1[78] ^ in2[78];
    assign G[41] = in1[77] & in2[77];
    assign P[41] = in1[77] ^ in2[77];
    assign G[42] = in1[76] & in2[76];
    assign P[42] = in1[76] ^ in2[76];
    assign G[43] = in1[75] & in2[75];
    assign P[43] = in1[75] ^ in2[75];
    assign G[44] = in1[74] & in2[74];
    assign P[44] = in1[74] ^ in2[74];
    assign G[45] = in1[73] & in2[73];
    assign P[45] = in1[73] ^ in2[73];
    assign G[46] = in1[72] & in2[72];
    assign P[46] = in1[72] ^ in2[72];
    assign G[47] = in1[71] & in2[71];
    assign P[47] = in1[71] ^ in2[71];
    assign G[48] = in1[70] & in2[70];
    assign P[48] = in1[70] ^ in2[70];
    assign G[49] = in1[69] & in2[69];
    assign P[49] = in1[69] ^ in2[69];
    assign G[50] = in1[68] & in2[68];
    assign P[50] = in1[68] ^ in2[68];
    assign G[51] = in1[67] & in2[67];
    assign P[51] = in1[67] ^ in2[67];
    assign G[52] = in1[66] & in2[66];
    assign P[52] = in1[66] ^ in2[66];
    assign G[53] = in1[65] & in2[65];
    assign P[53] = in1[65] ^ in2[65];
    assign G[54] = in1[64] & in2[64];
    assign P[54] = in1[64] ^ in2[64];
    assign G[55] = in1[63] & in2[63];
    assign P[55] = in1[63] ^ in2[63];
    assign G[56] = in1[62] & in2[62];
    assign P[56] = in1[62] ^ in2[62];
    assign G[57] = in1[61] & in2[61];
    assign P[57] = in1[61] ^ in2[61];
    assign G[58] = in1[60] & in2[60];
    assign P[58] = in1[60] ^ in2[60];
    assign G[59] = in1[59] & in2[59];
    assign P[59] = in1[59] ^ in2[59];
    assign G[60] = in1[58] & in2[58];
    assign P[60] = in1[58] ^ in2[58];
    assign G[61] = in1[57] & in2[57];
    assign P[61] = in1[57] ^ in2[57];
    assign G[62] = in1[56] & in2[56];
    assign P[62] = in1[56] ^ in2[56];
    assign G[63] = in1[55] & in2[55];
    assign P[63] = in1[55] ^ in2[55];
    assign G[64] = in1[54] & in2[54];
    assign P[64] = in1[54] ^ in2[54];
    assign G[65] = in1[53] & in2[53];
    assign P[65] = in1[53] ^ in2[53];
    assign G[66] = in1[52] & in2[52];
    assign P[66] = in1[52] ^ in2[52];
    assign G[67] = in1[51] & in2[51];
    assign P[67] = in1[51] ^ in2[51];
    assign G[68] = in1[50] & in2[50];
    assign P[68] = in1[50] ^ in2[50];
    assign G[69] = in1[49] & in2[49];
    assign P[69] = in1[49] ^ in2[49];
    assign G[70] = in1[48] & in2[48];
    assign P[70] = in1[48] ^ in2[48];
    assign G[71] = in1[47] & in2[47];
    assign P[71] = in1[47] ^ in2[47];
    assign G[72] = in1[46] & in2[46];
    assign P[72] = in1[46] ^ in2[46];
    assign G[73] = in1[45] & in2[45];
    assign P[73] = in1[45] ^ in2[45];
    assign G[74] = in1[44] & in2[44];
    assign P[74] = in1[44] ^ in2[44];
    assign G[75] = in1[43] & in2[43];
    assign P[75] = in1[43] ^ in2[43];
    assign G[76] = in1[42] & in2[42];
    assign P[76] = in1[42] ^ in2[42];
    assign G[77] = in1[41] & in2[41];
    assign P[77] = in1[41] ^ in2[41];
    assign G[78] = in1[40] & in2[40];
    assign P[78] = in1[40] ^ in2[40];
    assign G[79] = in1[39] & in2[39];
    assign P[79] = in1[39] ^ in2[39];
    assign G[80] = in1[38] & in2[38];
    assign P[80] = in1[38] ^ in2[38];
    assign G[81] = in1[37] & in2[37];
    assign P[81] = in1[37] ^ in2[37];
    assign G[82] = in1[36] & in2[36];
    assign P[82] = in1[36] ^ in2[36];
    assign G[83] = in1[35] & in2[35];
    assign P[83] = in1[35] ^ in2[35];
    assign G[84] = in1[34] & in2[34];
    assign P[84] = in1[34] ^ in2[34];
    assign G[85] = in1[33] & in2[33];
    assign P[85] = in1[33] ^ in2[33];
    assign G[86] = in1[32] & in2[32];
    assign P[86] = in1[32] ^ in2[32];
    assign G[87] = in1[31] & in2[31];
    assign P[87] = in1[31] ^ in2[31];
    assign G[88] = in1[30] & in2[30];
    assign P[88] = in1[30] ^ in2[30];
    assign G[89] = in1[29] & in2[29];
    assign P[89] = in1[29] ^ in2[29];
    assign G[90] = in1[28] & in2[28];
    assign P[90] = in1[28] ^ in2[28];
    assign G[91] = in1[27] & in2[27];
    assign P[91] = in1[27] ^ in2[27];
    assign G[92] = in1[26] & in2[26];
    assign P[92] = in1[26] ^ in2[26];
    assign G[93] = in1[25] & in2[25];
    assign P[93] = in1[25] ^ in2[25];
    assign G[94] = in1[24] & in2[24];
    assign P[94] = in1[24] ^ in2[24];
    assign G[95] = in1[23] & in2[23];
    assign P[95] = in1[23] ^ in2[23];
    assign G[96] = in1[22] & in2[22];
    assign P[96] = in1[22] ^ in2[22];
    assign G[97] = in1[21] & in2[21];
    assign P[97] = in1[21] ^ in2[21];
    assign G[98] = in1[20] & in2[20];
    assign P[98] = in1[20] ^ in2[20];
    assign G[99] = in1[19] & in2[19];
    assign P[99] = in1[19] ^ in2[19];
    assign G[100] = in1[18] & in2[18];
    assign P[100] = in1[18] ^ in2[18];
    assign G[101] = in1[17] & in2[17];
    assign P[101] = in1[17] ^ in2[17];
    assign G[102] = in1[16] & in2[16];
    assign P[102] = in1[16] ^ in2[16];
    assign G[103] = in1[15] & in2[15];
    assign P[103] = in1[15] ^ in2[15];
    assign G[104] = in1[14] & in2[14];
    assign P[104] = in1[14] ^ in2[14];
    assign G[105] = in1[13] & in2[13];
    assign P[105] = in1[13] ^ in2[13];
    assign G[106] = in1[12] & in2[12];
    assign P[106] = in1[12] ^ in2[12];
    assign G[107] = in1[11] & in2[11];
    assign P[107] = in1[11] ^ in2[11];
    assign G[108] = in1[10] & in2[10];
    assign P[108] = in1[10] ^ in2[10];
    assign G[109] = in1[9] & in2[9];
    assign P[109] = in1[9] ^ in2[9];
    assign G[110] = in1[8] & in2[8];
    assign P[110] = in1[8] ^ in2[8];
    assign G[111] = in1[7] & in2[7];
    assign P[111] = in1[7] ^ in2[7];
    assign G[112] = in1[6] & in2[6];
    assign P[112] = in1[6] ^ in2[6];
    assign G[113] = in1[5] & in2[5];
    assign P[113] = in1[5] ^ in2[5];
    assign G[114] = in1[4] & in2[4];
    assign P[114] = in1[4] ^ in2[4];
    assign G[115] = in1[3] & in2[3];
    assign P[115] = in1[3] ^ in2[3];
    assign G[116] = in1[2] & in2[2];
    assign P[116] = in1[2] ^ in2[2];
    assign G[117] = in1[1] & in2[1];
    assign P[117] = in1[1] ^ in2[1];
    assign G[118] = in1[0] & in2[0];
    assign P[118] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign cout = G[118] | (P[118] & C[118]);
    assign sum = P ^ C;
endmodule

module CLA_118(output [117:0] sum, output cout, input [117:0] in1, input [117:0] in2);

    wire[117:0] G;
    wire[117:0] C;
    wire[117:0] P;

    assign G[0] = in1[117] & in2[117];
    assign P[0] = in1[117] ^ in2[117];
    assign G[1] = in1[116] & in2[116];
    assign P[1] = in1[116] ^ in2[116];
    assign G[2] = in1[115] & in2[115];
    assign P[2] = in1[115] ^ in2[115];
    assign G[3] = in1[114] & in2[114];
    assign P[3] = in1[114] ^ in2[114];
    assign G[4] = in1[113] & in2[113];
    assign P[4] = in1[113] ^ in2[113];
    assign G[5] = in1[112] & in2[112];
    assign P[5] = in1[112] ^ in2[112];
    assign G[6] = in1[111] & in2[111];
    assign P[6] = in1[111] ^ in2[111];
    assign G[7] = in1[110] & in2[110];
    assign P[7] = in1[110] ^ in2[110];
    assign G[8] = in1[109] & in2[109];
    assign P[8] = in1[109] ^ in2[109];
    assign G[9] = in1[108] & in2[108];
    assign P[9] = in1[108] ^ in2[108];
    assign G[10] = in1[107] & in2[107];
    assign P[10] = in1[107] ^ in2[107];
    assign G[11] = in1[106] & in2[106];
    assign P[11] = in1[106] ^ in2[106];
    assign G[12] = in1[105] & in2[105];
    assign P[12] = in1[105] ^ in2[105];
    assign G[13] = in1[104] & in2[104];
    assign P[13] = in1[104] ^ in2[104];
    assign G[14] = in1[103] & in2[103];
    assign P[14] = in1[103] ^ in2[103];
    assign G[15] = in1[102] & in2[102];
    assign P[15] = in1[102] ^ in2[102];
    assign G[16] = in1[101] & in2[101];
    assign P[16] = in1[101] ^ in2[101];
    assign G[17] = in1[100] & in2[100];
    assign P[17] = in1[100] ^ in2[100];
    assign G[18] = in1[99] & in2[99];
    assign P[18] = in1[99] ^ in2[99];
    assign G[19] = in1[98] & in2[98];
    assign P[19] = in1[98] ^ in2[98];
    assign G[20] = in1[97] & in2[97];
    assign P[20] = in1[97] ^ in2[97];
    assign G[21] = in1[96] & in2[96];
    assign P[21] = in1[96] ^ in2[96];
    assign G[22] = in1[95] & in2[95];
    assign P[22] = in1[95] ^ in2[95];
    assign G[23] = in1[94] & in2[94];
    assign P[23] = in1[94] ^ in2[94];
    assign G[24] = in1[93] & in2[93];
    assign P[24] = in1[93] ^ in2[93];
    assign G[25] = in1[92] & in2[92];
    assign P[25] = in1[92] ^ in2[92];
    assign G[26] = in1[91] & in2[91];
    assign P[26] = in1[91] ^ in2[91];
    assign G[27] = in1[90] & in2[90];
    assign P[27] = in1[90] ^ in2[90];
    assign G[28] = in1[89] & in2[89];
    assign P[28] = in1[89] ^ in2[89];
    assign G[29] = in1[88] & in2[88];
    assign P[29] = in1[88] ^ in2[88];
    assign G[30] = in1[87] & in2[87];
    assign P[30] = in1[87] ^ in2[87];
    assign G[31] = in1[86] & in2[86];
    assign P[31] = in1[86] ^ in2[86];
    assign G[32] = in1[85] & in2[85];
    assign P[32] = in1[85] ^ in2[85];
    assign G[33] = in1[84] & in2[84];
    assign P[33] = in1[84] ^ in2[84];
    assign G[34] = in1[83] & in2[83];
    assign P[34] = in1[83] ^ in2[83];
    assign G[35] = in1[82] & in2[82];
    assign P[35] = in1[82] ^ in2[82];
    assign G[36] = in1[81] & in2[81];
    assign P[36] = in1[81] ^ in2[81];
    assign G[37] = in1[80] & in2[80];
    assign P[37] = in1[80] ^ in2[80];
    assign G[38] = in1[79] & in2[79];
    assign P[38] = in1[79] ^ in2[79];
    assign G[39] = in1[78] & in2[78];
    assign P[39] = in1[78] ^ in2[78];
    assign G[40] = in1[77] & in2[77];
    assign P[40] = in1[77] ^ in2[77];
    assign G[41] = in1[76] & in2[76];
    assign P[41] = in1[76] ^ in2[76];
    assign G[42] = in1[75] & in2[75];
    assign P[42] = in1[75] ^ in2[75];
    assign G[43] = in1[74] & in2[74];
    assign P[43] = in1[74] ^ in2[74];
    assign G[44] = in1[73] & in2[73];
    assign P[44] = in1[73] ^ in2[73];
    assign G[45] = in1[72] & in2[72];
    assign P[45] = in1[72] ^ in2[72];
    assign G[46] = in1[71] & in2[71];
    assign P[46] = in1[71] ^ in2[71];
    assign G[47] = in1[70] & in2[70];
    assign P[47] = in1[70] ^ in2[70];
    assign G[48] = in1[69] & in2[69];
    assign P[48] = in1[69] ^ in2[69];
    assign G[49] = in1[68] & in2[68];
    assign P[49] = in1[68] ^ in2[68];
    assign G[50] = in1[67] & in2[67];
    assign P[50] = in1[67] ^ in2[67];
    assign G[51] = in1[66] & in2[66];
    assign P[51] = in1[66] ^ in2[66];
    assign G[52] = in1[65] & in2[65];
    assign P[52] = in1[65] ^ in2[65];
    assign G[53] = in1[64] & in2[64];
    assign P[53] = in1[64] ^ in2[64];
    assign G[54] = in1[63] & in2[63];
    assign P[54] = in1[63] ^ in2[63];
    assign G[55] = in1[62] & in2[62];
    assign P[55] = in1[62] ^ in2[62];
    assign G[56] = in1[61] & in2[61];
    assign P[56] = in1[61] ^ in2[61];
    assign G[57] = in1[60] & in2[60];
    assign P[57] = in1[60] ^ in2[60];
    assign G[58] = in1[59] & in2[59];
    assign P[58] = in1[59] ^ in2[59];
    assign G[59] = in1[58] & in2[58];
    assign P[59] = in1[58] ^ in2[58];
    assign G[60] = in1[57] & in2[57];
    assign P[60] = in1[57] ^ in2[57];
    assign G[61] = in1[56] & in2[56];
    assign P[61] = in1[56] ^ in2[56];
    assign G[62] = in1[55] & in2[55];
    assign P[62] = in1[55] ^ in2[55];
    assign G[63] = in1[54] & in2[54];
    assign P[63] = in1[54] ^ in2[54];
    assign G[64] = in1[53] & in2[53];
    assign P[64] = in1[53] ^ in2[53];
    assign G[65] = in1[52] & in2[52];
    assign P[65] = in1[52] ^ in2[52];
    assign G[66] = in1[51] & in2[51];
    assign P[66] = in1[51] ^ in2[51];
    assign G[67] = in1[50] & in2[50];
    assign P[67] = in1[50] ^ in2[50];
    assign G[68] = in1[49] & in2[49];
    assign P[68] = in1[49] ^ in2[49];
    assign G[69] = in1[48] & in2[48];
    assign P[69] = in1[48] ^ in2[48];
    assign G[70] = in1[47] & in2[47];
    assign P[70] = in1[47] ^ in2[47];
    assign G[71] = in1[46] & in2[46];
    assign P[71] = in1[46] ^ in2[46];
    assign G[72] = in1[45] & in2[45];
    assign P[72] = in1[45] ^ in2[45];
    assign G[73] = in1[44] & in2[44];
    assign P[73] = in1[44] ^ in2[44];
    assign G[74] = in1[43] & in2[43];
    assign P[74] = in1[43] ^ in2[43];
    assign G[75] = in1[42] & in2[42];
    assign P[75] = in1[42] ^ in2[42];
    assign G[76] = in1[41] & in2[41];
    assign P[76] = in1[41] ^ in2[41];
    assign G[77] = in1[40] & in2[40];
    assign P[77] = in1[40] ^ in2[40];
    assign G[78] = in1[39] & in2[39];
    assign P[78] = in1[39] ^ in2[39];
    assign G[79] = in1[38] & in2[38];
    assign P[79] = in1[38] ^ in2[38];
    assign G[80] = in1[37] & in2[37];
    assign P[80] = in1[37] ^ in2[37];
    assign G[81] = in1[36] & in2[36];
    assign P[81] = in1[36] ^ in2[36];
    assign G[82] = in1[35] & in2[35];
    assign P[82] = in1[35] ^ in2[35];
    assign G[83] = in1[34] & in2[34];
    assign P[83] = in1[34] ^ in2[34];
    assign G[84] = in1[33] & in2[33];
    assign P[84] = in1[33] ^ in2[33];
    assign G[85] = in1[32] & in2[32];
    assign P[85] = in1[32] ^ in2[32];
    assign G[86] = in1[31] & in2[31];
    assign P[86] = in1[31] ^ in2[31];
    assign G[87] = in1[30] & in2[30];
    assign P[87] = in1[30] ^ in2[30];
    assign G[88] = in1[29] & in2[29];
    assign P[88] = in1[29] ^ in2[29];
    assign G[89] = in1[28] & in2[28];
    assign P[89] = in1[28] ^ in2[28];
    assign G[90] = in1[27] & in2[27];
    assign P[90] = in1[27] ^ in2[27];
    assign G[91] = in1[26] & in2[26];
    assign P[91] = in1[26] ^ in2[26];
    assign G[92] = in1[25] & in2[25];
    assign P[92] = in1[25] ^ in2[25];
    assign G[93] = in1[24] & in2[24];
    assign P[93] = in1[24] ^ in2[24];
    assign G[94] = in1[23] & in2[23];
    assign P[94] = in1[23] ^ in2[23];
    assign G[95] = in1[22] & in2[22];
    assign P[95] = in1[22] ^ in2[22];
    assign G[96] = in1[21] & in2[21];
    assign P[96] = in1[21] ^ in2[21];
    assign G[97] = in1[20] & in2[20];
    assign P[97] = in1[20] ^ in2[20];
    assign G[98] = in1[19] & in2[19];
    assign P[98] = in1[19] ^ in2[19];
    assign G[99] = in1[18] & in2[18];
    assign P[99] = in1[18] ^ in2[18];
    assign G[100] = in1[17] & in2[17];
    assign P[100] = in1[17] ^ in2[17];
    assign G[101] = in1[16] & in2[16];
    assign P[101] = in1[16] ^ in2[16];
    assign G[102] = in1[15] & in2[15];
    assign P[102] = in1[15] ^ in2[15];
    assign G[103] = in1[14] & in2[14];
    assign P[103] = in1[14] ^ in2[14];
    assign G[104] = in1[13] & in2[13];
    assign P[104] = in1[13] ^ in2[13];
    assign G[105] = in1[12] & in2[12];
    assign P[105] = in1[12] ^ in2[12];
    assign G[106] = in1[11] & in2[11];
    assign P[106] = in1[11] ^ in2[11];
    assign G[107] = in1[10] & in2[10];
    assign P[107] = in1[10] ^ in2[10];
    assign G[108] = in1[9] & in2[9];
    assign P[108] = in1[9] ^ in2[9];
    assign G[109] = in1[8] & in2[8];
    assign P[109] = in1[8] ^ in2[8];
    assign G[110] = in1[7] & in2[7];
    assign P[110] = in1[7] ^ in2[7];
    assign G[111] = in1[6] & in2[6];
    assign P[111] = in1[6] ^ in2[6];
    assign G[112] = in1[5] & in2[5];
    assign P[112] = in1[5] ^ in2[5];
    assign G[113] = in1[4] & in2[4];
    assign P[113] = in1[4] ^ in2[4];
    assign G[114] = in1[3] & in2[3];
    assign P[114] = in1[3] ^ in2[3];
    assign G[115] = in1[2] & in2[2];
    assign P[115] = in1[2] ^ in2[2];
    assign G[116] = in1[1] & in2[1];
    assign P[116] = in1[1] ^ in2[1];
    assign G[117] = in1[0] & in2[0];
    assign P[117] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign cout = G[117] | (P[117] & C[117]);
    assign sum = P ^ C;
endmodule

module CLA_117(output [116:0] sum, output cout, input [116:0] in1, input [116:0] in2);

    wire[116:0] G;
    wire[116:0] C;
    wire[116:0] P;

    assign G[0] = in1[116] & in2[116];
    assign P[0] = in1[116] ^ in2[116];
    assign G[1] = in1[115] & in2[115];
    assign P[1] = in1[115] ^ in2[115];
    assign G[2] = in1[114] & in2[114];
    assign P[2] = in1[114] ^ in2[114];
    assign G[3] = in1[113] & in2[113];
    assign P[3] = in1[113] ^ in2[113];
    assign G[4] = in1[112] & in2[112];
    assign P[4] = in1[112] ^ in2[112];
    assign G[5] = in1[111] & in2[111];
    assign P[5] = in1[111] ^ in2[111];
    assign G[6] = in1[110] & in2[110];
    assign P[6] = in1[110] ^ in2[110];
    assign G[7] = in1[109] & in2[109];
    assign P[7] = in1[109] ^ in2[109];
    assign G[8] = in1[108] & in2[108];
    assign P[8] = in1[108] ^ in2[108];
    assign G[9] = in1[107] & in2[107];
    assign P[9] = in1[107] ^ in2[107];
    assign G[10] = in1[106] & in2[106];
    assign P[10] = in1[106] ^ in2[106];
    assign G[11] = in1[105] & in2[105];
    assign P[11] = in1[105] ^ in2[105];
    assign G[12] = in1[104] & in2[104];
    assign P[12] = in1[104] ^ in2[104];
    assign G[13] = in1[103] & in2[103];
    assign P[13] = in1[103] ^ in2[103];
    assign G[14] = in1[102] & in2[102];
    assign P[14] = in1[102] ^ in2[102];
    assign G[15] = in1[101] & in2[101];
    assign P[15] = in1[101] ^ in2[101];
    assign G[16] = in1[100] & in2[100];
    assign P[16] = in1[100] ^ in2[100];
    assign G[17] = in1[99] & in2[99];
    assign P[17] = in1[99] ^ in2[99];
    assign G[18] = in1[98] & in2[98];
    assign P[18] = in1[98] ^ in2[98];
    assign G[19] = in1[97] & in2[97];
    assign P[19] = in1[97] ^ in2[97];
    assign G[20] = in1[96] & in2[96];
    assign P[20] = in1[96] ^ in2[96];
    assign G[21] = in1[95] & in2[95];
    assign P[21] = in1[95] ^ in2[95];
    assign G[22] = in1[94] & in2[94];
    assign P[22] = in1[94] ^ in2[94];
    assign G[23] = in1[93] & in2[93];
    assign P[23] = in1[93] ^ in2[93];
    assign G[24] = in1[92] & in2[92];
    assign P[24] = in1[92] ^ in2[92];
    assign G[25] = in1[91] & in2[91];
    assign P[25] = in1[91] ^ in2[91];
    assign G[26] = in1[90] & in2[90];
    assign P[26] = in1[90] ^ in2[90];
    assign G[27] = in1[89] & in2[89];
    assign P[27] = in1[89] ^ in2[89];
    assign G[28] = in1[88] & in2[88];
    assign P[28] = in1[88] ^ in2[88];
    assign G[29] = in1[87] & in2[87];
    assign P[29] = in1[87] ^ in2[87];
    assign G[30] = in1[86] & in2[86];
    assign P[30] = in1[86] ^ in2[86];
    assign G[31] = in1[85] & in2[85];
    assign P[31] = in1[85] ^ in2[85];
    assign G[32] = in1[84] & in2[84];
    assign P[32] = in1[84] ^ in2[84];
    assign G[33] = in1[83] & in2[83];
    assign P[33] = in1[83] ^ in2[83];
    assign G[34] = in1[82] & in2[82];
    assign P[34] = in1[82] ^ in2[82];
    assign G[35] = in1[81] & in2[81];
    assign P[35] = in1[81] ^ in2[81];
    assign G[36] = in1[80] & in2[80];
    assign P[36] = in1[80] ^ in2[80];
    assign G[37] = in1[79] & in2[79];
    assign P[37] = in1[79] ^ in2[79];
    assign G[38] = in1[78] & in2[78];
    assign P[38] = in1[78] ^ in2[78];
    assign G[39] = in1[77] & in2[77];
    assign P[39] = in1[77] ^ in2[77];
    assign G[40] = in1[76] & in2[76];
    assign P[40] = in1[76] ^ in2[76];
    assign G[41] = in1[75] & in2[75];
    assign P[41] = in1[75] ^ in2[75];
    assign G[42] = in1[74] & in2[74];
    assign P[42] = in1[74] ^ in2[74];
    assign G[43] = in1[73] & in2[73];
    assign P[43] = in1[73] ^ in2[73];
    assign G[44] = in1[72] & in2[72];
    assign P[44] = in1[72] ^ in2[72];
    assign G[45] = in1[71] & in2[71];
    assign P[45] = in1[71] ^ in2[71];
    assign G[46] = in1[70] & in2[70];
    assign P[46] = in1[70] ^ in2[70];
    assign G[47] = in1[69] & in2[69];
    assign P[47] = in1[69] ^ in2[69];
    assign G[48] = in1[68] & in2[68];
    assign P[48] = in1[68] ^ in2[68];
    assign G[49] = in1[67] & in2[67];
    assign P[49] = in1[67] ^ in2[67];
    assign G[50] = in1[66] & in2[66];
    assign P[50] = in1[66] ^ in2[66];
    assign G[51] = in1[65] & in2[65];
    assign P[51] = in1[65] ^ in2[65];
    assign G[52] = in1[64] & in2[64];
    assign P[52] = in1[64] ^ in2[64];
    assign G[53] = in1[63] & in2[63];
    assign P[53] = in1[63] ^ in2[63];
    assign G[54] = in1[62] & in2[62];
    assign P[54] = in1[62] ^ in2[62];
    assign G[55] = in1[61] & in2[61];
    assign P[55] = in1[61] ^ in2[61];
    assign G[56] = in1[60] & in2[60];
    assign P[56] = in1[60] ^ in2[60];
    assign G[57] = in1[59] & in2[59];
    assign P[57] = in1[59] ^ in2[59];
    assign G[58] = in1[58] & in2[58];
    assign P[58] = in1[58] ^ in2[58];
    assign G[59] = in1[57] & in2[57];
    assign P[59] = in1[57] ^ in2[57];
    assign G[60] = in1[56] & in2[56];
    assign P[60] = in1[56] ^ in2[56];
    assign G[61] = in1[55] & in2[55];
    assign P[61] = in1[55] ^ in2[55];
    assign G[62] = in1[54] & in2[54];
    assign P[62] = in1[54] ^ in2[54];
    assign G[63] = in1[53] & in2[53];
    assign P[63] = in1[53] ^ in2[53];
    assign G[64] = in1[52] & in2[52];
    assign P[64] = in1[52] ^ in2[52];
    assign G[65] = in1[51] & in2[51];
    assign P[65] = in1[51] ^ in2[51];
    assign G[66] = in1[50] & in2[50];
    assign P[66] = in1[50] ^ in2[50];
    assign G[67] = in1[49] & in2[49];
    assign P[67] = in1[49] ^ in2[49];
    assign G[68] = in1[48] & in2[48];
    assign P[68] = in1[48] ^ in2[48];
    assign G[69] = in1[47] & in2[47];
    assign P[69] = in1[47] ^ in2[47];
    assign G[70] = in1[46] & in2[46];
    assign P[70] = in1[46] ^ in2[46];
    assign G[71] = in1[45] & in2[45];
    assign P[71] = in1[45] ^ in2[45];
    assign G[72] = in1[44] & in2[44];
    assign P[72] = in1[44] ^ in2[44];
    assign G[73] = in1[43] & in2[43];
    assign P[73] = in1[43] ^ in2[43];
    assign G[74] = in1[42] & in2[42];
    assign P[74] = in1[42] ^ in2[42];
    assign G[75] = in1[41] & in2[41];
    assign P[75] = in1[41] ^ in2[41];
    assign G[76] = in1[40] & in2[40];
    assign P[76] = in1[40] ^ in2[40];
    assign G[77] = in1[39] & in2[39];
    assign P[77] = in1[39] ^ in2[39];
    assign G[78] = in1[38] & in2[38];
    assign P[78] = in1[38] ^ in2[38];
    assign G[79] = in1[37] & in2[37];
    assign P[79] = in1[37] ^ in2[37];
    assign G[80] = in1[36] & in2[36];
    assign P[80] = in1[36] ^ in2[36];
    assign G[81] = in1[35] & in2[35];
    assign P[81] = in1[35] ^ in2[35];
    assign G[82] = in1[34] & in2[34];
    assign P[82] = in1[34] ^ in2[34];
    assign G[83] = in1[33] & in2[33];
    assign P[83] = in1[33] ^ in2[33];
    assign G[84] = in1[32] & in2[32];
    assign P[84] = in1[32] ^ in2[32];
    assign G[85] = in1[31] & in2[31];
    assign P[85] = in1[31] ^ in2[31];
    assign G[86] = in1[30] & in2[30];
    assign P[86] = in1[30] ^ in2[30];
    assign G[87] = in1[29] & in2[29];
    assign P[87] = in1[29] ^ in2[29];
    assign G[88] = in1[28] & in2[28];
    assign P[88] = in1[28] ^ in2[28];
    assign G[89] = in1[27] & in2[27];
    assign P[89] = in1[27] ^ in2[27];
    assign G[90] = in1[26] & in2[26];
    assign P[90] = in1[26] ^ in2[26];
    assign G[91] = in1[25] & in2[25];
    assign P[91] = in1[25] ^ in2[25];
    assign G[92] = in1[24] & in2[24];
    assign P[92] = in1[24] ^ in2[24];
    assign G[93] = in1[23] & in2[23];
    assign P[93] = in1[23] ^ in2[23];
    assign G[94] = in1[22] & in2[22];
    assign P[94] = in1[22] ^ in2[22];
    assign G[95] = in1[21] & in2[21];
    assign P[95] = in1[21] ^ in2[21];
    assign G[96] = in1[20] & in2[20];
    assign P[96] = in1[20] ^ in2[20];
    assign G[97] = in1[19] & in2[19];
    assign P[97] = in1[19] ^ in2[19];
    assign G[98] = in1[18] & in2[18];
    assign P[98] = in1[18] ^ in2[18];
    assign G[99] = in1[17] & in2[17];
    assign P[99] = in1[17] ^ in2[17];
    assign G[100] = in1[16] & in2[16];
    assign P[100] = in1[16] ^ in2[16];
    assign G[101] = in1[15] & in2[15];
    assign P[101] = in1[15] ^ in2[15];
    assign G[102] = in1[14] & in2[14];
    assign P[102] = in1[14] ^ in2[14];
    assign G[103] = in1[13] & in2[13];
    assign P[103] = in1[13] ^ in2[13];
    assign G[104] = in1[12] & in2[12];
    assign P[104] = in1[12] ^ in2[12];
    assign G[105] = in1[11] & in2[11];
    assign P[105] = in1[11] ^ in2[11];
    assign G[106] = in1[10] & in2[10];
    assign P[106] = in1[10] ^ in2[10];
    assign G[107] = in1[9] & in2[9];
    assign P[107] = in1[9] ^ in2[9];
    assign G[108] = in1[8] & in2[8];
    assign P[108] = in1[8] ^ in2[8];
    assign G[109] = in1[7] & in2[7];
    assign P[109] = in1[7] ^ in2[7];
    assign G[110] = in1[6] & in2[6];
    assign P[110] = in1[6] ^ in2[6];
    assign G[111] = in1[5] & in2[5];
    assign P[111] = in1[5] ^ in2[5];
    assign G[112] = in1[4] & in2[4];
    assign P[112] = in1[4] ^ in2[4];
    assign G[113] = in1[3] & in2[3];
    assign P[113] = in1[3] ^ in2[3];
    assign G[114] = in1[2] & in2[2];
    assign P[114] = in1[2] ^ in2[2];
    assign G[115] = in1[1] & in2[1];
    assign P[115] = in1[1] ^ in2[1];
    assign G[116] = in1[0] & in2[0];
    assign P[116] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign cout = G[116] | (P[116] & C[116]);
    assign sum = P ^ C;
endmodule

module CLA_116(output [115:0] sum, output cout, input [115:0] in1, input [115:0] in2);

    wire[115:0] G;
    wire[115:0] C;
    wire[115:0] P;

    assign G[0] = in1[115] & in2[115];
    assign P[0] = in1[115] ^ in2[115];
    assign G[1] = in1[114] & in2[114];
    assign P[1] = in1[114] ^ in2[114];
    assign G[2] = in1[113] & in2[113];
    assign P[2] = in1[113] ^ in2[113];
    assign G[3] = in1[112] & in2[112];
    assign P[3] = in1[112] ^ in2[112];
    assign G[4] = in1[111] & in2[111];
    assign P[4] = in1[111] ^ in2[111];
    assign G[5] = in1[110] & in2[110];
    assign P[5] = in1[110] ^ in2[110];
    assign G[6] = in1[109] & in2[109];
    assign P[6] = in1[109] ^ in2[109];
    assign G[7] = in1[108] & in2[108];
    assign P[7] = in1[108] ^ in2[108];
    assign G[8] = in1[107] & in2[107];
    assign P[8] = in1[107] ^ in2[107];
    assign G[9] = in1[106] & in2[106];
    assign P[9] = in1[106] ^ in2[106];
    assign G[10] = in1[105] & in2[105];
    assign P[10] = in1[105] ^ in2[105];
    assign G[11] = in1[104] & in2[104];
    assign P[11] = in1[104] ^ in2[104];
    assign G[12] = in1[103] & in2[103];
    assign P[12] = in1[103] ^ in2[103];
    assign G[13] = in1[102] & in2[102];
    assign P[13] = in1[102] ^ in2[102];
    assign G[14] = in1[101] & in2[101];
    assign P[14] = in1[101] ^ in2[101];
    assign G[15] = in1[100] & in2[100];
    assign P[15] = in1[100] ^ in2[100];
    assign G[16] = in1[99] & in2[99];
    assign P[16] = in1[99] ^ in2[99];
    assign G[17] = in1[98] & in2[98];
    assign P[17] = in1[98] ^ in2[98];
    assign G[18] = in1[97] & in2[97];
    assign P[18] = in1[97] ^ in2[97];
    assign G[19] = in1[96] & in2[96];
    assign P[19] = in1[96] ^ in2[96];
    assign G[20] = in1[95] & in2[95];
    assign P[20] = in1[95] ^ in2[95];
    assign G[21] = in1[94] & in2[94];
    assign P[21] = in1[94] ^ in2[94];
    assign G[22] = in1[93] & in2[93];
    assign P[22] = in1[93] ^ in2[93];
    assign G[23] = in1[92] & in2[92];
    assign P[23] = in1[92] ^ in2[92];
    assign G[24] = in1[91] & in2[91];
    assign P[24] = in1[91] ^ in2[91];
    assign G[25] = in1[90] & in2[90];
    assign P[25] = in1[90] ^ in2[90];
    assign G[26] = in1[89] & in2[89];
    assign P[26] = in1[89] ^ in2[89];
    assign G[27] = in1[88] & in2[88];
    assign P[27] = in1[88] ^ in2[88];
    assign G[28] = in1[87] & in2[87];
    assign P[28] = in1[87] ^ in2[87];
    assign G[29] = in1[86] & in2[86];
    assign P[29] = in1[86] ^ in2[86];
    assign G[30] = in1[85] & in2[85];
    assign P[30] = in1[85] ^ in2[85];
    assign G[31] = in1[84] & in2[84];
    assign P[31] = in1[84] ^ in2[84];
    assign G[32] = in1[83] & in2[83];
    assign P[32] = in1[83] ^ in2[83];
    assign G[33] = in1[82] & in2[82];
    assign P[33] = in1[82] ^ in2[82];
    assign G[34] = in1[81] & in2[81];
    assign P[34] = in1[81] ^ in2[81];
    assign G[35] = in1[80] & in2[80];
    assign P[35] = in1[80] ^ in2[80];
    assign G[36] = in1[79] & in2[79];
    assign P[36] = in1[79] ^ in2[79];
    assign G[37] = in1[78] & in2[78];
    assign P[37] = in1[78] ^ in2[78];
    assign G[38] = in1[77] & in2[77];
    assign P[38] = in1[77] ^ in2[77];
    assign G[39] = in1[76] & in2[76];
    assign P[39] = in1[76] ^ in2[76];
    assign G[40] = in1[75] & in2[75];
    assign P[40] = in1[75] ^ in2[75];
    assign G[41] = in1[74] & in2[74];
    assign P[41] = in1[74] ^ in2[74];
    assign G[42] = in1[73] & in2[73];
    assign P[42] = in1[73] ^ in2[73];
    assign G[43] = in1[72] & in2[72];
    assign P[43] = in1[72] ^ in2[72];
    assign G[44] = in1[71] & in2[71];
    assign P[44] = in1[71] ^ in2[71];
    assign G[45] = in1[70] & in2[70];
    assign P[45] = in1[70] ^ in2[70];
    assign G[46] = in1[69] & in2[69];
    assign P[46] = in1[69] ^ in2[69];
    assign G[47] = in1[68] & in2[68];
    assign P[47] = in1[68] ^ in2[68];
    assign G[48] = in1[67] & in2[67];
    assign P[48] = in1[67] ^ in2[67];
    assign G[49] = in1[66] & in2[66];
    assign P[49] = in1[66] ^ in2[66];
    assign G[50] = in1[65] & in2[65];
    assign P[50] = in1[65] ^ in2[65];
    assign G[51] = in1[64] & in2[64];
    assign P[51] = in1[64] ^ in2[64];
    assign G[52] = in1[63] & in2[63];
    assign P[52] = in1[63] ^ in2[63];
    assign G[53] = in1[62] & in2[62];
    assign P[53] = in1[62] ^ in2[62];
    assign G[54] = in1[61] & in2[61];
    assign P[54] = in1[61] ^ in2[61];
    assign G[55] = in1[60] & in2[60];
    assign P[55] = in1[60] ^ in2[60];
    assign G[56] = in1[59] & in2[59];
    assign P[56] = in1[59] ^ in2[59];
    assign G[57] = in1[58] & in2[58];
    assign P[57] = in1[58] ^ in2[58];
    assign G[58] = in1[57] & in2[57];
    assign P[58] = in1[57] ^ in2[57];
    assign G[59] = in1[56] & in2[56];
    assign P[59] = in1[56] ^ in2[56];
    assign G[60] = in1[55] & in2[55];
    assign P[60] = in1[55] ^ in2[55];
    assign G[61] = in1[54] & in2[54];
    assign P[61] = in1[54] ^ in2[54];
    assign G[62] = in1[53] & in2[53];
    assign P[62] = in1[53] ^ in2[53];
    assign G[63] = in1[52] & in2[52];
    assign P[63] = in1[52] ^ in2[52];
    assign G[64] = in1[51] & in2[51];
    assign P[64] = in1[51] ^ in2[51];
    assign G[65] = in1[50] & in2[50];
    assign P[65] = in1[50] ^ in2[50];
    assign G[66] = in1[49] & in2[49];
    assign P[66] = in1[49] ^ in2[49];
    assign G[67] = in1[48] & in2[48];
    assign P[67] = in1[48] ^ in2[48];
    assign G[68] = in1[47] & in2[47];
    assign P[68] = in1[47] ^ in2[47];
    assign G[69] = in1[46] & in2[46];
    assign P[69] = in1[46] ^ in2[46];
    assign G[70] = in1[45] & in2[45];
    assign P[70] = in1[45] ^ in2[45];
    assign G[71] = in1[44] & in2[44];
    assign P[71] = in1[44] ^ in2[44];
    assign G[72] = in1[43] & in2[43];
    assign P[72] = in1[43] ^ in2[43];
    assign G[73] = in1[42] & in2[42];
    assign P[73] = in1[42] ^ in2[42];
    assign G[74] = in1[41] & in2[41];
    assign P[74] = in1[41] ^ in2[41];
    assign G[75] = in1[40] & in2[40];
    assign P[75] = in1[40] ^ in2[40];
    assign G[76] = in1[39] & in2[39];
    assign P[76] = in1[39] ^ in2[39];
    assign G[77] = in1[38] & in2[38];
    assign P[77] = in1[38] ^ in2[38];
    assign G[78] = in1[37] & in2[37];
    assign P[78] = in1[37] ^ in2[37];
    assign G[79] = in1[36] & in2[36];
    assign P[79] = in1[36] ^ in2[36];
    assign G[80] = in1[35] & in2[35];
    assign P[80] = in1[35] ^ in2[35];
    assign G[81] = in1[34] & in2[34];
    assign P[81] = in1[34] ^ in2[34];
    assign G[82] = in1[33] & in2[33];
    assign P[82] = in1[33] ^ in2[33];
    assign G[83] = in1[32] & in2[32];
    assign P[83] = in1[32] ^ in2[32];
    assign G[84] = in1[31] & in2[31];
    assign P[84] = in1[31] ^ in2[31];
    assign G[85] = in1[30] & in2[30];
    assign P[85] = in1[30] ^ in2[30];
    assign G[86] = in1[29] & in2[29];
    assign P[86] = in1[29] ^ in2[29];
    assign G[87] = in1[28] & in2[28];
    assign P[87] = in1[28] ^ in2[28];
    assign G[88] = in1[27] & in2[27];
    assign P[88] = in1[27] ^ in2[27];
    assign G[89] = in1[26] & in2[26];
    assign P[89] = in1[26] ^ in2[26];
    assign G[90] = in1[25] & in2[25];
    assign P[90] = in1[25] ^ in2[25];
    assign G[91] = in1[24] & in2[24];
    assign P[91] = in1[24] ^ in2[24];
    assign G[92] = in1[23] & in2[23];
    assign P[92] = in1[23] ^ in2[23];
    assign G[93] = in1[22] & in2[22];
    assign P[93] = in1[22] ^ in2[22];
    assign G[94] = in1[21] & in2[21];
    assign P[94] = in1[21] ^ in2[21];
    assign G[95] = in1[20] & in2[20];
    assign P[95] = in1[20] ^ in2[20];
    assign G[96] = in1[19] & in2[19];
    assign P[96] = in1[19] ^ in2[19];
    assign G[97] = in1[18] & in2[18];
    assign P[97] = in1[18] ^ in2[18];
    assign G[98] = in1[17] & in2[17];
    assign P[98] = in1[17] ^ in2[17];
    assign G[99] = in1[16] & in2[16];
    assign P[99] = in1[16] ^ in2[16];
    assign G[100] = in1[15] & in2[15];
    assign P[100] = in1[15] ^ in2[15];
    assign G[101] = in1[14] & in2[14];
    assign P[101] = in1[14] ^ in2[14];
    assign G[102] = in1[13] & in2[13];
    assign P[102] = in1[13] ^ in2[13];
    assign G[103] = in1[12] & in2[12];
    assign P[103] = in1[12] ^ in2[12];
    assign G[104] = in1[11] & in2[11];
    assign P[104] = in1[11] ^ in2[11];
    assign G[105] = in1[10] & in2[10];
    assign P[105] = in1[10] ^ in2[10];
    assign G[106] = in1[9] & in2[9];
    assign P[106] = in1[9] ^ in2[9];
    assign G[107] = in1[8] & in2[8];
    assign P[107] = in1[8] ^ in2[8];
    assign G[108] = in1[7] & in2[7];
    assign P[108] = in1[7] ^ in2[7];
    assign G[109] = in1[6] & in2[6];
    assign P[109] = in1[6] ^ in2[6];
    assign G[110] = in1[5] & in2[5];
    assign P[110] = in1[5] ^ in2[5];
    assign G[111] = in1[4] & in2[4];
    assign P[111] = in1[4] ^ in2[4];
    assign G[112] = in1[3] & in2[3];
    assign P[112] = in1[3] ^ in2[3];
    assign G[113] = in1[2] & in2[2];
    assign P[113] = in1[2] ^ in2[2];
    assign G[114] = in1[1] & in2[1];
    assign P[114] = in1[1] ^ in2[1];
    assign G[115] = in1[0] & in2[0];
    assign P[115] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign cout = G[115] | (P[115] & C[115]);
    assign sum = P ^ C;
endmodule

module CLA_115(output [114:0] sum, output cout, input [114:0] in1, input [114:0] in2);

    wire[114:0] G;
    wire[114:0] C;
    wire[114:0] P;

    assign G[0] = in1[114] & in2[114];
    assign P[0] = in1[114] ^ in2[114];
    assign G[1] = in1[113] & in2[113];
    assign P[1] = in1[113] ^ in2[113];
    assign G[2] = in1[112] & in2[112];
    assign P[2] = in1[112] ^ in2[112];
    assign G[3] = in1[111] & in2[111];
    assign P[3] = in1[111] ^ in2[111];
    assign G[4] = in1[110] & in2[110];
    assign P[4] = in1[110] ^ in2[110];
    assign G[5] = in1[109] & in2[109];
    assign P[5] = in1[109] ^ in2[109];
    assign G[6] = in1[108] & in2[108];
    assign P[6] = in1[108] ^ in2[108];
    assign G[7] = in1[107] & in2[107];
    assign P[7] = in1[107] ^ in2[107];
    assign G[8] = in1[106] & in2[106];
    assign P[8] = in1[106] ^ in2[106];
    assign G[9] = in1[105] & in2[105];
    assign P[9] = in1[105] ^ in2[105];
    assign G[10] = in1[104] & in2[104];
    assign P[10] = in1[104] ^ in2[104];
    assign G[11] = in1[103] & in2[103];
    assign P[11] = in1[103] ^ in2[103];
    assign G[12] = in1[102] & in2[102];
    assign P[12] = in1[102] ^ in2[102];
    assign G[13] = in1[101] & in2[101];
    assign P[13] = in1[101] ^ in2[101];
    assign G[14] = in1[100] & in2[100];
    assign P[14] = in1[100] ^ in2[100];
    assign G[15] = in1[99] & in2[99];
    assign P[15] = in1[99] ^ in2[99];
    assign G[16] = in1[98] & in2[98];
    assign P[16] = in1[98] ^ in2[98];
    assign G[17] = in1[97] & in2[97];
    assign P[17] = in1[97] ^ in2[97];
    assign G[18] = in1[96] & in2[96];
    assign P[18] = in1[96] ^ in2[96];
    assign G[19] = in1[95] & in2[95];
    assign P[19] = in1[95] ^ in2[95];
    assign G[20] = in1[94] & in2[94];
    assign P[20] = in1[94] ^ in2[94];
    assign G[21] = in1[93] & in2[93];
    assign P[21] = in1[93] ^ in2[93];
    assign G[22] = in1[92] & in2[92];
    assign P[22] = in1[92] ^ in2[92];
    assign G[23] = in1[91] & in2[91];
    assign P[23] = in1[91] ^ in2[91];
    assign G[24] = in1[90] & in2[90];
    assign P[24] = in1[90] ^ in2[90];
    assign G[25] = in1[89] & in2[89];
    assign P[25] = in1[89] ^ in2[89];
    assign G[26] = in1[88] & in2[88];
    assign P[26] = in1[88] ^ in2[88];
    assign G[27] = in1[87] & in2[87];
    assign P[27] = in1[87] ^ in2[87];
    assign G[28] = in1[86] & in2[86];
    assign P[28] = in1[86] ^ in2[86];
    assign G[29] = in1[85] & in2[85];
    assign P[29] = in1[85] ^ in2[85];
    assign G[30] = in1[84] & in2[84];
    assign P[30] = in1[84] ^ in2[84];
    assign G[31] = in1[83] & in2[83];
    assign P[31] = in1[83] ^ in2[83];
    assign G[32] = in1[82] & in2[82];
    assign P[32] = in1[82] ^ in2[82];
    assign G[33] = in1[81] & in2[81];
    assign P[33] = in1[81] ^ in2[81];
    assign G[34] = in1[80] & in2[80];
    assign P[34] = in1[80] ^ in2[80];
    assign G[35] = in1[79] & in2[79];
    assign P[35] = in1[79] ^ in2[79];
    assign G[36] = in1[78] & in2[78];
    assign P[36] = in1[78] ^ in2[78];
    assign G[37] = in1[77] & in2[77];
    assign P[37] = in1[77] ^ in2[77];
    assign G[38] = in1[76] & in2[76];
    assign P[38] = in1[76] ^ in2[76];
    assign G[39] = in1[75] & in2[75];
    assign P[39] = in1[75] ^ in2[75];
    assign G[40] = in1[74] & in2[74];
    assign P[40] = in1[74] ^ in2[74];
    assign G[41] = in1[73] & in2[73];
    assign P[41] = in1[73] ^ in2[73];
    assign G[42] = in1[72] & in2[72];
    assign P[42] = in1[72] ^ in2[72];
    assign G[43] = in1[71] & in2[71];
    assign P[43] = in1[71] ^ in2[71];
    assign G[44] = in1[70] & in2[70];
    assign P[44] = in1[70] ^ in2[70];
    assign G[45] = in1[69] & in2[69];
    assign P[45] = in1[69] ^ in2[69];
    assign G[46] = in1[68] & in2[68];
    assign P[46] = in1[68] ^ in2[68];
    assign G[47] = in1[67] & in2[67];
    assign P[47] = in1[67] ^ in2[67];
    assign G[48] = in1[66] & in2[66];
    assign P[48] = in1[66] ^ in2[66];
    assign G[49] = in1[65] & in2[65];
    assign P[49] = in1[65] ^ in2[65];
    assign G[50] = in1[64] & in2[64];
    assign P[50] = in1[64] ^ in2[64];
    assign G[51] = in1[63] & in2[63];
    assign P[51] = in1[63] ^ in2[63];
    assign G[52] = in1[62] & in2[62];
    assign P[52] = in1[62] ^ in2[62];
    assign G[53] = in1[61] & in2[61];
    assign P[53] = in1[61] ^ in2[61];
    assign G[54] = in1[60] & in2[60];
    assign P[54] = in1[60] ^ in2[60];
    assign G[55] = in1[59] & in2[59];
    assign P[55] = in1[59] ^ in2[59];
    assign G[56] = in1[58] & in2[58];
    assign P[56] = in1[58] ^ in2[58];
    assign G[57] = in1[57] & in2[57];
    assign P[57] = in1[57] ^ in2[57];
    assign G[58] = in1[56] & in2[56];
    assign P[58] = in1[56] ^ in2[56];
    assign G[59] = in1[55] & in2[55];
    assign P[59] = in1[55] ^ in2[55];
    assign G[60] = in1[54] & in2[54];
    assign P[60] = in1[54] ^ in2[54];
    assign G[61] = in1[53] & in2[53];
    assign P[61] = in1[53] ^ in2[53];
    assign G[62] = in1[52] & in2[52];
    assign P[62] = in1[52] ^ in2[52];
    assign G[63] = in1[51] & in2[51];
    assign P[63] = in1[51] ^ in2[51];
    assign G[64] = in1[50] & in2[50];
    assign P[64] = in1[50] ^ in2[50];
    assign G[65] = in1[49] & in2[49];
    assign P[65] = in1[49] ^ in2[49];
    assign G[66] = in1[48] & in2[48];
    assign P[66] = in1[48] ^ in2[48];
    assign G[67] = in1[47] & in2[47];
    assign P[67] = in1[47] ^ in2[47];
    assign G[68] = in1[46] & in2[46];
    assign P[68] = in1[46] ^ in2[46];
    assign G[69] = in1[45] & in2[45];
    assign P[69] = in1[45] ^ in2[45];
    assign G[70] = in1[44] & in2[44];
    assign P[70] = in1[44] ^ in2[44];
    assign G[71] = in1[43] & in2[43];
    assign P[71] = in1[43] ^ in2[43];
    assign G[72] = in1[42] & in2[42];
    assign P[72] = in1[42] ^ in2[42];
    assign G[73] = in1[41] & in2[41];
    assign P[73] = in1[41] ^ in2[41];
    assign G[74] = in1[40] & in2[40];
    assign P[74] = in1[40] ^ in2[40];
    assign G[75] = in1[39] & in2[39];
    assign P[75] = in1[39] ^ in2[39];
    assign G[76] = in1[38] & in2[38];
    assign P[76] = in1[38] ^ in2[38];
    assign G[77] = in1[37] & in2[37];
    assign P[77] = in1[37] ^ in2[37];
    assign G[78] = in1[36] & in2[36];
    assign P[78] = in1[36] ^ in2[36];
    assign G[79] = in1[35] & in2[35];
    assign P[79] = in1[35] ^ in2[35];
    assign G[80] = in1[34] & in2[34];
    assign P[80] = in1[34] ^ in2[34];
    assign G[81] = in1[33] & in2[33];
    assign P[81] = in1[33] ^ in2[33];
    assign G[82] = in1[32] & in2[32];
    assign P[82] = in1[32] ^ in2[32];
    assign G[83] = in1[31] & in2[31];
    assign P[83] = in1[31] ^ in2[31];
    assign G[84] = in1[30] & in2[30];
    assign P[84] = in1[30] ^ in2[30];
    assign G[85] = in1[29] & in2[29];
    assign P[85] = in1[29] ^ in2[29];
    assign G[86] = in1[28] & in2[28];
    assign P[86] = in1[28] ^ in2[28];
    assign G[87] = in1[27] & in2[27];
    assign P[87] = in1[27] ^ in2[27];
    assign G[88] = in1[26] & in2[26];
    assign P[88] = in1[26] ^ in2[26];
    assign G[89] = in1[25] & in2[25];
    assign P[89] = in1[25] ^ in2[25];
    assign G[90] = in1[24] & in2[24];
    assign P[90] = in1[24] ^ in2[24];
    assign G[91] = in1[23] & in2[23];
    assign P[91] = in1[23] ^ in2[23];
    assign G[92] = in1[22] & in2[22];
    assign P[92] = in1[22] ^ in2[22];
    assign G[93] = in1[21] & in2[21];
    assign P[93] = in1[21] ^ in2[21];
    assign G[94] = in1[20] & in2[20];
    assign P[94] = in1[20] ^ in2[20];
    assign G[95] = in1[19] & in2[19];
    assign P[95] = in1[19] ^ in2[19];
    assign G[96] = in1[18] & in2[18];
    assign P[96] = in1[18] ^ in2[18];
    assign G[97] = in1[17] & in2[17];
    assign P[97] = in1[17] ^ in2[17];
    assign G[98] = in1[16] & in2[16];
    assign P[98] = in1[16] ^ in2[16];
    assign G[99] = in1[15] & in2[15];
    assign P[99] = in1[15] ^ in2[15];
    assign G[100] = in1[14] & in2[14];
    assign P[100] = in1[14] ^ in2[14];
    assign G[101] = in1[13] & in2[13];
    assign P[101] = in1[13] ^ in2[13];
    assign G[102] = in1[12] & in2[12];
    assign P[102] = in1[12] ^ in2[12];
    assign G[103] = in1[11] & in2[11];
    assign P[103] = in1[11] ^ in2[11];
    assign G[104] = in1[10] & in2[10];
    assign P[104] = in1[10] ^ in2[10];
    assign G[105] = in1[9] & in2[9];
    assign P[105] = in1[9] ^ in2[9];
    assign G[106] = in1[8] & in2[8];
    assign P[106] = in1[8] ^ in2[8];
    assign G[107] = in1[7] & in2[7];
    assign P[107] = in1[7] ^ in2[7];
    assign G[108] = in1[6] & in2[6];
    assign P[108] = in1[6] ^ in2[6];
    assign G[109] = in1[5] & in2[5];
    assign P[109] = in1[5] ^ in2[5];
    assign G[110] = in1[4] & in2[4];
    assign P[110] = in1[4] ^ in2[4];
    assign G[111] = in1[3] & in2[3];
    assign P[111] = in1[3] ^ in2[3];
    assign G[112] = in1[2] & in2[2];
    assign P[112] = in1[2] ^ in2[2];
    assign G[113] = in1[1] & in2[1];
    assign P[113] = in1[1] ^ in2[1];
    assign G[114] = in1[0] & in2[0];
    assign P[114] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign cout = G[114] | (P[114] & C[114]);
    assign sum = P ^ C;
endmodule

module CLA_114(output [113:0] sum, output cout, input [113:0] in1, input [113:0] in2);

    wire[113:0] G;
    wire[113:0] C;
    wire[113:0] P;

    assign G[0] = in1[113] & in2[113];
    assign P[0] = in1[113] ^ in2[113];
    assign G[1] = in1[112] & in2[112];
    assign P[1] = in1[112] ^ in2[112];
    assign G[2] = in1[111] & in2[111];
    assign P[2] = in1[111] ^ in2[111];
    assign G[3] = in1[110] & in2[110];
    assign P[3] = in1[110] ^ in2[110];
    assign G[4] = in1[109] & in2[109];
    assign P[4] = in1[109] ^ in2[109];
    assign G[5] = in1[108] & in2[108];
    assign P[5] = in1[108] ^ in2[108];
    assign G[6] = in1[107] & in2[107];
    assign P[6] = in1[107] ^ in2[107];
    assign G[7] = in1[106] & in2[106];
    assign P[7] = in1[106] ^ in2[106];
    assign G[8] = in1[105] & in2[105];
    assign P[8] = in1[105] ^ in2[105];
    assign G[9] = in1[104] & in2[104];
    assign P[9] = in1[104] ^ in2[104];
    assign G[10] = in1[103] & in2[103];
    assign P[10] = in1[103] ^ in2[103];
    assign G[11] = in1[102] & in2[102];
    assign P[11] = in1[102] ^ in2[102];
    assign G[12] = in1[101] & in2[101];
    assign P[12] = in1[101] ^ in2[101];
    assign G[13] = in1[100] & in2[100];
    assign P[13] = in1[100] ^ in2[100];
    assign G[14] = in1[99] & in2[99];
    assign P[14] = in1[99] ^ in2[99];
    assign G[15] = in1[98] & in2[98];
    assign P[15] = in1[98] ^ in2[98];
    assign G[16] = in1[97] & in2[97];
    assign P[16] = in1[97] ^ in2[97];
    assign G[17] = in1[96] & in2[96];
    assign P[17] = in1[96] ^ in2[96];
    assign G[18] = in1[95] & in2[95];
    assign P[18] = in1[95] ^ in2[95];
    assign G[19] = in1[94] & in2[94];
    assign P[19] = in1[94] ^ in2[94];
    assign G[20] = in1[93] & in2[93];
    assign P[20] = in1[93] ^ in2[93];
    assign G[21] = in1[92] & in2[92];
    assign P[21] = in1[92] ^ in2[92];
    assign G[22] = in1[91] & in2[91];
    assign P[22] = in1[91] ^ in2[91];
    assign G[23] = in1[90] & in2[90];
    assign P[23] = in1[90] ^ in2[90];
    assign G[24] = in1[89] & in2[89];
    assign P[24] = in1[89] ^ in2[89];
    assign G[25] = in1[88] & in2[88];
    assign P[25] = in1[88] ^ in2[88];
    assign G[26] = in1[87] & in2[87];
    assign P[26] = in1[87] ^ in2[87];
    assign G[27] = in1[86] & in2[86];
    assign P[27] = in1[86] ^ in2[86];
    assign G[28] = in1[85] & in2[85];
    assign P[28] = in1[85] ^ in2[85];
    assign G[29] = in1[84] & in2[84];
    assign P[29] = in1[84] ^ in2[84];
    assign G[30] = in1[83] & in2[83];
    assign P[30] = in1[83] ^ in2[83];
    assign G[31] = in1[82] & in2[82];
    assign P[31] = in1[82] ^ in2[82];
    assign G[32] = in1[81] & in2[81];
    assign P[32] = in1[81] ^ in2[81];
    assign G[33] = in1[80] & in2[80];
    assign P[33] = in1[80] ^ in2[80];
    assign G[34] = in1[79] & in2[79];
    assign P[34] = in1[79] ^ in2[79];
    assign G[35] = in1[78] & in2[78];
    assign P[35] = in1[78] ^ in2[78];
    assign G[36] = in1[77] & in2[77];
    assign P[36] = in1[77] ^ in2[77];
    assign G[37] = in1[76] & in2[76];
    assign P[37] = in1[76] ^ in2[76];
    assign G[38] = in1[75] & in2[75];
    assign P[38] = in1[75] ^ in2[75];
    assign G[39] = in1[74] & in2[74];
    assign P[39] = in1[74] ^ in2[74];
    assign G[40] = in1[73] & in2[73];
    assign P[40] = in1[73] ^ in2[73];
    assign G[41] = in1[72] & in2[72];
    assign P[41] = in1[72] ^ in2[72];
    assign G[42] = in1[71] & in2[71];
    assign P[42] = in1[71] ^ in2[71];
    assign G[43] = in1[70] & in2[70];
    assign P[43] = in1[70] ^ in2[70];
    assign G[44] = in1[69] & in2[69];
    assign P[44] = in1[69] ^ in2[69];
    assign G[45] = in1[68] & in2[68];
    assign P[45] = in1[68] ^ in2[68];
    assign G[46] = in1[67] & in2[67];
    assign P[46] = in1[67] ^ in2[67];
    assign G[47] = in1[66] & in2[66];
    assign P[47] = in1[66] ^ in2[66];
    assign G[48] = in1[65] & in2[65];
    assign P[48] = in1[65] ^ in2[65];
    assign G[49] = in1[64] & in2[64];
    assign P[49] = in1[64] ^ in2[64];
    assign G[50] = in1[63] & in2[63];
    assign P[50] = in1[63] ^ in2[63];
    assign G[51] = in1[62] & in2[62];
    assign P[51] = in1[62] ^ in2[62];
    assign G[52] = in1[61] & in2[61];
    assign P[52] = in1[61] ^ in2[61];
    assign G[53] = in1[60] & in2[60];
    assign P[53] = in1[60] ^ in2[60];
    assign G[54] = in1[59] & in2[59];
    assign P[54] = in1[59] ^ in2[59];
    assign G[55] = in1[58] & in2[58];
    assign P[55] = in1[58] ^ in2[58];
    assign G[56] = in1[57] & in2[57];
    assign P[56] = in1[57] ^ in2[57];
    assign G[57] = in1[56] & in2[56];
    assign P[57] = in1[56] ^ in2[56];
    assign G[58] = in1[55] & in2[55];
    assign P[58] = in1[55] ^ in2[55];
    assign G[59] = in1[54] & in2[54];
    assign P[59] = in1[54] ^ in2[54];
    assign G[60] = in1[53] & in2[53];
    assign P[60] = in1[53] ^ in2[53];
    assign G[61] = in1[52] & in2[52];
    assign P[61] = in1[52] ^ in2[52];
    assign G[62] = in1[51] & in2[51];
    assign P[62] = in1[51] ^ in2[51];
    assign G[63] = in1[50] & in2[50];
    assign P[63] = in1[50] ^ in2[50];
    assign G[64] = in1[49] & in2[49];
    assign P[64] = in1[49] ^ in2[49];
    assign G[65] = in1[48] & in2[48];
    assign P[65] = in1[48] ^ in2[48];
    assign G[66] = in1[47] & in2[47];
    assign P[66] = in1[47] ^ in2[47];
    assign G[67] = in1[46] & in2[46];
    assign P[67] = in1[46] ^ in2[46];
    assign G[68] = in1[45] & in2[45];
    assign P[68] = in1[45] ^ in2[45];
    assign G[69] = in1[44] & in2[44];
    assign P[69] = in1[44] ^ in2[44];
    assign G[70] = in1[43] & in2[43];
    assign P[70] = in1[43] ^ in2[43];
    assign G[71] = in1[42] & in2[42];
    assign P[71] = in1[42] ^ in2[42];
    assign G[72] = in1[41] & in2[41];
    assign P[72] = in1[41] ^ in2[41];
    assign G[73] = in1[40] & in2[40];
    assign P[73] = in1[40] ^ in2[40];
    assign G[74] = in1[39] & in2[39];
    assign P[74] = in1[39] ^ in2[39];
    assign G[75] = in1[38] & in2[38];
    assign P[75] = in1[38] ^ in2[38];
    assign G[76] = in1[37] & in2[37];
    assign P[76] = in1[37] ^ in2[37];
    assign G[77] = in1[36] & in2[36];
    assign P[77] = in1[36] ^ in2[36];
    assign G[78] = in1[35] & in2[35];
    assign P[78] = in1[35] ^ in2[35];
    assign G[79] = in1[34] & in2[34];
    assign P[79] = in1[34] ^ in2[34];
    assign G[80] = in1[33] & in2[33];
    assign P[80] = in1[33] ^ in2[33];
    assign G[81] = in1[32] & in2[32];
    assign P[81] = in1[32] ^ in2[32];
    assign G[82] = in1[31] & in2[31];
    assign P[82] = in1[31] ^ in2[31];
    assign G[83] = in1[30] & in2[30];
    assign P[83] = in1[30] ^ in2[30];
    assign G[84] = in1[29] & in2[29];
    assign P[84] = in1[29] ^ in2[29];
    assign G[85] = in1[28] & in2[28];
    assign P[85] = in1[28] ^ in2[28];
    assign G[86] = in1[27] & in2[27];
    assign P[86] = in1[27] ^ in2[27];
    assign G[87] = in1[26] & in2[26];
    assign P[87] = in1[26] ^ in2[26];
    assign G[88] = in1[25] & in2[25];
    assign P[88] = in1[25] ^ in2[25];
    assign G[89] = in1[24] & in2[24];
    assign P[89] = in1[24] ^ in2[24];
    assign G[90] = in1[23] & in2[23];
    assign P[90] = in1[23] ^ in2[23];
    assign G[91] = in1[22] & in2[22];
    assign P[91] = in1[22] ^ in2[22];
    assign G[92] = in1[21] & in2[21];
    assign P[92] = in1[21] ^ in2[21];
    assign G[93] = in1[20] & in2[20];
    assign P[93] = in1[20] ^ in2[20];
    assign G[94] = in1[19] & in2[19];
    assign P[94] = in1[19] ^ in2[19];
    assign G[95] = in1[18] & in2[18];
    assign P[95] = in1[18] ^ in2[18];
    assign G[96] = in1[17] & in2[17];
    assign P[96] = in1[17] ^ in2[17];
    assign G[97] = in1[16] & in2[16];
    assign P[97] = in1[16] ^ in2[16];
    assign G[98] = in1[15] & in2[15];
    assign P[98] = in1[15] ^ in2[15];
    assign G[99] = in1[14] & in2[14];
    assign P[99] = in1[14] ^ in2[14];
    assign G[100] = in1[13] & in2[13];
    assign P[100] = in1[13] ^ in2[13];
    assign G[101] = in1[12] & in2[12];
    assign P[101] = in1[12] ^ in2[12];
    assign G[102] = in1[11] & in2[11];
    assign P[102] = in1[11] ^ in2[11];
    assign G[103] = in1[10] & in2[10];
    assign P[103] = in1[10] ^ in2[10];
    assign G[104] = in1[9] & in2[9];
    assign P[104] = in1[9] ^ in2[9];
    assign G[105] = in1[8] & in2[8];
    assign P[105] = in1[8] ^ in2[8];
    assign G[106] = in1[7] & in2[7];
    assign P[106] = in1[7] ^ in2[7];
    assign G[107] = in1[6] & in2[6];
    assign P[107] = in1[6] ^ in2[6];
    assign G[108] = in1[5] & in2[5];
    assign P[108] = in1[5] ^ in2[5];
    assign G[109] = in1[4] & in2[4];
    assign P[109] = in1[4] ^ in2[4];
    assign G[110] = in1[3] & in2[3];
    assign P[110] = in1[3] ^ in2[3];
    assign G[111] = in1[2] & in2[2];
    assign P[111] = in1[2] ^ in2[2];
    assign G[112] = in1[1] & in2[1];
    assign P[112] = in1[1] ^ in2[1];
    assign G[113] = in1[0] & in2[0];
    assign P[113] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign cout = G[113] | (P[113] & C[113]);
    assign sum = P ^ C;
endmodule

module CLA_113(output [112:0] sum, output cout, input [112:0] in1, input [112:0] in2);

    wire[112:0] G;
    wire[112:0] C;
    wire[112:0] P;

    assign G[0] = in1[112] & in2[112];
    assign P[0] = in1[112] ^ in2[112];
    assign G[1] = in1[111] & in2[111];
    assign P[1] = in1[111] ^ in2[111];
    assign G[2] = in1[110] & in2[110];
    assign P[2] = in1[110] ^ in2[110];
    assign G[3] = in1[109] & in2[109];
    assign P[3] = in1[109] ^ in2[109];
    assign G[4] = in1[108] & in2[108];
    assign P[4] = in1[108] ^ in2[108];
    assign G[5] = in1[107] & in2[107];
    assign P[5] = in1[107] ^ in2[107];
    assign G[6] = in1[106] & in2[106];
    assign P[6] = in1[106] ^ in2[106];
    assign G[7] = in1[105] & in2[105];
    assign P[7] = in1[105] ^ in2[105];
    assign G[8] = in1[104] & in2[104];
    assign P[8] = in1[104] ^ in2[104];
    assign G[9] = in1[103] & in2[103];
    assign P[9] = in1[103] ^ in2[103];
    assign G[10] = in1[102] & in2[102];
    assign P[10] = in1[102] ^ in2[102];
    assign G[11] = in1[101] & in2[101];
    assign P[11] = in1[101] ^ in2[101];
    assign G[12] = in1[100] & in2[100];
    assign P[12] = in1[100] ^ in2[100];
    assign G[13] = in1[99] & in2[99];
    assign P[13] = in1[99] ^ in2[99];
    assign G[14] = in1[98] & in2[98];
    assign P[14] = in1[98] ^ in2[98];
    assign G[15] = in1[97] & in2[97];
    assign P[15] = in1[97] ^ in2[97];
    assign G[16] = in1[96] & in2[96];
    assign P[16] = in1[96] ^ in2[96];
    assign G[17] = in1[95] & in2[95];
    assign P[17] = in1[95] ^ in2[95];
    assign G[18] = in1[94] & in2[94];
    assign P[18] = in1[94] ^ in2[94];
    assign G[19] = in1[93] & in2[93];
    assign P[19] = in1[93] ^ in2[93];
    assign G[20] = in1[92] & in2[92];
    assign P[20] = in1[92] ^ in2[92];
    assign G[21] = in1[91] & in2[91];
    assign P[21] = in1[91] ^ in2[91];
    assign G[22] = in1[90] & in2[90];
    assign P[22] = in1[90] ^ in2[90];
    assign G[23] = in1[89] & in2[89];
    assign P[23] = in1[89] ^ in2[89];
    assign G[24] = in1[88] & in2[88];
    assign P[24] = in1[88] ^ in2[88];
    assign G[25] = in1[87] & in2[87];
    assign P[25] = in1[87] ^ in2[87];
    assign G[26] = in1[86] & in2[86];
    assign P[26] = in1[86] ^ in2[86];
    assign G[27] = in1[85] & in2[85];
    assign P[27] = in1[85] ^ in2[85];
    assign G[28] = in1[84] & in2[84];
    assign P[28] = in1[84] ^ in2[84];
    assign G[29] = in1[83] & in2[83];
    assign P[29] = in1[83] ^ in2[83];
    assign G[30] = in1[82] & in2[82];
    assign P[30] = in1[82] ^ in2[82];
    assign G[31] = in1[81] & in2[81];
    assign P[31] = in1[81] ^ in2[81];
    assign G[32] = in1[80] & in2[80];
    assign P[32] = in1[80] ^ in2[80];
    assign G[33] = in1[79] & in2[79];
    assign P[33] = in1[79] ^ in2[79];
    assign G[34] = in1[78] & in2[78];
    assign P[34] = in1[78] ^ in2[78];
    assign G[35] = in1[77] & in2[77];
    assign P[35] = in1[77] ^ in2[77];
    assign G[36] = in1[76] & in2[76];
    assign P[36] = in1[76] ^ in2[76];
    assign G[37] = in1[75] & in2[75];
    assign P[37] = in1[75] ^ in2[75];
    assign G[38] = in1[74] & in2[74];
    assign P[38] = in1[74] ^ in2[74];
    assign G[39] = in1[73] & in2[73];
    assign P[39] = in1[73] ^ in2[73];
    assign G[40] = in1[72] & in2[72];
    assign P[40] = in1[72] ^ in2[72];
    assign G[41] = in1[71] & in2[71];
    assign P[41] = in1[71] ^ in2[71];
    assign G[42] = in1[70] & in2[70];
    assign P[42] = in1[70] ^ in2[70];
    assign G[43] = in1[69] & in2[69];
    assign P[43] = in1[69] ^ in2[69];
    assign G[44] = in1[68] & in2[68];
    assign P[44] = in1[68] ^ in2[68];
    assign G[45] = in1[67] & in2[67];
    assign P[45] = in1[67] ^ in2[67];
    assign G[46] = in1[66] & in2[66];
    assign P[46] = in1[66] ^ in2[66];
    assign G[47] = in1[65] & in2[65];
    assign P[47] = in1[65] ^ in2[65];
    assign G[48] = in1[64] & in2[64];
    assign P[48] = in1[64] ^ in2[64];
    assign G[49] = in1[63] & in2[63];
    assign P[49] = in1[63] ^ in2[63];
    assign G[50] = in1[62] & in2[62];
    assign P[50] = in1[62] ^ in2[62];
    assign G[51] = in1[61] & in2[61];
    assign P[51] = in1[61] ^ in2[61];
    assign G[52] = in1[60] & in2[60];
    assign P[52] = in1[60] ^ in2[60];
    assign G[53] = in1[59] & in2[59];
    assign P[53] = in1[59] ^ in2[59];
    assign G[54] = in1[58] & in2[58];
    assign P[54] = in1[58] ^ in2[58];
    assign G[55] = in1[57] & in2[57];
    assign P[55] = in1[57] ^ in2[57];
    assign G[56] = in1[56] & in2[56];
    assign P[56] = in1[56] ^ in2[56];
    assign G[57] = in1[55] & in2[55];
    assign P[57] = in1[55] ^ in2[55];
    assign G[58] = in1[54] & in2[54];
    assign P[58] = in1[54] ^ in2[54];
    assign G[59] = in1[53] & in2[53];
    assign P[59] = in1[53] ^ in2[53];
    assign G[60] = in1[52] & in2[52];
    assign P[60] = in1[52] ^ in2[52];
    assign G[61] = in1[51] & in2[51];
    assign P[61] = in1[51] ^ in2[51];
    assign G[62] = in1[50] & in2[50];
    assign P[62] = in1[50] ^ in2[50];
    assign G[63] = in1[49] & in2[49];
    assign P[63] = in1[49] ^ in2[49];
    assign G[64] = in1[48] & in2[48];
    assign P[64] = in1[48] ^ in2[48];
    assign G[65] = in1[47] & in2[47];
    assign P[65] = in1[47] ^ in2[47];
    assign G[66] = in1[46] & in2[46];
    assign P[66] = in1[46] ^ in2[46];
    assign G[67] = in1[45] & in2[45];
    assign P[67] = in1[45] ^ in2[45];
    assign G[68] = in1[44] & in2[44];
    assign P[68] = in1[44] ^ in2[44];
    assign G[69] = in1[43] & in2[43];
    assign P[69] = in1[43] ^ in2[43];
    assign G[70] = in1[42] & in2[42];
    assign P[70] = in1[42] ^ in2[42];
    assign G[71] = in1[41] & in2[41];
    assign P[71] = in1[41] ^ in2[41];
    assign G[72] = in1[40] & in2[40];
    assign P[72] = in1[40] ^ in2[40];
    assign G[73] = in1[39] & in2[39];
    assign P[73] = in1[39] ^ in2[39];
    assign G[74] = in1[38] & in2[38];
    assign P[74] = in1[38] ^ in2[38];
    assign G[75] = in1[37] & in2[37];
    assign P[75] = in1[37] ^ in2[37];
    assign G[76] = in1[36] & in2[36];
    assign P[76] = in1[36] ^ in2[36];
    assign G[77] = in1[35] & in2[35];
    assign P[77] = in1[35] ^ in2[35];
    assign G[78] = in1[34] & in2[34];
    assign P[78] = in1[34] ^ in2[34];
    assign G[79] = in1[33] & in2[33];
    assign P[79] = in1[33] ^ in2[33];
    assign G[80] = in1[32] & in2[32];
    assign P[80] = in1[32] ^ in2[32];
    assign G[81] = in1[31] & in2[31];
    assign P[81] = in1[31] ^ in2[31];
    assign G[82] = in1[30] & in2[30];
    assign P[82] = in1[30] ^ in2[30];
    assign G[83] = in1[29] & in2[29];
    assign P[83] = in1[29] ^ in2[29];
    assign G[84] = in1[28] & in2[28];
    assign P[84] = in1[28] ^ in2[28];
    assign G[85] = in1[27] & in2[27];
    assign P[85] = in1[27] ^ in2[27];
    assign G[86] = in1[26] & in2[26];
    assign P[86] = in1[26] ^ in2[26];
    assign G[87] = in1[25] & in2[25];
    assign P[87] = in1[25] ^ in2[25];
    assign G[88] = in1[24] & in2[24];
    assign P[88] = in1[24] ^ in2[24];
    assign G[89] = in1[23] & in2[23];
    assign P[89] = in1[23] ^ in2[23];
    assign G[90] = in1[22] & in2[22];
    assign P[90] = in1[22] ^ in2[22];
    assign G[91] = in1[21] & in2[21];
    assign P[91] = in1[21] ^ in2[21];
    assign G[92] = in1[20] & in2[20];
    assign P[92] = in1[20] ^ in2[20];
    assign G[93] = in1[19] & in2[19];
    assign P[93] = in1[19] ^ in2[19];
    assign G[94] = in1[18] & in2[18];
    assign P[94] = in1[18] ^ in2[18];
    assign G[95] = in1[17] & in2[17];
    assign P[95] = in1[17] ^ in2[17];
    assign G[96] = in1[16] & in2[16];
    assign P[96] = in1[16] ^ in2[16];
    assign G[97] = in1[15] & in2[15];
    assign P[97] = in1[15] ^ in2[15];
    assign G[98] = in1[14] & in2[14];
    assign P[98] = in1[14] ^ in2[14];
    assign G[99] = in1[13] & in2[13];
    assign P[99] = in1[13] ^ in2[13];
    assign G[100] = in1[12] & in2[12];
    assign P[100] = in1[12] ^ in2[12];
    assign G[101] = in1[11] & in2[11];
    assign P[101] = in1[11] ^ in2[11];
    assign G[102] = in1[10] & in2[10];
    assign P[102] = in1[10] ^ in2[10];
    assign G[103] = in1[9] & in2[9];
    assign P[103] = in1[9] ^ in2[9];
    assign G[104] = in1[8] & in2[8];
    assign P[104] = in1[8] ^ in2[8];
    assign G[105] = in1[7] & in2[7];
    assign P[105] = in1[7] ^ in2[7];
    assign G[106] = in1[6] & in2[6];
    assign P[106] = in1[6] ^ in2[6];
    assign G[107] = in1[5] & in2[5];
    assign P[107] = in1[5] ^ in2[5];
    assign G[108] = in1[4] & in2[4];
    assign P[108] = in1[4] ^ in2[4];
    assign G[109] = in1[3] & in2[3];
    assign P[109] = in1[3] ^ in2[3];
    assign G[110] = in1[2] & in2[2];
    assign P[110] = in1[2] ^ in2[2];
    assign G[111] = in1[1] & in2[1];
    assign P[111] = in1[1] ^ in2[1];
    assign G[112] = in1[0] & in2[0];
    assign P[112] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign cout = G[112] | (P[112] & C[112]);
    assign sum = P ^ C;
endmodule

module CLA_112(output [111:0] sum, output cout, input [111:0] in1, input [111:0] in2);

    wire[111:0] G;
    wire[111:0] C;
    wire[111:0] P;

    assign G[0] = in1[111] & in2[111];
    assign P[0] = in1[111] ^ in2[111];
    assign G[1] = in1[110] & in2[110];
    assign P[1] = in1[110] ^ in2[110];
    assign G[2] = in1[109] & in2[109];
    assign P[2] = in1[109] ^ in2[109];
    assign G[3] = in1[108] & in2[108];
    assign P[3] = in1[108] ^ in2[108];
    assign G[4] = in1[107] & in2[107];
    assign P[4] = in1[107] ^ in2[107];
    assign G[5] = in1[106] & in2[106];
    assign P[5] = in1[106] ^ in2[106];
    assign G[6] = in1[105] & in2[105];
    assign P[6] = in1[105] ^ in2[105];
    assign G[7] = in1[104] & in2[104];
    assign P[7] = in1[104] ^ in2[104];
    assign G[8] = in1[103] & in2[103];
    assign P[8] = in1[103] ^ in2[103];
    assign G[9] = in1[102] & in2[102];
    assign P[9] = in1[102] ^ in2[102];
    assign G[10] = in1[101] & in2[101];
    assign P[10] = in1[101] ^ in2[101];
    assign G[11] = in1[100] & in2[100];
    assign P[11] = in1[100] ^ in2[100];
    assign G[12] = in1[99] & in2[99];
    assign P[12] = in1[99] ^ in2[99];
    assign G[13] = in1[98] & in2[98];
    assign P[13] = in1[98] ^ in2[98];
    assign G[14] = in1[97] & in2[97];
    assign P[14] = in1[97] ^ in2[97];
    assign G[15] = in1[96] & in2[96];
    assign P[15] = in1[96] ^ in2[96];
    assign G[16] = in1[95] & in2[95];
    assign P[16] = in1[95] ^ in2[95];
    assign G[17] = in1[94] & in2[94];
    assign P[17] = in1[94] ^ in2[94];
    assign G[18] = in1[93] & in2[93];
    assign P[18] = in1[93] ^ in2[93];
    assign G[19] = in1[92] & in2[92];
    assign P[19] = in1[92] ^ in2[92];
    assign G[20] = in1[91] & in2[91];
    assign P[20] = in1[91] ^ in2[91];
    assign G[21] = in1[90] & in2[90];
    assign P[21] = in1[90] ^ in2[90];
    assign G[22] = in1[89] & in2[89];
    assign P[22] = in1[89] ^ in2[89];
    assign G[23] = in1[88] & in2[88];
    assign P[23] = in1[88] ^ in2[88];
    assign G[24] = in1[87] & in2[87];
    assign P[24] = in1[87] ^ in2[87];
    assign G[25] = in1[86] & in2[86];
    assign P[25] = in1[86] ^ in2[86];
    assign G[26] = in1[85] & in2[85];
    assign P[26] = in1[85] ^ in2[85];
    assign G[27] = in1[84] & in2[84];
    assign P[27] = in1[84] ^ in2[84];
    assign G[28] = in1[83] & in2[83];
    assign P[28] = in1[83] ^ in2[83];
    assign G[29] = in1[82] & in2[82];
    assign P[29] = in1[82] ^ in2[82];
    assign G[30] = in1[81] & in2[81];
    assign P[30] = in1[81] ^ in2[81];
    assign G[31] = in1[80] & in2[80];
    assign P[31] = in1[80] ^ in2[80];
    assign G[32] = in1[79] & in2[79];
    assign P[32] = in1[79] ^ in2[79];
    assign G[33] = in1[78] & in2[78];
    assign P[33] = in1[78] ^ in2[78];
    assign G[34] = in1[77] & in2[77];
    assign P[34] = in1[77] ^ in2[77];
    assign G[35] = in1[76] & in2[76];
    assign P[35] = in1[76] ^ in2[76];
    assign G[36] = in1[75] & in2[75];
    assign P[36] = in1[75] ^ in2[75];
    assign G[37] = in1[74] & in2[74];
    assign P[37] = in1[74] ^ in2[74];
    assign G[38] = in1[73] & in2[73];
    assign P[38] = in1[73] ^ in2[73];
    assign G[39] = in1[72] & in2[72];
    assign P[39] = in1[72] ^ in2[72];
    assign G[40] = in1[71] & in2[71];
    assign P[40] = in1[71] ^ in2[71];
    assign G[41] = in1[70] & in2[70];
    assign P[41] = in1[70] ^ in2[70];
    assign G[42] = in1[69] & in2[69];
    assign P[42] = in1[69] ^ in2[69];
    assign G[43] = in1[68] & in2[68];
    assign P[43] = in1[68] ^ in2[68];
    assign G[44] = in1[67] & in2[67];
    assign P[44] = in1[67] ^ in2[67];
    assign G[45] = in1[66] & in2[66];
    assign P[45] = in1[66] ^ in2[66];
    assign G[46] = in1[65] & in2[65];
    assign P[46] = in1[65] ^ in2[65];
    assign G[47] = in1[64] & in2[64];
    assign P[47] = in1[64] ^ in2[64];
    assign G[48] = in1[63] & in2[63];
    assign P[48] = in1[63] ^ in2[63];
    assign G[49] = in1[62] & in2[62];
    assign P[49] = in1[62] ^ in2[62];
    assign G[50] = in1[61] & in2[61];
    assign P[50] = in1[61] ^ in2[61];
    assign G[51] = in1[60] & in2[60];
    assign P[51] = in1[60] ^ in2[60];
    assign G[52] = in1[59] & in2[59];
    assign P[52] = in1[59] ^ in2[59];
    assign G[53] = in1[58] & in2[58];
    assign P[53] = in1[58] ^ in2[58];
    assign G[54] = in1[57] & in2[57];
    assign P[54] = in1[57] ^ in2[57];
    assign G[55] = in1[56] & in2[56];
    assign P[55] = in1[56] ^ in2[56];
    assign G[56] = in1[55] & in2[55];
    assign P[56] = in1[55] ^ in2[55];
    assign G[57] = in1[54] & in2[54];
    assign P[57] = in1[54] ^ in2[54];
    assign G[58] = in1[53] & in2[53];
    assign P[58] = in1[53] ^ in2[53];
    assign G[59] = in1[52] & in2[52];
    assign P[59] = in1[52] ^ in2[52];
    assign G[60] = in1[51] & in2[51];
    assign P[60] = in1[51] ^ in2[51];
    assign G[61] = in1[50] & in2[50];
    assign P[61] = in1[50] ^ in2[50];
    assign G[62] = in1[49] & in2[49];
    assign P[62] = in1[49] ^ in2[49];
    assign G[63] = in1[48] & in2[48];
    assign P[63] = in1[48] ^ in2[48];
    assign G[64] = in1[47] & in2[47];
    assign P[64] = in1[47] ^ in2[47];
    assign G[65] = in1[46] & in2[46];
    assign P[65] = in1[46] ^ in2[46];
    assign G[66] = in1[45] & in2[45];
    assign P[66] = in1[45] ^ in2[45];
    assign G[67] = in1[44] & in2[44];
    assign P[67] = in1[44] ^ in2[44];
    assign G[68] = in1[43] & in2[43];
    assign P[68] = in1[43] ^ in2[43];
    assign G[69] = in1[42] & in2[42];
    assign P[69] = in1[42] ^ in2[42];
    assign G[70] = in1[41] & in2[41];
    assign P[70] = in1[41] ^ in2[41];
    assign G[71] = in1[40] & in2[40];
    assign P[71] = in1[40] ^ in2[40];
    assign G[72] = in1[39] & in2[39];
    assign P[72] = in1[39] ^ in2[39];
    assign G[73] = in1[38] & in2[38];
    assign P[73] = in1[38] ^ in2[38];
    assign G[74] = in1[37] & in2[37];
    assign P[74] = in1[37] ^ in2[37];
    assign G[75] = in1[36] & in2[36];
    assign P[75] = in1[36] ^ in2[36];
    assign G[76] = in1[35] & in2[35];
    assign P[76] = in1[35] ^ in2[35];
    assign G[77] = in1[34] & in2[34];
    assign P[77] = in1[34] ^ in2[34];
    assign G[78] = in1[33] & in2[33];
    assign P[78] = in1[33] ^ in2[33];
    assign G[79] = in1[32] & in2[32];
    assign P[79] = in1[32] ^ in2[32];
    assign G[80] = in1[31] & in2[31];
    assign P[80] = in1[31] ^ in2[31];
    assign G[81] = in1[30] & in2[30];
    assign P[81] = in1[30] ^ in2[30];
    assign G[82] = in1[29] & in2[29];
    assign P[82] = in1[29] ^ in2[29];
    assign G[83] = in1[28] & in2[28];
    assign P[83] = in1[28] ^ in2[28];
    assign G[84] = in1[27] & in2[27];
    assign P[84] = in1[27] ^ in2[27];
    assign G[85] = in1[26] & in2[26];
    assign P[85] = in1[26] ^ in2[26];
    assign G[86] = in1[25] & in2[25];
    assign P[86] = in1[25] ^ in2[25];
    assign G[87] = in1[24] & in2[24];
    assign P[87] = in1[24] ^ in2[24];
    assign G[88] = in1[23] & in2[23];
    assign P[88] = in1[23] ^ in2[23];
    assign G[89] = in1[22] & in2[22];
    assign P[89] = in1[22] ^ in2[22];
    assign G[90] = in1[21] & in2[21];
    assign P[90] = in1[21] ^ in2[21];
    assign G[91] = in1[20] & in2[20];
    assign P[91] = in1[20] ^ in2[20];
    assign G[92] = in1[19] & in2[19];
    assign P[92] = in1[19] ^ in2[19];
    assign G[93] = in1[18] & in2[18];
    assign P[93] = in1[18] ^ in2[18];
    assign G[94] = in1[17] & in2[17];
    assign P[94] = in1[17] ^ in2[17];
    assign G[95] = in1[16] & in2[16];
    assign P[95] = in1[16] ^ in2[16];
    assign G[96] = in1[15] & in2[15];
    assign P[96] = in1[15] ^ in2[15];
    assign G[97] = in1[14] & in2[14];
    assign P[97] = in1[14] ^ in2[14];
    assign G[98] = in1[13] & in2[13];
    assign P[98] = in1[13] ^ in2[13];
    assign G[99] = in1[12] & in2[12];
    assign P[99] = in1[12] ^ in2[12];
    assign G[100] = in1[11] & in2[11];
    assign P[100] = in1[11] ^ in2[11];
    assign G[101] = in1[10] & in2[10];
    assign P[101] = in1[10] ^ in2[10];
    assign G[102] = in1[9] & in2[9];
    assign P[102] = in1[9] ^ in2[9];
    assign G[103] = in1[8] & in2[8];
    assign P[103] = in1[8] ^ in2[8];
    assign G[104] = in1[7] & in2[7];
    assign P[104] = in1[7] ^ in2[7];
    assign G[105] = in1[6] & in2[6];
    assign P[105] = in1[6] ^ in2[6];
    assign G[106] = in1[5] & in2[5];
    assign P[106] = in1[5] ^ in2[5];
    assign G[107] = in1[4] & in2[4];
    assign P[107] = in1[4] ^ in2[4];
    assign G[108] = in1[3] & in2[3];
    assign P[108] = in1[3] ^ in2[3];
    assign G[109] = in1[2] & in2[2];
    assign P[109] = in1[2] ^ in2[2];
    assign G[110] = in1[1] & in2[1];
    assign P[110] = in1[1] ^ in2[1];
    assign G[111] = in1[0] & in2[0];
    assign P[111] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign cout = G[111] | (P[111] & C[111]);
    assign sum = P ^ C;
endmodule

module CLA_111(output [110:0] sum, output cout, input [110:0] in1, input [110:0] in2);

    wire[110:0] G;
    wire[110:0] C;
    wire[110:0] P;

    assign G[0] = in1[110] & in2[110];
    assign P[0] = in1[110] ^ in2[110];
    assign G[1] = in1[109] & in2[109];
    assign P[1] = in1[109] ^ in2[109];
    assign G[2] = in1[108] & in2[108];
    assign P[2] = in1[108] ^ in2[108];
    assign G[3] = in1[107] & in2[107];
    assign P[3] = in1[107] ^ in2[107];
    assign G[4] = in1[106] & in2[106];
    assign P[4] = in1[106] ^ in2[106];
    assign G[5] = in1[105] & in2[105];
    assign P[5] = in1[105] ^ in2[105];
    assign G[6] = in1[104] & in2[104];
    assign P[6] = in1[104] ^ in2[104];
    assign G[7] = in1[103] & in2[103];
    assign P[7] = in1[103] ^ in2[103];
    assign G[8] = in1[102] & in2[102];
    assign P[8] = in1[102] ^ in2[102];
    assign G[9] = in1[101] & in2[101];
    assign P[9] = in1[101] ^ in2[101];
    assign G[10] = in1[100] & in2[100];
    assign P[10] = in1[100] ^ in2[100];
    assign G[11] = in1[99] & in2[99];
    assign P[11] = in1[99] ^ in2[99];
    assign G[12] = in1[98] & in2[98];
    assign P[12] = in1[98] ^ in2[98];
    assign G[13] = in1[97] & in2[97];
    assign P[13] = in1[97] ^ in2[97];
    assign G[14] = in1[96] & in2[96];
    assign P[14] = in1[96] ^ in2[96];
    assign G[15] = in1[95] & in2[95];
    assign P[15] = in1[95] ^ in2[95];
    assign G[16] = in1[94] & in2[94];
    assign P[16] = in1[94] ^ in2[94];
    assign G[17] = in1[93] & in2[93];
    assign P[17] = in1[93] ^ in2[93];
    assign G[18] = in1[92] & in2[92];
    assign P[18] = in1[92] ^ in2[92];
    assign G[19] = in1[91] & in2[91];
    assign P[19] = in1[91] ^ in2[91];
    assign G[20] = in1[90] & in2[90];
    assign P[20] = in1[90] ^ in2[90];
    assign G[21] = in1[89] & in2[89];
    assign P[21] = in1[89] ^ in2[89];
    assign G[22] = in1[88] & in2[88];
    assign P[22] = in1[88] ^ in2[88];
    assign G[23] = in1[87] & in2[87];
    assign P[23] = in1[87] ^ in2[87];
    assign G[24] = in1[86] & in2[86];
    assign P[24] = in1[86] ^ in2[86];
    assign G[25] = in1[85] & in2[85];
    assign P[25] = in1[85] ^ in2[85];
    assign G[26] = in1[84] & in2[84];
    assign P[26] = in1[84] ^ in2[84];
    assign G[27] = in1[83] & in2[83];
    assign P[27] = in1[83] ^ in2[83];
    assign G[28] = in1[82] & in2[82];
    assign P[28] = in1[82] ^ in2[82];
    assign G[29] = in1[81] & in2[81];
    assign P[29] = in1[81] ^ in2[81];
    assign G[30] = in1[80] & in2[80];
    assign P[30] = in1[80] ^ in2[80];
    assign G[31] = in1[79] & in2[79];
    assign P[31] = in1[79] ^ in2[79];
    assign G[32] = in1[78] & in2[78];
    assign P[32] = in1[78] ^ in2[78];
    assign G[33] = in1[77] & in2[77];
    assign P[33] = in1[77] ^ in2[77];
    assign G[34] = in1[76] & in2[76];
    assign P[34] = in1[76] ^ in2[76];
    assign G[35] = in1[75] & in2[75];
    assign P[35] = in1[75] ^ in2[75];
    assign G[36] = in1[74] & in2[74];
    assign P[36] = in1[74] ^ in2[74];
    assign G[37] = in1[73] & in2[73];
    assign P[37] = in1[73] ^ in2[73];
    assign G[38] = in1[72] & in2[72];
    assign P[38] = in1[72] ^ in2[72];
    assign G[39] = in1[71] & in2[71];
    assign P[39] = in1[71] ^ in2[71];
    assign G[40] = in1[70] & in2[70];
    assign P[40] = in1[70] ^ in2[70];
    assign G[41] = in1[69] & in2[69];
    assign P[41] = in1[69] ^ in2[69];
    assign G[42] = in1[68] & in2[68];
    assign P[42] = in1[68] ^ in2[68];
    assign G[43] = in1[67] & in2[67];
    assign P[43] = in1[67] ^ in2[67];
    assign G[44] = in1[66] & in2[66];
    assign P[44] = in1[66] ^ in2[66];
    assign G[45] = in1[65] & in2[65];
    assign P[45] = in1[65] ^ in2[65];
    assign G[46] = in1[64] & in2[64];
    assign P[46] = in1[64] ^ in2[64];
    assign G[47] = in1[63] & in2[63];
    assign P[47] = in1[63] ^ in2[63];
    assign G[48] = in1[62] & in2[62];
    assign P[48] = in1[62] ^ in2[62];
    assign G[49] = in1[61] & in2[61];
    assign P[49] = in1[61] ^ in2[61];
    assign G[50] = in1[60] & in2[60];
    assign P[50] = in1[60] ^ in2[60];
    assign G[51] = in1[59] & in2[59];
    assign P[51] = in1[59] ^ in2[59];
    assign G[52] = in1[58] & in2[58];
    assign P[52] = in1[58] ^ in2[58];
    assign G[53] = in1[57] & in2[57];
    assign P[53] = in1[57] ^ in2[57];
    assign G[54] = in1[56] & in2[56];
    assign P[54] = in1[56] ^ in2[56];
    assign G[55] = in1[55] & in2[55];
    assign P[55] = in1[55] ^ in2[55];
    assign G[56] = in1[54] & in2[54];
    assign P[56] = in1[54] ^ in2[54];
    assign G[57] = in1[53] & in2[53];
    assign P[57] = in1[53] ^ in2[53];
    assign G[58] = in1[52] & in2[52];
    assign P[58] = in1[52] ^ in2[52];
    assign G[59] = in1[51] & in2[51];
    assign P[59] = in1[51] ^ in2[51];
    assign G[60] = in1[50] & in2[50];
    assign P[60] = in1[50] ^ in2[50];
    assign G[61] = in1[49] & in2[49];
    assign P[61] = in1[49] ^ in2[49];
    assign G[62] = in1[48] & in2[48];
    assign P[62] = in1[48] ^ in2[48];
    assign G[63] = in1[47] & in2[47];
    assign P[63] = in1[47] ^ in2[47];
    assign G[64] = in1[46] & in2[46];
    assign P[64] = in1[46] ^ in2[46];
    assign G[65] = in1[45] & in2[45];
    assign P[65] = in1[45] ^ in2[45];
    assign G[66] = in1[44] & in2[44];
    assign P[66] = in1[44] ^ in2[44];
    assign G[67] = in1[43] & in2[43];
    assign P[67] = in1[43] ^ in2[43];
    assign G[68] = in1[42] & in2[42];
    assign P[68] = in1[42] ^ in2[42];
    assign G[69] = in1[41] & in2[41];
    assign P[69] = in1[41] ^ in2[41];
    assign G[70] = in1[40] & in2[40];
    assign P[70] = in1[40] ^ in2[40];
    assign G[71] = in1[39] & in2[39];
    assign P[71] = in1[39] ^ in2[39];
    assign G[72] = in1[38] & in2[38];
    assign P[72] = in1[38] ^ in2[38];
    assign G[73] = in1[37] & in2[37];
    assign P[73] = in1[37] ^ in2[37];
    assign G[74] = in1[36] & in2[36];
    assign P[74] = in1[36] ^ in2[36];
    assign G[75] = in1[35] & in2[35];
    assign P[75] = in1[35] ^ in2[35];
    assign G[76] = in1[34] & in2[34];
    assign P[76] = in1[34] ^ in2[34];
    assign G[77] = in1[33] & in2[33];
    assign P[77] = in1[33] ^ in2[33];
    assign G[78] = in1[32] & in2[32];
    assign P[78] = in1[32] ^ in2[32];
    assign G[79] = in1[31] & in2[31];
    assign P[79] = in1[31] ^ in2[31];
    assign G[80] = in1[30] & in2[30];
    assign P[80] = in1[30] ^ in2[30];
    assign G[81] = in1[29] & in2[29];
    assign P[81] = in1[29] ^ in2[29];
    assign G[82] = in1[28] & in2[28];
    assign P[82] = in1[28] ^ in2[28];
    assign G[83] = in1[27] & in2[27];
    assign P[83] = in1[27] ^ in2[27];
    assign G[84] = in1[26] & in2[26];
    assign P[84] = in1[26] ^ in2[26];
    assign G[85] = in1[25] & in2[25];
    assign P[85] = in1[25] ^ in2[25];
    assign G[86] = in1[24] & in2[24];
    assign P[86] = in1[24] ^ in2[24];
    assign G[87] = in1[23] & in2[23];
    assign P[87] = in1[23] ^ in2[23];
    assign G[88] = in1[22] & in2[22];
    assign P[88] = in1[22] ^ in2[22];
    assign G[89] = in1[21] & in2[21];
    assign P[89] = in1[21] ^ in2[21];
    assign G[90] = in1[20] & in2[20];
    assign P[90] = in1[20] ^ in2[20];
    assign G[91] = in1[19] & in2[19];
    assign P[91] = in1[19] ^ in2[19];
    assign G[92] = in1[18] & in2[18];
    assign P[92] = in1[18] ^ in2[18];
    assign G[93] = in1[17] & in2[17];
    assign P[93] = in1[17] ^ in2[17];
    assign G[94] = in1[16] & in2[16];
    assign P[94] = in1[16] ^ in2[16];
    assign G[95] = in1[15] & in2[15];
    assign P[95] = in1[15] ^ in2[15];
    assign G[96] = in1[14] & in2[14];
    assign P[96] = in1[14] ^ in2[14];
    assign G[97] = in1[13] & in2[13];
    assign P[97] = in1[13] ^ in2[13];
    assign G[98] = in1[12] & in2[12];
    assign P[98] = in1[12] ^ in2[12];
    assign G[99] = in1[11] & in2[11];
    assign P[99] = in1[11] ^ in2[11];
    assign G[100] = in1[10] & in2[10];
    assign P[100] = in1[10] ^ in2[10];
    assign G[101] = in1[9] & in2[9];
    assign P[101] = in1[9] ^ in2[9];
    assign G[102] = in1[8] & in2[8];
    assign P[102] = in1[8] ^ in2[8];
    assign G[103] = in1[7] & in2[7];
    assign P[103] = in1[7] ^ in2[7];
    assign G[104] = in1[6] & in2[6];
    assign P[104] = in1[6] ^ in2[6];
    assign G[105] = in1[5] & in2[5];
    assign P[105] = in1[5] ^ in2[5];
    assign G[106] = in1[4] & in2[4];
    assign P[106] = in1[4] ^ in2[4];
    assign G[107] = in1[3] & in2[3];
    assign P[107] = in1[3] ^ in2[3];
    assign G[108] = in1[2] & in2[2];
    assign P[108] = in1[2] ^ in2[2];
    assign G[109] = in1[1] & in2[1];
    assign P[109] = in1[1] ^ in2[1];
    assign G[110] = in1[0] & in2[0];
    assign P[110] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign cout = G[110] | (P[110] & C[110]);
    assign sum = P ^ C;
endmodule

module CLA_110(output [109:0] sum, output cout, input [109:0] in1, input [109:0] in2);

    wire[109:0] G;
    wire[109:0] C;
    wire[109:0] P;

    assign G[0] = in1[109] & in2[109];
    assign P[0] = in1[109] ^ in2[109];
    assign G[1] = in1[108] & in2[108];
    assign P[1] = in1[108] ^ in2[108];
    assign G[2] = in1[107] & in2[107];
    assign P[2] = in1[107] ^ in2[107];
    assign G[3] = in1[106] & in2[106];
    assign P[3] = in1[106] ^ in2[106];
    assign G[4] = in1[105] & in2[105];
    assign P[4] = in1[105] ^ in2[105];
    assign G[5] = in1[104] & in2[104];
    assign P[5] = in1[104] ^ in2[104];
    assign G[6] = in1[103] & in2[103];
    assign P[6] = in1[103] ^ in2[103];
    assign G[7] = in1[102] & in2[102];
    assign P[7] = in1[102] ^ in2[102];
    assign G[8] = in1[101] & in2[101];
    assign P[8] = in1[101] ^ in2[101];
    assign G[9] = in1[100] & in2[100];
    assign P[9] = in1[100] ^ in2[100];
    assign G[10] = in1[99] & in2[99];
    assign P[10] = in1[99] ^ in2[99];
    assign G[11] = in1[98] & in2[98];
    assign P[11] = in1[98] ^ in2[98];
    assign G[12] = in1[97] & in2[97];
    assign P[12] = in1[97] ^ in2[97];
    assign G[13] = in1[96] & in2[96];
    assign P[13] = in1[96] ^ in2[96];
    assign G[14] = in1[95] & in2[95];
    assign P[14] = in1[95] ^ in2[95];
    assign G[15] = in1[94] & in2[94];
    assign P[15] = in1[94] ^ in2[94];
    assign G[16] = in1[93] & in2[93];
    assign P[16] = in1[93] ^ in2[93];
    assign G[17] = in1[92] & in2[92];
    assign P[17] = in1[92] ^ in2[92];
    assign G[18] = in1[91] & in2[91];
    assign P[18] = in1[91] ^ in2[91];
    assign G[19] = in1[90] & in2[90];
    assign P[19] = in1[90] ^ in2[90];
    assign G[20] = in1[89] & in2[89];
    assign P[20] = in1[89] ^ in2[89];
    assign G[21] = in1[88] & in2[88];
    assign P[21] = in1[88] ^ in2[88];
    assign G[22] = in1[87] & in2[87];
    assign P[22] = in1[87] ^ in2[87];
    assign G[23] = in1[86] & in2[86];
    assign P[23] = in1[86] ^ in2[86];
    assign G[24] = in1[85] & in2[85];
    assign P[24] = in1[85] ^ in2[85];
    assign G[25] = in1[84] & in2[84];
    assign P[25] = in1[84] ^ in2[84];
    assign G[26] = in1[83] & in2[83];
    assign P[26] = in1[83] ^ in2[83];
    assign G[27] = in1[82] & in2[82];
    assign P[27] = in1[82] ^ in2[82];
    assign G[28] = in1[81] & in2[81];
    assign P[28] = in1[81] ^ in2[81];
    assign G[29] = in1[80] & in2[80];
    assign P[29] = in1[80] ^ in2[80];
    assign G[30] = in1[79] & in2[79];
    assign P[30] = in1[79] ^ in2[79];
    assign G[31] = in1[78] & in2[78];
    assign P[31] = in1[78] ^ in2[78];
    assign G[32] = in1[77] & in2[77];
    assign P[32] = in1[77] ^ in2[77];
    assign G[33] = in1[76] & in2[76];
    assign P[33] = in1[76] ^ in2[76];
    assign G[34] = in1[75] & in2[75];
    assign P[34] = in1[75] ^ in2[75];
    assign G[35] = in1[74] & in2[74];
    assign P[35] = in1[74] ^ in2[74];
    assign G[36] = in1[73] & in2[73];
    assign P[36] = in1[73] ^ in2[73];
    assign G[37] = in1[72] & in2[72];
    assign P[37] = in1[72] ^ in2[72];
    assign G[38] = in1[71] & in2[71];
    assign P[38] = in1[71] ^ in2[71];
    assign G[39] = in1[70] & in2[70];
    assign P[39] = in1[70] ^ in2[70];
    assign G[40] = in1[69] & in2[69];
    assign P[40] = in1[69] ^ in2[69];
    assign G[41] = in1[68] & in2[68];
    assign P[41] = in1[68] ^ in2[68];
    assign G[42] = in1[67] & in2[67];
    assign P[42] = in1[67] ^ in2[67];
    assign G[43] = in1[66] & in2[66];
    assign P[43] = in1[66] ^ in2[66];
    assign G[44] = in1[65] & in2[65];
    assign P[44] = in1[65] ^ in2[65];
    assign G[45] = in1[64] & in2[64];
    assign P[45] = in1[64] ^ in2[64];
    assign G[46] = in1[63] & in2[63];
    assign P[46] = in1[63] ^ in2[63];
    assign G[47] = in1[62] & in2[62];
    assign P[47] = in1[62] ^ in2[62];
    assign G[48] = in1[61] & in2[61];
    assign P[48] = in1[61] ^ in2[61];
    assign G[49] = in1[60] & in2[60];
    assign P[49] = in1[60] ^ in2[60];
    assign G[50] = in1[59] & in2[59];
    assign P[50] = in1[59] ^ in2[59];
    assign G[51] = in1[58] & in2[58];
    assign P[51] = in1[58] ^ in2[58];
    assign G[52] = in1[57] & in2[57];
    assign P[52] = in1[57] ^ in2[57];
    assign G[53] = in1[56] & in2[56];
    assign P[53] = in1[56] ^ in2[56];
    assign G[54] = in1[55] & in2[55];
    assign P[54] = in1[55] ^ in2[55];
    assign G[55] = in1[54] & in2[54];
    assign P[55] = in1[54] ^ in2[54];
    assign G[56] = in1[53] & in2[53];
    assign P[56] = in1[53] ^ in2[53];
    assign G[57] = in1[52] & in2[52];
    assign P[57] = in1[52] ^ in2[52];
    assign G[58] = in1[51] & in2[51];
    assign P[58] = in1[51] ^ in2[51];
    assign G[59] = in1[50] & in2[50];
    assign P[59] = in1[50] ^ in2[50];
    assign G[60] = in1[49] & in2[49];
    assign P[60] = in1[49] ^ in2[49];
    assign G[61] = in1[48] & in2[48];
    assign P[61] = in1[48] ^ in2[48];
    assign G[62] = in1[47] & in2[47];
    assign P[62] = in1[47] ^ in2[47];
    assign G[63] = in1[46] & in2[46];
    assign P[63] = in1[46] ^ in2[46];
    assign G[64] = in1[45] & in2[45];
    assign P[64] = in1[45] ^ in2[45];
    assign G[65] = in1[44] & in2[44];
    assign P[65] = in1[44] ^ in2[44];
    assign G[66] = in1[43] & in2[43];
    assign P[66] = in1[43] ^ in2[43];
    assign G[67] = in1[42] & in2[42];
    assign P[67] = in1[42] ^ in2[42];
    assign G[68] = in1[41] & in2[41];
    assign P[68] = in1[41] ^ in2[41];
    assign G[69] = in1[40] & in2[40];
    assign P[69] = in1[40] ^ in2[40];
    assign G[70] = in1[39] & in2[39];
    assign P[70] = in1[39] ^ in2[39];
    assign G[71] = in1[38] & in2[38];
    assign P[71] = in1[38] ^ in2[38];
    assign G[72] = in1[37] & in2[37];
    assign P[72] = in1[37] ^ in2[37];
    assign G[73] = in1[36] & in2[36];
    assign P[73] = in1[36] ^ in2[36];
    assign G[74] = in1[35] & in2[35];
    assign P[74] = in1[35] ^ in2[35];
    assign G[75] = in1[34] & in2[34];
    assign P[75] = in1[34] ^ in2[34];
    assign G[76] = in1[33] & in2[33];
    assign P[76] = in1[33] ^ in2[33];
    assign G[77] = in1[32] & in2[32];
    assign P[77] = in1[32] ^ in2[32];
    assign G[78] = in1[31] & in2[31];
    assign P[78] = in1[31] ^ in2[31];
    assign G[79] = in1[30] & in2[30];
    assign P[79] = in1[30] ^ in2[30];
    assign G[80] = in1[29] & in2[29];
    assign P[80] = in1[29] ^ in2[29];
    assign G[81] = in1[28] & in2[28];
    assign P[81] = in1[28] ^ in2[28];
    assign G[82] = in1[27] & in2[27];
    assign P[82] = in1[27] ^ in2[27];
    assign G[83] = in1[26] & in2[26];
    assign P[83] = in1[26] ^ in2[26];
    assign G[84] = in1[25] & in2[25];
    assign P[84] = in1[25] ^ in2[25];
    assign G[85] = in1[24] & in2[24];
    assign P[85] = in1[24] ^ in2[24];
    assign G[86] = in1[23] & in2[23];
    assign P[86] = in1[23] ^ in2[23];
    assign G[87] = in1[22] & in2[22];
    assign P[87] = in1[22] ^ in2[22];
    assign G[88] = in1[21] & in2[21];
    assign P[88] = in1[21] ^ in2[21];
    assign G[89] = in1[20] & in2[20];
    assign P[89] = in1[20] ^ in2[20];
    assign G[90] = in1[19] & in2[19];
    assign P[90] = in1[19] ^ in2[19];
    assign G[91] = in1[18] & in2[18];
    assign P[91] = in1[18] ^ in2[18];
    assign G[92] = in1[17] & in2[17];
    assign P[92] = in1[17] ^ in2[17];
    assign G[93] = in1[16] & in2[16];
    assign P[93] = in1[16] ^ in2[16];
    assign G[94] = in1[15] & in2[15];
    assign P[94] = in1[15] ^ in2[15];
    assign G[95] = in1[14] & in2[14];
    assign P[95] = in1[14] ^ in2[14];
    assign G[96] = in1[13] & in2[13];
    assign P[96] = in1[13] ^ in2[13];
    assign G[97] = in1[12] & in2[12];
    assign P[97] = in1[12] ^ in2[12];
    assign G[98] = in1[11] & in2[11];
    assign P[98] = in1[11] ^ in2[11];
    assign G[99] = in1[10] & in2[10];
    assign P[99] = in1[10] ^ in2[10];
    assign G[100] = in1[9] & in2[9];
    assign P[100] = in1[9] ^ in2[9];
    assign G[101] = in1[8] & in2[8];
    assign P[101] = in1[8] ^ in2[8];
    assign G[102] = in1[7] & in2[7];
    assign P[102] = in1[7] ^ in2[7];
    assign G[103] = in1[6] & in2[6];
    assign P[103] = in1[6] ^ in2[6];
    assign G[104] = in1[5] & in2[5];
    assign P[104] = in1[5] ^ in2[5];
    assign G[105] = in1[4] & in2[4];
    assign P[105] = in1[4] ^ in2[4];
    assign G[106] = in1[3] & in2[3];
    assign P[106] = in1[3] ^ in2[3];
    assign G[107] = in1[2] & in2[2];
    assign P[107] = in1[2] ^ in2[2];
    assign G[108] = in1[1] & in2[1];
    assign P[108] = in1[1] ^ in2[1];
    assign G[109] = in1[0] & in2[0];
    assign P[109] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign cout = G[109] | (P[109] & C[109]);
    assign sum = P ^ C;
endmodule

module CLA_109(output [108:0] sum, output cout, input [108:0] in1, input [108:0] in2);

    wire[108:0] G;
    wire[108:0] C;
    wire[108:0] P;

    assign G[0] = in1[108] & in2[108];
    assign P[0] = in1[108] ^ in2[108];
    assign G[1] = in1[107] & in2[107];
    assign P[1] = in1[107] ^ in2[107];
    assign G[2] = in1[106] & in2[106];
    assign P[2] = in1[106] ^ in2[106];
    assign G[3] = in1[105] & in2[105];
    assign P[3] = in1[105] ^ in2[105];
    assign G[4] = in1[104] & in2[104];
    assign P[4] = in1[104] ^ in2[104];
    assign G[5] = in1[103] & in2[103];
    assign P[5] = in1[103] ^ in2[103];
    assign G[6] = in1[102] & in2[102];
    assign P[6] = in1[102] ^ in2[102];
    assign G[7] = in1[101] & in2[101];
    assign P[7] = in1[101] ^ in2[101];
    assign G[8] = in1[100] & in2[100];
    assign P[8] = in1[100] ^ in2[100];
    assign G[9] = in1[99] & in2[99];
    assign P[9] = in1[99] ^ in2[99];
    assign G[10] = in1[98] & in2[98];
    assign P[10] = in1[98] ^ in2[98];
    assign G[11] = in1[97] & in2[97];
    assign P[11] = in1[97] ^ in2[97];
    assign G[12] = in1[96] & in2[96];
    assign P[12] = in1[96] ^ in2[96];
    assign G[13] = in1[95] & in2[95];
    assign P[13] = in1[95] ^ in2[95];
    assign G[14] = in1[94] & in2[94];
    assign P[14] = in1[94] ^ in2[94];
    assign G[15] = in1[93] & in2[93];
    assign P[15] = in1[93] ^ in2[93];
    assign G[16] = in1[92] & in2[92];
    assign P[16] = in1[92] ^ in2[92];
    assign G[17] = in1[91] & in2[91];
    assign P[17] = in1[91] ^ in2[91];
    assign G[18] = in1[90] & in2[90];
    assign P[18] = in1[90] ^ in2[90];
    assign G[19] = in1[89] & in2[89];
    assign P[19] = in1[89] ^ in2[89];
    assign G[20] = in1[88] & in2[88];
    assign P[20] = in1[88] ^ in2[88];
    assign G[21] = in1[87] & in2[87];
    assign P[21] = in1[87] ^ in2[87];
    assign G[22] = in1[86] & in2[86];
    assign P[22] = in1[86] ^ in2[86];
    assign G[23] = in1[85] & in2[85];
    assign P[23] = in1[85] ^ in2[85];
    assign G[24] = in1[84] & in2[84];
    assign P[24] = in1[84] ^ in2[84];
    assign G[25] = in1[83] & in2[83];
    assign P[25] = in1[83] ^ in2[83];
    assign G[26] = in1[82] & in2[82];
    assign P[26] = in1[82] ^ in2[82];
    assign G[27] = in1[81] & in2[81];
    assign P[27] = in1[81] ^ in2[81];
    assign G[28] = in1[80] & in2[80];
    assign P[28] = in1[80] ^ in2[80];
    assign G[29] = in1[79] & in2[79];
    assign P[29] = in1[79] ^ in2[79];
    assign G[30] = in1[78] & in2[78];
    assign P[30] = in1[78] ^ in2[78];
    assign G[31] = in1[77] & in2[77];
    assign P[31] = in1[77] ^ in2[77];
    assign G[32] = in1[76] & in2[76];
    assign P[32] = in1[76] ^ in2[76];
    assign G[33] = in1[75] & in2[75];
    assign P[33] = in1[75] ^ in2[75];
    assign G[34] = in1[74] & in2[74];
    assign P[34] = in1[74] ^ in2[74];
    assign G[35] = in1[73] & in2[73];
    assign P[35] = in1[73] ^ in2[73];
    assign G[36] = in1[72] & in2[72];
    assign P[36] = in1[72] ^ in2[72];
    assign G[37] = in1[71] & in2[71];
    assign P[37] = in1[71] ^ in2[71];
    assign G[38] = in1[70] & in2[70];
    assign P[38] = in1[70] ^ in2[70];
    assign G[39] = in1[69] & in2[69];
    assign P[39] = in1[69] ^ in2[69];
    assign G[40] = in1[68] & in2[68];
    assign P[40] = in1[68] ^ in2[68];
    assign G[41] = in1[67] & in2[67];
    assign P[41] = in1[67] ^ in2[67];
    assign G[42] = in1[66] & in2[66];
    assign P[42] = in1[66] ^ in2[66];
    assign G[43] = in1[65] & in2[65];
    assign P[43] = in1[65] ^ in2[65];
    assign G[44] = in1[64] & in2[64];
    assign P[44] = in1[64] ^ in2[64];
    assign G[45] = in1[63] & in2[63];
    assign P[45] = in1[63] ^ in2[63];
    assign G[46] = in1[62] & in2[62];
    assign P[46] = in1[62] ^ in2[62];
    assign G[47] = in1[61] & in2[61];
    assign P[47] = in1[61] ^ in2[61];
    assign G[48] = in1[60] & in2[60];
    assign P[48] = in1[60] ^ in2[60];
    assign G[49] = in1[59] & in2[59];
    assign P[49] = in1[59] ^ in2[59];
    assign G[50] = in1[58] & in2[58];
    assign P[50] = in1[58] ^ in2[58];
    assign G[51] = in1[57] & in2[57];
    assign P[51] = in1[57] ^ in2[57];
    assign G[52] = in1[56] & in2[56];
    assign P[52] = in1[56] ^ in2[56];
    assign G[53] = in1[55] & in2[55];
    assign P[53] = in1[55] ^ in2[55];
    assign G[54] = in1[54] & in2[54];
    assign P[54] = in1[54] ^ in2[54];
    assign G[55] = in1[53] & in2[53];
    assign P[55] = in1[53] ^ in2[53];
    assign G[56] = in1[52] & in2[52];
    assign P[56] = in1[52] ^ in2[52];
    assign G[57] = in1[51] & in2[51];
    assign P[57] = in1[51] ^ in2[51];
    assign G[58] = in1[50] & in2[50];
    assign P[58] = in1[50] ^ in2[50];
    assign G[59] = in1[49] & in2[49];
    assign P[59] = in1[49] ^ in2[49];
    assign G[60] = in1[48] & in2[48];
    assign P[60] = in1[48] ^ in2[48];
    assign G[61] = in1[47] & in2[47];
    assign P[61] = in1[47] ^ in2[47];
    assign G[62] = in1[46] & in2[46];
    assign P[62] = in1[46] ^ in2[46];
    assign G[63] = in1[45] & in2[45];
    assign P[63] = in1[45] ^ in2[45];
    assign G[64] = in1[44] & in2[44];
    assign P[64] = in1[44] ^ in2[44];
    assign G[65] = in1[43] & in2[43];
    assign P[65] = in1[43] ^ in2[43];
    assign G[66] = in1[42] & in2[42];
    assign P[66] = in1[42] ^ in2[42];
    assign G[67] = in1[41] & in2[41];
    assign P[67] = in1[41] ^ in2[41];
    assign G[68] = in1[40] & in2[40];
    assign P[68] = in1[40] ^ in2[40];
    assign G[69] = in1[39] & in2[39];
    assign P[69] = in1[39] ^ in2[39];
    assign G[70] = in1[38] & in2[38];
    assign P[70] = in1[38] ^ in2[38];
    assign G[71] = in1[37] & in2[37];
    assign P[71] = in1[37] ^ in2[37];
    assign G[72] = in1[36] & in2[36];
    assign P[72] = in1[36] ^ in2[36];
    assign G[73] = in1[35] & in2[35];
    assign P[73] = in1[35] ^ in2[35];
    assign G[74] = in1[34] & in2[34];
    assign P[74] = in1[34] ^ in2[34];
    assign G[75] = in1[33] & in2[33];
    assign P[75] = in1[33] ^ in2[33];
    assign G[76] = in1[32] & in2[32];
    assign P[76] = in1[32] ^ in2[32];
    assign G[77] = in1[31] & in2[31];
    assign P[77] = in1[31] ^ in2[31];
    assign G[78] = in1[30] & in2[30];
    assign P[78] = in1[30] ^ in2[30];
    assign G[79] = in1[29] & in2[29];
    assign P[79] = in1[29] ^ in2[29];
    assign G[80] = in1[28] & in2[28];
    assign P[80] = in1[28] ^ in2[28];
    assign G[81] = in1[27] & in2[27];
    assign P[81] = in1[27] ^ in2[27];
    assign G[82] = in1[26] & in2[26];
    assign P[82] = in1[26] ^ in2[26];
    assign G[83] = in1[25] & in2[25];
    assign P[83] = in1[25] ^ in2[25];
    assign G[84] = in1[24] & in2[24];
    assign P[84] = in1[24] ^ in2[24];
    assign G[85] = in1[23] & in2[23];
    assign P[85] = in1[23] ^ in2[23];
    assign G[86] = in1[22] & in2[22];
    assign P[86] = in1[22] ^ in2[22];
    assign G[87] = in1[21] & in2[21];
    assign P[87] = in1[21] ^ in2[21];
    assign G[88] = in1[20] & in2[20];
    assign P[88] = in1[20] ^ in2[20];
    assign G[89] = in1[19] & in2[19];
    assign P[89] = in1[19] ^ in2[19];
    assign G[90] = in1[18] & in2[18];
    assign P[90] = in1[18] ^ in2[18];
    assign G[91] = in1[17] & in2[17];
    assign P[91] = in1[17] ^ in2[17];
    assign G[92] = in1[16] & in2[16];
    assign P[92] = in1[16] ^ in2[16];
    assign G[93] = in1[15] & in2[15];
    assign P[93] = in1[15] ^ in2[15];
    assign G[94] = in1[14] & in2[14];
    assign P[94] = in1[14] ^ in2[14];
    assign G[95] = in1[13] & in2[13];
    assign P[95] = in1[13] ^ in2[13];
    assign G[96] = in1[12] & in2[12];
    assign P[96] = in1[12] ^ in2[12];
    assign G[97] = in1[11] & in2[11];
    assign P[97] = in1[11] ^ in2[11];
    assign G[98] = in1[10] & in2[10];
    assign P[98] = in1[10] ^ in2[10];
    assign G[99] = in1[9] & in2[9];
    assign P[99] = in1[9] ^ in2[9];
    assign G[100] = in1[8] & in2[8];
    assign P[100] = in1[8] ^ in2[8];
    assign G[101] = in1[7] & in2[7];
    assign P[101] = in1[7] ^ in2[7];
    assign G[102] = in1[6] & in2[6];
    assign P[102] = in1[6] ^ in2[6];
    assign G[103] = in1[5] & in2[5];
    assign P[103] = in1[5] ^ in2[5];
    assign G[104] = in1[4] & in2[4];
    assign P[104] = in1[4] ^ in2[4];
    assign G[105] = in1[3] & in2[3];
    assign P[105] = in1[3] ^ in2[3];
    assign G[106] = in1[2] & in2[2];
    assign P[106] = in1[2] ^ in2[2];
    assign G[107] = in1[1] & in2[1];
    assign P[107] = in1[1] ^ in2[1];
    assign G[108] = in1[0] & in2[0];
    assign P[108] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign cout = G[108] | (P[108] & C[108]);
    assign sum = P ^ C;
endmodule

module CLA_108(output [107:0] sum, output cout, input [107:0] in1, input [107:0] in2);

    wire[107:0] G;
    wire[107:0] C;
    wire[107:0] P;

    assign G[0] = in1[107] & in2[107];
    assign P[0] = in1[107] ^ in2[107];
    assign G[1] = in1[106] & in2[106];
    assign P[1] = in1[106] ^ in2[106];
    assign G[2] = in1[105] & in2[105];
    assign P[2] = in1[105] ^ in2[105];
    assign G[3] = in1[104] & in2[104];
    assign P[3] = in1[104] ^ in2[104];
    assign G[4] = in1[103] & in2[103];
    assign P[4] = in1[103] ^ in2[103];
    assign G[5] = in1[102] & in2[102];
    assign P[5] = in1[102] ^ in2[102];
    assign G[6] = in1[101] & in2[101];
    assign P[6] = in1[101] ^ in2[101];
    assign G[7] = in1[100] & in2[100];
    assign P[7] = in1[100] ^ in2[100];
    assign G[8] = in1[99] & in2[99];
    assign P[8] = in1[99] ^ in2[99];
    assign G[9] = in1[98] & in2[98];
    assign P[9] = in1[98] ^ in2[98];
    assign G[10] = in1[97] & in2[97];
    assign P[10] = in1[97] ^ in2[97];
    assign G[11] = in1[96] & in2[96];
    assign P[11] = in1[96] ^ in2[96];
    assign G[12] = in1[95] & in2[95];
    assign P[12] = in1[95] ^ in2[95];
    assign G[13] = in1[94] & in2[94];
    assign P[13] = in1[94] ^ in2[94];
    assign G[14] = in1[93] & in2[93];
    assign P[14] = in1[93] ^ in2[93];
    assign G[15] = in1[92] & in2[92];
    assign P[15] = in1[92] ^ in2[92];
    assign G[16] = in1[91] & in2[91];
    assign P[16] = in1[91] ^ in2[91];
    assign G[17] = in1[90] & in2[90];
    assign P[17] = in1[90] ^ in2[90];
    assign G[18] = in1[89] & in2[89];
    assign P[18] = in1[89] ^ in2[89];
    assign G[19] = in1[88] & in2[88];
    assign P[19] = in1[88] ^ in2[88];
    assign G[20] = in1[87] & in2[87];
    assign P[20] = in1[87] ^ in2[87];
    assign G[21] = in1[86] & in2[86];
    assign P[21] = in1[86] ^ in2[86];
    assign G[22] = in1[85] & in2[85];
    assign P[22] = in1[85] ^ in2[85];
    assign G[23] = in1[84] & in2[84];
    assign P[23] = in1[84] ^ in2[84];
    assign G[24] = in1[83] & in2[83];
    assign P[24] = in1[83] ^ in2[83];
    assign G[25] = in1[82] & in2[82];
    assign P[25] = in1[82] ^ in2[82];
    assign G[26] = in1[81] & in2[81];
    assign P[26] = in1[81] ^ in2[81];
    assign G[27] = in1[80] & in2[80];
    assign P[27] = in1[80] ^ in2[80];
    assign G[28] = in1[79] & in2[79];
    assign P[28] = in1[79] ^ in2[79];
    assign G[29] = in1[78] & in2[78];
    assign P[29] = in1[78] ^ in2[78];
    assign G[30] = in1[77] & in2[77];
    assign P[30] = in1[77] ^ in2[77];
    assign G[31] = in1[76] & in2[76];
    assign P[31] = in1[76] ^ in2[76];
    assign G[32] = in1[75] & in2[75];
    assign P[32] = in1[75] ^ in2[75];
    assign G[33] = in1[74] & in2[74];
    assign P[33] = in1[74] ^ in2[74];
    assign G[34] = in1[73] & in2[73];
    assign P[34] = in1[73] ^ in2[73];
    assign G[35] = in1[72] & in2[72];
    assign P[35] = in1[72] ^ in2[72];
    assign G[36] = in1[71] & in2[71];
    assign P[36] = in1[71] ^ in2[71];
    assign G[37] = in1[70] & in2[70];
    assign P[37] = in1[70] ^ in2[70];
    assign G[38] = in1[69] & in2[69];
    assign P[38] = in1[69] ^ in2[69];
    assign G[39] = in1[68] & in2[68];
    assign P[39] = in1[68] ^ in2[68];
    assign G[40] = in1[67] & in2[67];
    assign P[40] = in1[67] ^ in2[67];
    assign G[41] = in1[66] & in2[66];
    assign P[41] = in1[66] ^ in2[66];
    assign G[42] = in1[65] & in2[65];
    assign P[42] = in1[65] ^ in2[65];
    assign G[43] = in1[64] & in2[64];
    assign P[43] = in1[64] ^ in2[64];
    assign G[44] = in1[63] & in2[63];
    assign P[44] = in1[63] ^ in2[63];
    assign G[45] = in1[62] & in2[62];
    assign P[45] = in1[62] ^ in2[62];
    assign G[46] = in1[61] & in2[61];
    assign P[46] = in1[61] ^ in2[61];
    assign G[47] = in1[60] & in2[60];
    assign P[47] = in1[60] ^ in2[60];
    assign G[48] = in1[59] & in2[59];
    assign P[48] = in1[59] ^ in2[59];
    assign G[49] = in1[58] & in2[58];
    assign P[49] = in1[58] ^ in2[58];
    assign G[50] = in1[57] & in2[57];
    assign P[50] = in1[57] ^ in2[57];
    assign G[51] = in1[56] & in2[56];
    assign P[51] = in1[56] ^ in2[56];
    assign G[52] = in1[55] & in2[55];
    assign P[52] = in1[55] ^ in2[55];
    assign G[53] = in1[54] & in2[54];
    assign P[53] = in1[54] ^ in2[54];
    assign G[54] = in1[53] & in2[53];
    assign P[54] = in1[53] ^ in2[53];
    assign G[55] = in1[52] & in2[52];
    assign P[55] = in1[52] ^ in2[52];
    assign G[56] = in1[51] & in2[51];
    assign P[56] = in1[51] ^ in2[51];
    assign G[57] = in1[50] & in2[50];
    assign P[57] = in1[50] ^ in2[50];
    assign G[58] = in1[49] & in2[49];
    assign P[58] = in1[49] ^ in2[49];
    assign G[59] = in1[48] & in2[48];
    assign P[59] = in1[48] ^ in2[48];
    assign G[60] = in1[47] & in2[47];
    assign P[60] = in1[47] ^ in2[47];
    assign G[61] = in1[46] & in2[46];
    assign P[61] = in1[46] ^ in2[46];
    assign G[62] = in1[45] & in2[45];
    assign P[62] = in1[45] ^ in2[45];
    assign G[63] = in1[44] & in2[44];
    assign P[63] = in1[44] ^ in2[44];
    assign G[64] = in1[43] & in2[43];
    assign P[64] = in1[43] ^ in2[43];
    assign G[65] = in1[42] & in2[42];
    assign P[65] = in1[42] ^ in2[42];
    assign G[66] = in1[41] & in2[41];
    assign P[66] = in1[41] ^ in2[41];
    assign G[67] = in1[40] & in2[40];
    assign P[67] = in1[40] ^ in2[40];
    assign G[68] = in1[39] & in2[39];
    assign P[68] = in1[39] ^ in2[39];
    assign G[69] = in1[38] & in2[38];
    assign P[69] = in1[38] ^ in2[38];
    assign G[70] = in1[37] & in2[37];
    assign P[70] = in1[37] ^ in2[37];
    assign G[71] = in1[36] & in2[36];
    assign P[71] = in1[36] ^ in2[36];
    assign G[72] = in1[35] & in2[35];
    assign P[72] = in1[35] ^ in2[35];
    assign G[73] = in1[34] & in2[34];
    assign P[73] = in1[34] ^ in2[34];
    assign G[74] = in1[33] & in2[33];
    assign P[74] = in1[33] ^ in2[33];
    assign G[75] = in1[32] & in2[32];
    assign P[75] = in1[32] ^ in2[32];
    assign G[76] = in1[31] & in2[31];
    assign P[76] = in1[31] ^ in2[31];
    assign G[77] = in1[30] & in2[30];
    assign P[77] = in1[30] ^ in2[30];
    assign G[78] = in1[29] & in2[29];
    assign P[78] = in1[29] ^ in2[29];
    assign G[79] = in1[28] & in2[28];
    assign P[79] = in1[28] ^ in2[28];
    assign G[80] = in1[27] & in2[27];
    assign P[80] = in1[27] ^ in2[27];
    assign G[81] = in1[26] & in2[26];
    assign P[81] = in1[26] ^ in2[26];
    assign G[82] = in1[25] & in2[25];
    assign P[82] = in1[25] ^ in2[25];
    assign G[83] = in1[24] & in2[24];
    assign P[83] = in1[24] ^ in2[24];
    assign G[84] = in1[23] & in2[23];
    assign P[84] = in1[23] ^ in2[23];
    assign G[85] = in1[22] & in2[22];
    assign P[85] = in1[22] ^ in2[22];
    assign G[86] = in1[21] & in2[21];
    assign P[86] = in1[21] ^ in2[21];
    assign G[87] = in1[20] & in2[20];
    assign P[87] = in1[20] ^ in2[20];
    assign G[88] = in1[19] & in2[19];
    assign P[88] = in1[19] ^ in2[19];
    assign G[89] = in1[18] & in2[18];
    assign P[89] = in1[18] ^ in2[18];
    assign G[90] = in1[17] & in2[17];
    assign P[90] = in1[17] ^ in2[17];
    assign G[91] = in1[16] & in2[16];
    assign P[91] = in1[16] ^ in2[16];
    assign G[92] = in1[15] & in2[15];
    assign P[92] = in1[15] ^ in2[15];
    assign G[93] = in1[14] & in2[14];
    assign P[93] = in1[14] ^ in2[14];
    assign G[94] = in1[13] & in2[13];
    assign P[94] = in1[13] ^ in2[13];
    assign G[95] = in1[12] & in2[12];
    assign P[95] = in1[12] ^ in2[12];
    assign G[96] = in1[11] & in2[11];
    assign P[96] = in1[11] ^ in2[11];
    assign G[97] = in1[10] & in2[10];
    assign P[97] = in1[10] ^ in2[10];
    assign G[98] = in1[9] & in2[9];
    assign P[98] = in1[9] ^ in2[9];
    assign G[99] = in1[8] & in2[8];
    assign P[99] = in1[8] ^ in2[8];
    assign G[100] = in1[7] & in2[7];
    assign P[100] = in1[7] ^ in2[7];
    assign G[101] = in1[6] & in2[6];
    assign P[101] = in1[6] ^ in2[6];
    assign G[102] = in1[5] & in2[5];
    assign P[102] = in1[5] ^ in2[5];
    assign G[103] = in1[4] & in2[4];
    assign P[103] = in1[4] ^ in2[4];
    assign G[104] = in1[3] & in2[3];
    assign P[104] = in1[3] ^ in2[3];
    assign G[105] = in1[2] & in2[2];
    assign P[105] = in1[2] ^ in2[2];
    assign G[106] = in1[1] & in2[1];
    assign P[106] = in1[1] ^ in2[1];
    assign G[107] = in1[0] & in2[0];
    assign P[107] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign cout = G[107] | (P[107] & C[107]);
    assign sum = P ^ C;
endmodule

module CLA_107(output [106:0] sum, output cout, input [106:0] in1, input [106:0] in2);

    wire[106:0] G;
    wire[106:0] C;
    wire[106:0] P;

    assign G[0] = in1[106] & in2[106];
    assign P[0] = in1[106] ^ in2[106];
    assign G[1] = in1[105] & in2[105];
    assign P[1] = in1[105] ^ in2[105];
    assign G[2] = in1[104] & in2[104];
    assign P[2] = in1[104] ^ in2[104];
    assign G[3] = in1[103] & in2[103];
    assign P[3] = in1[103] ^ in2[103];
    assign G[4] = in1[102] & in2[102];
    assign P[4] = in1[102] ^ in2[102];
    assign G[5] = in1[101] & in2[101];
    assign P[5] = in1[101] ^ in2[101];
    assign G[6] = in1[100] & in2[100];
    assign P[6] = in1[100] ^ in2[100];
    assign G[7] = in1[99] & in2[99];
    assign P[7] = in1[99] ^ in2[99];
    assign G[8] = in1[98] & in2[98];
    assign P[8] = in1[98] ^ in2[98];
    assign G[9] = in1[97] & in2[97];
    assign P[9] = in1[97] ^ in2[97];
    assign G[10] = in1[96] & in2[96];
    assign P[10] = in1[96] ^ in2[96];
    assign G[11] = in1[95] & in2[95];
    assign P[11] = in1[95] ^ in2[95];
    assign G[12] = in1[94] & in2[94];
    assign P[12] = in1[94] ^ in2[94];
    assign G[13] = in1[93] & in2[93];
    assign P[13] = in1[93] ^ in2[93];
    assign G[14] = in1[92] & in2[92];
    assign P[14] = in1[92] ^ in2[92];
    assign G[15] = in1[91] & in2[91];
    assign P[15] = in1[91] ^ in2[91];
    assign G[16] = in1[90] & in2[90];
    assign P[16] = in1[90] ^ in2[90];
    assign G[17] = in1[89] & in2[89];
    assign P[17] = in1[89] ^ in2[89];
    assign G[18] = in1[88] & in2[88];
    assign P[18] = in1[88] ^ in2[88];
    assign G[19] = in1[87] & in2[87];
    assign P[19] = in1[87] ^ in2[87];
    assign G[20] = in1[86] & in2[86];
    assign P[20] = in1[86] ^ in2[86];
    assign G[21] = in1[85] & in2[85];
    assign P[21] = in1[85] ^ in2[85];
    assign G[22] = in1[84] & in2[84];
    assign P[22] = in1[84] ^ in2[84];
    assign G[23] = in1[83] & in2[83];
    assign P[23] = in1[83] ^ in2[83];
    assign G[24] = in1[82] & in2[82];
    assign P[24] = in1[82] ^ in2[82];
    assign G[25] = in1[81] & in2[81];
    assign P[25] = in1[81] ^ in2[81];
    assign G[26] = in1[80] & in2[80];
    assign P[26] = in1[80] ^ in2[80];
    assign G[27] = in1[79] & in2[79];
    assign P[27] = in1[79] ^ in2[79];
    assign G[28] = in1[78] & in2[78];
    assign P[28] = in1[78] ^ in2[78];
    assign G[29] = in1[77] & in2[77];
    assign P[29] = in1[77] ^ in2[77];
    assign G[30] = in1[76] & in2[76];
    assign P[30] = in1[76] ^ in2[76];
    assign G[31] = in1[75] & in2[75];
    assign P[31] = in1[75] ^ in2[75];
    assign G[32] = in1[74] & in2[74];
    assign P[32] = in1[74] ^ in2[74];
    assign G[33] = in1[73] & in2[73];
    assign P[33] = in1[73] ^ in2[73];
    assign G[34] = in1[72] & in2[72];
    assign P[34] = in1[72] ^ in2[72];
    assign G[35] = in1[71] & in2[71];
    assign P[35] = in1[71] ^ in2[71];
    assign G[36] = in1[70] & in2[70];
    assign P[36] = in1[70] ^ in2[70];
    assign G[37] = in1[69] & in2[69];
    assign P[37] = in1[69] ^ in2[69];
    assign G[38] = in1[68] & in2[68];
    assign P[38] = in1[68] ^ in2[68];
    assign G[39] = in1[67] & in2[67];
    assign P[39] = in1[67] ^ in2[67];
    assign G[40] = in1[66] & in2[66];
    assign P[40] = in1[66] ^ in2[66];
    assign G[41] = in1[65] & in2[65];
    assign P[41] = in1[65] ^ in2[65];
    assign G[42] = in1[64] & in2[64];
    assign P[42] = in1[64] ^ in2[64];
    assign G[43] = in1[63] & in2[63];
    assign P[43] = in1[63] ^ in2[63];
    assign G[44] = in1[62] & in2[62];
    assign P[44] = in1[62] ^ in2[62];
    assign G[45] = in1[61] & in2[61];
    assign P[45] = in1[61] ^ in2[61];
    assign G[46] = in1[60] & in2[60];
    assign P[46] = in1[60] ^ in2[60];
    assign G[47] = in1[59] & in2[59];
    assign P[47] = in1[59] ^ in2[59];
    assign G[48] = in1[58] & in2[58];
    assign P[48] = in1[58] ^ in2[58];
    assign G[49] = in1[57] & in2[57];
    assign P[49] = in1[57] ^ in2[57];
    assign G[50] = in1[56] & in2[56];
    assign P[50] = in1[56] ^ in2[56];
    assign G[51] = in1[55] & in2[55];
    assign P[51] = in1[55] ^ in2[55];
    assign G[52] = in1[54] & in2[54];
    assign P[52] = in1[54] ^ in2[54];
    assign G[53] = in1[53] & in2[53];
    assign P[53] = in1[53] ^ in2[53];
    assign G[54] = in1[52] & in2[52];
    assign P[54] = in1[52] ^ in2[52];
    assign G[55] = in1[51] & in2[51];
    assign P[55] = in1[51] ^ in2[51];
    assign G[56] = in1[50] & in2[50];
    assign P[56] = in1[50] ^ in2[50];
    assign G[57] = in1[49] & in2[49];
    assign P[57] = in1[49] ^ in2[49];
    assign G[58] = in1[48] & in2[48];
    assign P[58] = in1[48] ^ in2[48];
    assign G[59] = in1[47] & in2[47];
    assign P[59] = in1[47] ^ in2[47];
    assign G[60] = in1[46] & in2[46];
    assign P[60] = in1[46] ^ in2[46];
    assign G[61] = in1[45] & in2[45];
    assign P[61] = in1[45] ^ in2[45];
    assign G[62] = in1[44] & in2[44];
    assign P[62] = in1[44] ^ in2[44];
    assign G[63] = in1[43] & in2[43];
    assign P[63] = in1[43] ^ in2[43];
    assign G[64] = in1[42] & in2[42];
    assign P[64] = in1[42] ^ in2[42];
    assign G[65] = in1[41] & in2[41];
    assign P[65] = in1[41] ^ in2[41];
    assign G[66] = in1[40] & in2[40];
    assign P[66] = in1[40] ^ in2[40];
    assign G[67] = in1[39] & in2[39];
    assign P[67] = in1[39] ^ in2[39];
    assign G[68] = in1[38] & in2[38];
    assign P[68] = in1[38] ^ in2[38];
    assign G[69] = in1[37] & in2[37];
    assign P[69] = in1[37] ^ in2[37];
    assign G[70] = in1[36] & in2[36];
    assign P[70] = in1[36] ^ in2[36];
    assign G[71] = in1[35] & in2[35];
    assign P[71] = in1[35] ^ in2[35];
    assign G[72] = in1[34] & in2[34];
    assign P[72] = in1[34] ^ in2[34];
    assign G[73] = in1[33] & in2[33];
    assign P[73] = in1[33] ^ in2[33];
    assign G[74] = in1[32] & in2[32];
    assign P[74] = in1[32] ^ in2[32];
    assign G[75] = in1[31] & in2[31];
    assign P[75] = in1[31] ^ in2[31];
    assign G[76] = in1[30] & in2[30];
    assign P[76] = in1[30] ^ in2[30];
    assign G[77] = in1[29] & in2[29];
    assign P[77] = in1[29] ^ in2[29];
    assign G[78] = in1[28] & in2[28];
    assign P[78] = in1[28] ^ in2[28];
    assign G[79] = in1[27] & in2[27];
    assign P[79] = in1[27] ^ in2[27];
    assign G[80] = in1[26] & in2[26];
    assign P[80] = in1[26] ^ in2[26];
    assign G[81] = in1[25] & in2[25];
    assign P[81] = in1[25] ^ in2[25];
    assign G[82] = in1[24] & in2[24];
    assign P[82] = in1[24] ^ in2[24];
    assign G[83] = in1[23] & in2[23];
    assign P[83] = in1[23] ^ in2[23];
    assign G[84] = in1[22] & in2[22];
    assign P[84] = in1[22] ^ in2[22];
    assign G[85] = in1[21] & in2[21];
    assign P[85] = in1[21] ^ in2[21];
    assign G[86] = in1[20] & in2[20];
    assign P[86] = in1[20] ^ in2[20];
    assign G[87] = in1[19] & in2[19];
    assign P[87] = in1[19] ^ in2[19];
    assign G[88] = in1[18] & in2[18];
    assign P[88] = in1[18] ^ in2[18];
    assign G[89] = in1[17] & in2[17];
    assign P[89] = in1[17] ^ in2[17];
    assign G[90] = in1[16] & in2[16];
    assign P[90] = in1[16] ^ in2[16];
    assign G[91] = in1[15] & in2[15];
    assign P[91] = in1[15] ^ in2[15];
    assign G[92] = in1[14] & in2[14];
    assign P[92] = in1[14] ^ in2[14];
    assign G[93] = in1[13] & in2[13];
    assign P[93] = in1[13] ^ in2[13];
    assign G[94] = in1[12] & in2[12];
    assign P[94] = in1[12] ^ in2[12];
    assign G[95] = in1[11] & in2[11];
    assign P[95] = in1[11] ^ in2[11];
    assign G[96] = in1[10] & in2[10];
    assign P[96] = in1[10] ^ in2[10];
    assign G[97] = in1[9] & in2[9];
    assign P[97] = in1[9] ^ in2[9];
    assign G[98] = in1[8] & in2[8];
    assign P[98] = in1[8] ^ in2[8];
    assign G[99] = in1[7] & in2[7];
    assign P[99] = in1[7] ^ in2[7];
    assign G[100] = in1[6] & in2[6];
    assign P[100] = in1[6] ^ in2[6];
    assign G[101] = in1[5] & in2[5];
    assign P[101] = in1[5] ^ in2[5];
    assign G[102] = in1[4] & in2[4];
    assign P[102] = in1[4] ^ in2[4];
    assign G[103] = in1[3] & in2[3];
    assign P[103] = in1[3] ^ in2[3];
    assign G[104] = in1[2] & in2[2];
    assign P[104] = in1[2] ^ in2[2];
    assign G[105] = in1[1] & in2[1];
    assign P[105] = in1[1] ^ in2[1];
    assign G[106] = in1[0] & in2[0];
    assign P[106] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign cout = G[106] | (P[106] & C[106]);
    assign sum = P ^ C;
endmodule

module CLA_106(output [105:0] sum, output cout, input [105:0] in1, input [105:0] in2);

    wire[105:0] G;
    wire[105:0] C;
    wire[105:0] P;

    assign G[0] = in1[105] & in2[105];
    assign P[0] = in1[105] ^ in2[105];
    assign G[1] = in1[104] & in2[104];
    assign P[1] = in1[104] ^ in2[104];
    assign G[2] = in1[103] & in2[103];
    assign P[2] = in1[103] ^ in2[103];
    assign G[3] = in1[102] & in2[102];
    assign P[3] = in1[102] ^ in2[102];
    assign G[4] = in1[101] & in2[101];
    assign P[4] = in1[101] ^ in2[101];
    assign G[5] = in1[100] & in2[100];
    assign P[5] = in1[100] ^ in2[100];
    assign G[6] = in1[99] & in2[99];
    assign P[6] = in1[99] ^ in2[99];
    assign G[7] = in1[98] & in2[98];
    assign P[7] = in1[98] ^ in2[98];
    assign G[8] = in1[97] & in2[97];
    assign P[8] = in1[97] ^ in2[97];
    assign G[9] = in1[96] & in2[96];
    assign P[9] = in1[96] ^ in2[96];
    assign G[10] = in1[95] & in2[95];
    assign P[10] = in1[95] ^ in2[95];
    assign G[11] = in1[94] & in2[94];
    assign P[11] = in1[94] ^ in2[94];
    assign G[12] = in1[93] & in2[93];
    assign P[12] = in1[93] ^ in2[93];
    assign G[13] = in1[92] & in2[92];
    assign P[13] = in1[92] ^ in2[92];
    assign G[14] = in1[91] & in2[91];
    assign P[14] = in1[91] ^ in2[91];
    assign G[15] = in1[90] & in2[90];
    assign P[15] = in1[90] ^ in2[90];
    assign G[16] = in1[89] & in2[89];
    assign P[16] = in1[89] ^ in2[89];
    assign G[17] = in1[88] & in2[88];
    assign P[17] = in1[88] ^ in2[88];
    assign G[18] = in1[87] & in2[87];
    assign P[18] = in1[87] ^ in2[87];
    assign G[19] = in1[86] & in2[86];
    assign P[19] = in1[86] ^ in2[86];
    assign G[20] = in1[85] & in2[85];
    assign P[20] = in1[85] ^ in2[85];
    assign G[21] = in1[84] & in2[84];
    assign P[21] = in1[84] ^ in2[84];
    assign G[22] = in1[83] & in2[83];
    assign P[22] = in1[83] ^ in2[83];
    assign G[23] = in1[82] & in2[82];
    assign P[23] = in1[82] ^ in2[82];
    assign G[24] = in1[81] & in2[81];
    assign P[24] = in1[81] ^ in2[81];
    assign G[25] = in1[80] & in2[80];
    assign P[25] = in1[80] ^ in2[80];
    assign G[26] = in1[79] & in2[79];
    assign P[26] = in1[79] ^ in2[79];
    assign G[27] = in1[78] & in2[78];
    assign P[27] = in1[78] ^ in2[78];
    assign G[28] = in1[77] & in2[77];
    assign P[28] = in1[77] ^ in2[77];
    assign G[29] = in1[76] & in2[76];
    assign P[29] = in1[76] ^ in2[76];
    assign G[30] = in1[75] & in2[75];
    assign P[30] = in1[75] ^ in2[75];
    assign G[31] = in1[74] & in2[74];
    assign P[31] = in1[74] ^ in2[74];
    assign G[32] = in1[73] & in2[73];
    assign P[32] = in1[73] ^ in2[73];
    assign G[33] = in1[72] & in2[72];
    assign P[33] = in1[72] ^ in2[72];
    assign G[34] = in1[71] & in2[71];
    assign P[34] = in1[71] ^ in2[71];
    assign G[35] = in1[70] & in2[70];
    assign P[35] = in1[70] ^ in2[70];
    assign G[36] = in1[69] & in2[69];
    assign P[36] = in1[69] ^ in2[69];
    assign G[37] = in1[68] & in2[68];
    assign P[37] = in1[68] ^ in2[68];
    assign G[38] = in1[67] & in2[67];
    assign P[38] = in1[67] ^ in2[67];
    assign G[39] = in1[66] & in2[66];
    assign P[39] = in1[66] ^ in2[66];
    assign G[40] = in1[65] & in2[65];
    assign P[40] = in1[65] ^ in2[65];
    assign G[41] = in1[64] & in2[64];
    assign P[41] = in1[64] ^ in2[64];
    assign G[42] = in1[63] & in2[63];
    assign P[42] = in1[63] ^ in2[63];
    assign G[43] = in1[62] & in2[62];
    assign P[43] = in1[62] ^ in2[62];
    assign G[44] = in1[61] & in2[61];
    assign P[44] = in1[61] ^ in2[61];
    assign G[45] = in1[60] & in2[60];
    assign P[45] = in1[60] ^ in2[60];
    assign G[46] = in1[59] & in2[59];
    assign P[46] = in1[59] ^ in2[59];
    assign G[47] = in1[58] & in2[58];
    assign P[47] = in1[58] ^ in2[58];
    assign G[48] = in1[57] & in2[57];
    assign P[48] = in1[57] ^ in2[57];
    assign G[49] = in1[56] & in2[56];
    assign P[49] = in1[56] ^ in2[56];
    assign G[50] = in1[55] & in2[55];
    assign P[50] = in1[55] ^ in2[55];
    assign G[51] = in1[54] & in2[54];
    assign P[51] = in1[54] ^ in2[54];
    assign G[52] = in1[53] & in2[53];
    assign P[52] = in1[53] ^ in2[53];
    assign G[53] = in1[52] & in2[52];
    assign P[53] = in1[52] ^ in2[52];
    assign G[54] = in1[51] & in2[51];
    assign P[54] = in1[51] ^ in2[51];
    assign G[55] = in1[50] & in2[50];
    assign P[55] = in1[50] ^ in2[50];
    assign G[56] = in1[49] & in2[49];
    assign P[56] = in1[49] ^ in2[49];
    assign G[57] = in1[48] & in2[48];
    assign P[57] = in1[48] ^ in2[48];
    assign G[58] = in1[47] & in2[47];
    assign P[58] = in1[47] ^ in2[47];
    assign G[59] = in1[46] & in2[46];
    assign P[59] = in1[46] ^ in2[46];
    assign G[60] = in1[45] & in2[45];
    assign P[60] = in1[45] ^ in2[45];
    assign G[61] = in1[44] & in2[44];
    assign P[61] = in1[44] ^ in2[44];
    assign G[62] = in1[43] & in2[43];
    assign P[62] = in1[43] ^ in2[43];
    assign G[63] = in1[42] & in2[42];
    assign P[63] = in1[42] ^ in2[42];
    assign G[64] = in1[41] & in2[41];
    assign P[64] = in1[41] ^ in2[41];
    assign G[65] = in1[40] & in2[40];
    assign P[65] = in1[40] ^ in2[40];
    assign G[66] = in1[39] & in2[39];
    assign P[66] = in1[39] ^ in2[39];
    assign G[67] = in1[38] & in2[38];
    assign P[67] = in1[38] ^ in2[38];
    assign G[68] = in1[37] & in2[37];
    assign P[68] = in1[37] ^ in2[37];
    assign G[69] = in1[36] & in2[36];
    assign P[69] = in1[36] ^ in2[36];
    assign G[70] = in1[35] & in2[35];
    assign P[70] = in1[35] ^ in2[35];
    assign G[71] = in1[34] & in2[34];
    assign P[71] = in1[34] ^ in2[34];
    assign G[72] = in1[33] & in2[33];
    assign P[72] = in1[33] ^ in2[33];
    assign G[73] = in1[32] & in2[32];
    assign P[73] = in1[32] ^ in2[32];
    assign G[74] = in1[31] & in2[31];
    assign P[74] = in1[31] ^ in2[31];
    assign G[75] = in1[30] & in2[30];
    assign P[75] = in1[30] ^ in2[30];
    assign G[76] = in1[29] & in2[29];
    assign P[76] = in1[29] ^ in2[29];
    assign G[77] = in1[28] & in2[28];
    assign P[77] = in1[28] ^ in2[28];
    assign G[78] = in1[27] & in2[27];
    assign P[78] = in1[27] ^ in2[27];
    assign G[79] = in1[26] & in2[26];
    assign P[79] = in1[26] ^ in2[26];
    assign G[80] = in1[25] & in2[25];
    assign P[80] = in1[25] ^ in2[25];
    assign G[81] = in1[24] & in2[24];
    assign P[81] = in1[24] ^ in2[24];
    assign G[82] = in1[23] & in2[23];
    assign P[82] = in1[23] ^ in2[23];
    assign G[83] = in1[22] & in2[22];
    assign P[83] = in1[22] ^ in2[22];
    assign G[84] = in1[21] & in2[21];
    assign P[84] = in1[21] ^ in2[21];
    assign G[85] = in1[20] & in2[20];
    assign P[85] = in1[20] ^ in2[20];
    assign G[86] = in1[19] & in2[19];
    assign P[86] = in1[19] ^ in2[19];
    assign G[87] = in1[18] & in2[18];
    assign P[87] = in1[18] ^ in2[18];
    assign G[88] = in1[17] & in2[17];
    assign P[88] = in1[17] ^ in2[17];
    assign G[89] = in1[16] & in2[16];
    assign P[89] = in1[16] ^ in2[16];
    assign G[90] = in1[15] & in2[15];
    assign P[90] = in1[15] ^ in2[15];
    assign G[91] = in1[14] & in2[14];
    assign P[91] = in1[14] ^ in2[14];
    assign G[92] = in1[13] & in2[13];
    assign P[92] = in1[13] ^ in2[13];
    assign G[93] = in1[12] & in2[12];
    assign P[93] = in1[12] ^ in2[12];
    assign G[94] = in1[11] & in2[11];
    assign P[94] = in1[11] ^ in2[11];
    assign G[95] = in1[10] & in2[10];
    assign P[95] = in1[10] ^ in2[10];
    assign G[96] = in1[9] & in2[9];
    assign P[96] = in1[9] ^ in2[9];
    assign G[97] = in1[8] & in2[8];
    assign P[97] = in1[8] ^ in2[8];
    assign G[98] = in1[7] & in2[7];
    assign P[98] = in1[7] ^ in2[7];
    assign G[99] = in1[6] & in2[6];
    assign P[99] = in1[6] ^ in2[6];
    assign G[100] = in1[5] & in2[5];
    assign P[100] = in1[5] ^ in2[5];
    assign G[101] = in1[4] & in2[4];
    assign P[101] = in1[4] ^ in2[4];
    assign G[102] = in1[3] & in2[3];
    assign P[102] = in1[3] ^ in2[3];
    assign G[103] = in1[2] & in2[2];
    assign P[103] = in1[2] ^ in2[2];
    assign G[104] = in1[1] & in2[1];
    assign P[104] = in1[1] ^ in2[1];
    assign G[105] = in1[0] & in2[0];
    assign P[105] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign cout = G[105] | (P[105] & C[105]);
    assign sum = P ^ C;
endmodule

module CLA_105(output [104:0] sum, output cout, input [104:0] in1, input [104:0] in2);

    wire[104:0] G;
    wire[104:0] C;
    wire[104:0] P;

    assign G[0] = in1[104] & in2[104];
    assign P[0] = in1[104] ^ in2[104];
    assign G[1] = in1[103] & in2[103];
    assign P[1] = in1[103] ^ in2[103];
    assign G[2] = in1[102] & in2[102];
    assign P[2] = in1[102] ^ in2[102];
    assign G[3] = in1[101] & in2[101];
    assign P[3] = in1[101] ^ in2[101];
    assign G[4] = in1[100] & in2[100];
    assign P[4] = in1[100] ^ in2[100];
    assign G[5] = in1[99] & in2[99];
    assign P[5] = in1[99] ^ in2[99];
    assign G[6] = in1[98] & in2[98];
    assign P[6] = in1[98] ^ in2[98];
    assign G[7] = in1[97] & in2[97];
    assign P[7] = in1[97] ^ in2[97];
    assign G[8] = in1[96] & in2[96];
    assign P[8] = in1[96] ^ in2[96];
    assign G[9] = in1[95] & in2[95];
    assign P[9] = in1[95] ^ in2[95];
    assign G[10] = in1[94] & in2[94];
    assign P[10] = in1[94] ^ in2[94];
    assign G[11] = in1[93] & in2[93];
    assign P[11] = in1[93] ^ in2[93];
    assign G[12] = in1[92] & in2[92];
    assign P[12] = in1[92] ^ in2[92];
    assign G[13] = in1[91] & in2[91];
    assign P[13] = in1[91] ^ in2[91];
    assign G[14] = in1[90] & in2[90];
    assign P[14] = in1[90] ^ in2[90];
    assign G[15] = in1[89] & in2[89];
    assign P[15] = in1[89] ^ in2[89];
    assign G[16] = in1[88] & in2[88];
    assign P[16] = in1[88] ^ in2[88];
    assign G[17] = in1[87] & in2[87];
    assign P[17] = in1[87] ^ in2[87];
    assign G[18] = in1[86] & in2[86];
    assign P[18] = in1[86] ^ in2[86];
    assign G[19] = in1[85] & in2[85];
    assign P[19] = in1[85] ^ in2[85];
    assign G[20] = in1[84] & in2[84];
    assign P[20] = in1[84] ^ in2[84];
    assign G[21] = in1[83] & in2[83];
    assign P[21] = in1[83] ^ in2[83];
    assign G[22] = in1[82] & in2[82];
    assign P[22] = in1[82] ^ in2[82];
    assign G[23] = in1[81] & in2[81];
    assign P[23] = in1[81] ^ in2[81];
    assign G[24] = in1[80] & in2[80];
    assign P[24] = in1[80] ^ in2[80];
    assign G[25] = in1[79] & in2[79];
    assign P[25] = in1[79] ^ in2[79];
    assign G[26] = in1[78] & in2[78];
    assign P[26] = in1[78] ^ in2[78];
    assign G[27] = in1[77] & in2[77];
    assign P[27] = in1[77] ^ in2[77];
    assign G[28] = in1[76] & in2[76];
    assign P[28] = in1[76] ^ in2[76];
    assign G[29] = in1[75] & in2[75];
    assign P[29] = in1[75] ^ in2[75];
    assign G[30] = in1[74] & in2[74];
    assign P[30] = in1[74] ^ in2[74];
    assign G[31] = in1[73] & in2[73];
    assign P[31] = in1[73] ^ in2[73];
    assign G[32] = in1[72] & in2[72];
    assign P[32] = in1[72] ^ in2[72];
    assign G[33] = in1[71] & in2[71];
    assign P[33] = in1[71] ^ in2[71];
    assign G[34] = in1[70] & in2[70];
    assign P[34] = in1[70] ^ in2[70];
    assign G[35] = in1[69] & in2[69];
    assign P[35] = in1[69] ^ in2[69];
    assign G[36] = in1[68] & in2[68];
    assign P[36] = in1[68] ^ in2[68];
    assign G[37] = in1[67] & in2[67];
    assign P[37] = in1[67] ^ in2[67];
    assign G[38] = in1[66] & in2[66];
    assign P[38] = in1[66] ^ in2[66];
    assign G[39] = in1[65] & in2[65];
    assign P[39] = in1[65] ^ in2[65];
    assign G[40] = in1[64] & in2[64];
    assign P[40] = in1[64] ^ in2[64];
    assign G[41] = in1[63] & in2[63];
    assign P[41] = in1[63] ^ in2[63];
    assign G[42] = in1[62] & in2[62];
    assign P[42] = in1[62] ^ in2[62];
    assign G[43] = in1[61] & in2[61];
    assign P[43] = in1[61] ^ in2[61];
    assign G[44] = in1[60] & in2[60];
    assign P[44] = in1[60] ^ in2[60];
    assign G[45] = in1[59] & in2[59];
    assign P[45] = in1[59] ^ in2[59];
    assign G[46] = in1[58] & in2[58];
    assign P[46] = in1[58] ^ in2[58];
    assign G[47] = in1[57] & in2[57];
    assign P[47] = in1[57] ^ in2[57];
    assign G[48] = in1[56] & in2[56];
    assign P[48] = in1[56] ^ in2[56];
    assign G[49] = in1[55] & in2[55];
    assign P[49] = in1[55] ^ in2[55];
    assign G[50] = in1[54] & in2[54];
    assign P[50] = in1[54] ^ in2[54];
    assign G[51] = in1[53] & in2[53];
    assign P[51] = in1[53] ^ in2[53];
    assign G[52] = in1[52] & in2[52];
    assign P[52] = in1[52] ^ in2[52];
    assign G[53] = in1[51] & in2[51];
    assign P[53] = in1[51] ^ in2[51];
    assign G[54] = in1[50] & in2[50];
    assign P[54] = in1[50] ^ in2[50];
    assign G[55] = in1[49] & in2[49];
    assign P[55] = in1[49] ^ in2[49];
    assign G[56] = in1[48] & in2[48];
    assign P[56] = in1[48] ^ in2[48];
    assign G[57] = in1[47] & in2[47];
    assign P[57] = in1[47] ^ in2[47];
    assign G[58] = in1[46] & in2[46];
    assign P[58] = in1[46] ^ in2[46];
    assign G[59] = in1[45] & in2[45];
    assign P[59] = in1[45] ^ in2[45];
    assign G[60] = in1[44] & in2[44];
    assign P[60] = in1[44] ^ in2[44];
    assign G[61] = in1[43] & in2[43];
    assign P[61] = in1[43] ^ in2[43];
    assign G[62] = in1[42] & in2[42];
    assign P[62] = in1[42] ^ in2[42];
    assign G[63] = in1[41] & in2[41];
    assign P[63] = in1[41] ^ in2[41];
    assign G[64] = in1[40] & in2[40];
    assign P[64] = in1[40] ^ in2[40];
    assign G[65] = in1[39] & in2[39];
    assign P[65] = in1[39] ^ in2[39];
    assign G[66] = in1[38] & in2[38];
    assign P[66] = in1[38] ^ in2[38];
    assign G[67] = in1[37] & in2[37];
    assign P[67] = in1[37] ^ in2[37];
    assign G[68] = in1[36] & in2[36];
    assign P[68] = in1[36] ^ in2[36];
    assign G[69] = in1[35] & in2[35];
    assign P[69] = in1[35] ^ in2[35];
    assign G[70] = in1[34] & in2[34];
    assign P[70] = in1[34] ^ in2[34];
    assign G[71] = in1[33] & in2[33];
    assign P[71] = in1[33] ^ in2[33];
    assign G[72] = in1[32] & in2[32];
    assign P[72] = in1[32] ^ in2[32];
    assign G[73] = in1[31] & in2[31];
    assign P[73] = in1[31] ^ in2[31];
    assign G[74] = in1[30] & in2[30];
    assign P[74] = in1[30] ^ in2[30];
    assign G[75] = in1[29] & in2[29];
    assign P[75] = in1[29] ^ in2[29];
    assign G[76] = in1[28] & in2[28];
    assign P[76] = in1[28] ^ in2[28];
    assign G[77] = in1[27] & in2[27];
    assign P[77] = in1[27] ^ in2[27];
    assign G[78] = in1[26] & in2[26];
    assign P[78] = in1[26] ^ in2[26];
    assign G[79] = in1[25] & in2[25];
    assign P[79] = in1[25] ^ in2[25];
    assign G[80] = in1[24] & in2[24];
    assign P[80] = in1[24] ^ in2[24];
    assign G[81] = in1[23] & in2[23];
    assign P[81] = in1[23] ^ in2[23];
    assign G[82] = in1[22] & in2[22];
    assign P[82] = in1[22] ^ in2[22];
    assign G[83] = in1[21] & in2[21];
    assign P[83] = in1[21] ^ in2[21];
    assign G[84] = in1[20] & in2[20];
    assign P[84] = in1[20] ^ in2[20];
    assign G[85] = in1[19] & in2[19];
    assign P[85] = in1[19] ^ in2[19];
    assign G[86] = in1[18] & in2[18];
    assign P[86] = in1[18] ^ in2[18];
    assign G[87] = in1[17] & in2[17];
    assign P[87] = in1[17] ^ in2[17];
    assign G[88] = in1[16] & in2[16];
    assign P[88] = in1[16] ^ in2[16];
    assign G[89] = in1[15] & in2[15];
    assign P[89] = in1[15] ^ in2[15];
    assign G[90] = in1[14] & in2[14];
    assign P[90] = in1[14] ^ in2[14];
    assign G[91] = in1[13] & in2[13];
    assign P[91] = in1[13] ^ in2[13];
    assign G[92] = in1[12] & in2[12];
    assign P[92] = in1[12] ^ in2[12];
    assign G[93] = in1[11] & in2[11];
    assign P[93] = in1[11] ^ in2[11];
    assign G[94] = in1[10] & in2[10];
    assign P[94] = in1[10] ^ in2[10];
    assign G[95] = in1[9] & in2[9];
    assign P[95] = in1[9] ^ in2[9];
    assign G[96] = in1[8] & in2[8];
    assign P[96] = in1[8] ^ in2[8];
    assign G[97] = in1[7] & in2[7];
    assign P[97] = in1[7] ^ in2[7];
    assign G[98] = in1[6] & in2[6];
    assign P[98] = in1[6] ^ in2[6];
    assign G[99] = in1[5] & in2[5];
    assign P[99] = in1[5] ^ in2[5];
    assign G[100] = in1[4] & in2[4];
    assign P[100] = in1[4] ^ in2[4];
    assign G[101] = in1[3] & in2[3];
    assign P[101] = in1[3] ^ in2[3];
    assign G[102] = in1[2] & in2[2];
    assign P[102] = in1[2] ^ in2[2];
    assign G[103] = in1[1] & in2[1];
    assign P[103] = in1[1] ^ in2[1];
    assign G[104] = in1[0] & in2[0];
    assign P[104] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign cout = G[104] | (P[104] & C[104]);
    assign sum = P ^ C;
endmodule

module CLA_104(output [103:0] sum, output cout, input [103:0] in1, input [103:0] in2);

    wire[103:0] G;
    wire[103:0] C;
    wire[103:0] P;

    assign G[0] = in1[103] & in2[103];
    assign P[0] = in1[103] ^ in2[103];
    assign G[1] = in1[102] & in2[102];
    assign P[1] = in1[102] ^ in2[102];
    assign G[2] = in1[101] & in2[101];
    assign P[2] = in1[101] ^ in2[101];
    assign G[3] = in1[100] & in2[100];
    assign P[3] = in1[100] ^ in2[100];
    assign G[4] = in1[99] & in2[99];
    assign P[4] = in1[99] ^ in2[99];
    assign G[5] = in1[98] & in2[98];
    assign P[5] = in1[98] ^ in2[98];
    assign G[6] = in1[97] & in2[97];
    assign P[6] = in1[97] ^ in2[97];
    assign G[7] = in1[96] & in2[96];
    assign P[7] = in1[96] ^ in2[96];
    assign G[8] = in1[95] & in2[95];
    assign P[8] = in1[95] ^ in2[95];
    assign G[9] = in1[94] & in2[94];
    assign P[9] = in1[94] ^ in2[94];
    assign G[10] = in1[93] & in2[93];
    assign P[10] = in1[93] ^ in2[93];
    assign G[11] = in1[92] & in2[92];
    assign P[11] = in1[92] ^ in2[92];
    assign G[12] = in1[91] & in2[91];
    assign P[12] = in1[91] ^ in2[91];
    assign G[13] = in1[90] & in2[90];
    assign P[13] = in1[90] ^ in2[90];
    assign G[14] = in1[89] & in2[89];
    assign P[14] = in1[89] ^ in2[89];
    assign G[15] = in1[88] & in2[88];
    assign P[15] = in1[88] ^ in2[88];
    assign G[16] = in1[87] & in2[87];
    assign P[16] = in1[87] ^ in2[87];
    assign G[17] = in1[86] & in2[86];
    assign P[17] = in1[86] ^ in2[86];
    assign G[18] = in1[85] & in2[85];
    assign P[18] = in1[85] ^ in2[85];
    assign G[19] = in1[84] & in2[84];
    assign P[19] = in1[84] ^ in2[84];
    assign G[20] = in1[83] & in2[83];
    assign P[20] = in1[83] ^ in2[83];
    assign G[21] = in1[82] & in2[82];
    assign P[21] = in1[82] ^ in2[82];
    assign G[22] = in1[81] & in2[81];
    assign P[22] = in1[81] ^ in2[81];
    assign G[23] = in1[80] & in2[80];
    assign P[23] = in1[80] ^ in2[80];
    assign G[24] = in1[79] & in2[79];
    assign P[24] = in1[79] ^ in2[79];
    assign G[25] = in1[78] & in2[78];
    assign P[25] = in1[78] ^ in2[78];
    assign G[26] = in1[77] & in2[77];
    assign P[26] = in1[77] ^ in2[77];
    assign G[27] = in1[76] & in2[76];
    assign P[27] = in1[76] ^ in2[76];
    assign G[28] = in1[75] & in2[75];
    assign P[28] = in1[75] ^ in2[75];
    assign G[29] = in1[74] & in2[74];
    assign P[29] = in1[74] ^ in2[74];
    assign G[30] = in1[73] & in2[73];
    assign P[30] = in1[73] ^ in2[73];
    assign G[31] = in1[72] & in2[72];
    assign P[31] = in1[72] ^ in2[72];
    assign G[32] = in1[71] & in2[71];
    assign P[32] = in1[71] ^ in2[71];
    assign G[33] = in1[70] & in2[70];
    assign P[33] = in1[70] ^ in2[70];
    assign G[34] = in1[69] & in2[69];
    assign P[34] = in1[69] ^ in2[69];
    assign G[35] = in1[68] & in2[68];
    assign P[35] = in1[68] ^ in2[68];
    assign G[36] = in1[67] & in2[67];
    assign P[36] = in1[67] ^ in2[67];
    assign G[37] = in1[66] & in2[66];
    assign P[37] = in1[66] ^ in2[66];
    assign G[38] = in1[65] & in2[65];
    assign P[38] = in1[65] ^ in2[65];
    assign G[39] = in1[64] & in2[64];
    assign P[39] = in1[64] ^ in2[64];
    assign G[40] = in1[63] & in2[63];
    assign P[40] = in1[63] ^ in2[63];
    assign G[41] = in1[62] & in2[62];
    assign P[41] = in1[62] ^ in2[62];
    assign G[42] = in1[61] & in2[61];
    assign P[42] = in1[61] ^ in2[61];
    assign G[43] = in1[60] & in2[60];
    assign P[43] = in1[60] ^ in2[60];
    assign G[44] = in1[59] & in2[59];
    assign P[44] = in1[59] ^ in2[59];
    assign G[45] = in1[58] & in2[58];
    assign P[45] = in1[58] ^ in2[58];
    assign G[46] = in1[57] & in2[57];
    assign P[46] = in1[57] ^ in2[57];
    assign G[47] = in1[56] & in2[56];
    assign P[47] = in1[56] ^ in2[56];
    assign G[48] = in1[55] & in2[55];
    assign P[48] = in1[55] ^ in2[55];
    assign G[49] = in1[54] & in2[54];
    assign P[49] = in1[54] ^ in2[54];
    assign G[50] = in1[53] & in2[53];
    assign P[50] = in1[53] ^ in2[53];
    assign G[51] = in1[52] & in2[52];
    assign P[51] = in1[52] ^ in2[52];
    assign G[52] = in1[51] & in2[51];
    assign P[52] = in1[51] ^ in2[51];
    assign G[53] = in1[50] & in2[50];
    assign P[53] = in1[50] ^ in2[50];
    assign G[54] = in1[49] & in2[49];
    assign P[54] = in1[49] ^ in2[49];
    assign G[55] = in1[48] & in2[48];
    assign P[55] = in1[48] ^ in2[48];
    assign G[56] = in1[47] & in2[47];
    assign P[56] = in1[47] ^ in2[47];
    assign G[57] = in1[46] & in2[46];
    assign P[57] = in1[46] ^ in2[46];
    assign G[58] = in1[45] & in2[45];
    assign P[58] = in1[45] ^ in2[45];
    assign G[59] = in1[44] & in2[44];
    assign P[59] = in1[44] ^ in2[44];
    assign G[60] = in1[43] & in2[43];
    assign P[60] = in1[43] ^ in2[43];
    assign G[61] = in1[42] & in2[42];
    assign P[61] = in1[42] ^ in2[42];
    assign G[62] = in1[41] & in2[41];
    assign P[62] = in1[41] ^ in2[41];
    assign G[63] = in1[40] & in2[40];
    assign P[63] = in1[40] ^ in2[40];
    assign G[64] = in1[39] & in2[39];
    assign P[64] = in1[39] ^ in2[39];
    assign G[65] = in1[38] & in2[38];
    assign P[65] = in1[38] ^ in2[38];
    assign G[66] = in1[37] & in2[37];
    assign P[66] = in1[37] ^ in2[37];
    assign G[67] = in1[36] & in2[36];
    assign P[67] = in1[36] ^ in2[36];
    assign G[68] = in1[35] & in2[35];
    assign P[68] = in1[35] ^ in2[35];
    assign G[69] = in1[34] & in2[34];
    assign P[69] = in1[34] ^ in2[34];
    assign G[70] = in1[33] & in2[33];
    assign P[70] = in1[33] ^ in2[33];
    assign G[71] = in1[32] & in2[32];
    assign P[71] = in1[32] ^ in2[32];
    assign G[72] = in1[31] & in2[31];
    assign P[72] = in1[31] ^ in2[31];
    assign G[73] = in1[30] & in2[30];
    assign P[73] = in1[30] ^ in2[30];
    assign G[74] = in1[29] & in2[29];
    assign P[74] = in1[29] ^ in2[29];
    assign G[75] = in1[28] & in2[28];
    assign P[75] = in1[28] ^ in2[28];
    assign G[76] = in1[27] & in2[27];
    assign P[76] = in1[27] ^ in2[27];
    assign G[77] = in1[26] & in2[26];
    assign P[77] = in1[26] ^ in2[26];
    assign G[78] = in1[25] & in2[25];
    assign P[78] = in1[25] ^ in2[25];
    assign G[79] = in1[24] & in2[24];
    assign P[79] = in1[24] ^ in2[24];
    assign G[80] = in1[23] & in2[23];
    assign P[80] = in1[23] ^ in2[23];
    assign G[81] = in1[22] & in2[22];
    assign P[81] = in1[22] ^ in2[22];
    assign G[82] = in1[21] & in2[21];
    assign P[82] = in1[21] ^ in2[21];
    assign G[83] = in1[20] & in2[20];
    assign P[83] = in1[20] ^ in2[20];
    assign G[84] = in1[19] & in2[19];
    assign P[84] = in1[19] ^ in2[19];
    assign G[85] = in1[18] & in2[18];
    assign P[85] = in1[18] ^ in2[18];
    assign G[86] = in1[17] & in2[17];
    assign P[86] = in1[17] ^ in2[17];
    assign G[87] = in1[16] & in2[16];
    assign P[87] = in1[16] ^ in2[16];
    assign G[88] = in1[15] & in2[15];
    assign P[88] = in1[15] ^ in2[15];
    assign G[89] = in1[14] & in2[14];
    assign P[89] = in1[14] ^ in2[14];
    assign G[90] = in1[13] & in2[13];
    assign P[90] = in1[13] ^ in2[13];
    assign G[91] = in1[12] & in2[12];
    assign P[91] = in1[12] ^ in2[12];
    assign G[92] = in1[11] & in2[11];
    assign P[92] = in1[11] ^ in2[11];
    assign G[93] = in1[10] & in2[10];
    assign P[93] = in1[10] ^ in2[10];
    assign G[94] = in1[9] & in2[9];
    assign P[94] = in1[9] ^ in2[9];
    assign G[95] = in1[8] & in2[8];
    assign P[95] = in1[8] ^ in2[8];
    assign G[96] = in1[7] & in2[7];
    assign P[96] = in1[7] ^ in2[7];
    assign G[97] = in1[6] & in2[6];
    assign P[97] = in1[6] ^ in2[6];
    assign G[98] = in1[5] & in2[5];
    assign P[98] = in1[5] ^ in2[5];
    assign G[99] = in1[4] & in2[4];
    assign P[99] = in1[4] ^ in2[4];
    assign G[100] = in1[3] & in2[3];
    assign P[100] = in1[3] ^ in2[3];
    assign G[101] = in1[2] & in2[2];
    assign P[101] = in1[2] ^ in2[2];
    assign G[102] = in1[1] & in2[1];
    assign P[102] = in1[1] ^ in2[1];
    assign G[103] = in1[0] & in2[0];
    assign P[103] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign cout = G[103] | (P[103] & C[103]);
    assign sum = P ^ C;
endmodule

module CLA_103(output [102:0] sum, output cout, input [102:0] in1, input [102:0] in2);

    wire[102:0] G;
    wire[102:0] C;
    wire[102:0] P;

    assign G[0] = in1[102] & in2[102];
    assign P[0] = in1[102] ^ in2[102];
    assign G[1] = in1[101] & in2[101];
    assign P[1] = in1[101] ^ in2[101];
    assign G[2] = in1[100] & in2[100];
    assign P[2] = in1[100] ^ in2[100];
    assign G[3] = in1[99] & in2[99];
    assign P[3] = in1[99] ^ in2[99];
    assign G[4] = in1[98] & in2[98];
    assign P[4] = in1[98] ^ in2[98];
    assign G[5] = in1[97] & in2[97];
    assign P[5] = in1[97] ^ in2[97];
    assign G[6] = in1[96] & in2[96];
    assign P[6] = in1[96] ^ in2[96];
    assign G[7] = in1[95] & in2[95];
    assign P[7] = in1[95] ^ in2[95];
    assign G[8] = in1[94] & in2[94];
    assign P[8] = in1[94] ^ in2[94];
    assign G[9] = in1[93] & in2[93];
    assign P[9] = in1[93] ^ in2[93];
    assign G[10] = in1[92] & in2[92];
    assign P[10] = in1[92] ^ in2[92];
    assign G[11] = in1[91] & in2[91];
    assign P[11] = in1[91] ^ in2[91];
    assign G[12] = in1[90] & in2[90];
    assign P[12] = in1[90] ^ in2[90];
    assign G[13] = in1[89] & in2[89];
    assign P[13] = in1[89] ^ in2[89];
    assign G[14] = in1[88] & in2[88];
    assign P[14] = in1[88] ^ in2[88];
    assign G[15] = in1[87] & in2[87];
    assign P[15] = in1[87] ^ in2[87];
    assign G[16] = in1[86] & in2[86];
    assign P[16] = in1[86] ^ in2[86];
    assign G[17] = in1[85] & in2[85];
    assign P[17] = in1[85] ^ in2[85];
    assign G[18] = in1[84] & in2[84];
    assign P[18] = in1[84] ^ in2[84];
    assign G[19] = in1[83] & in2[83];
    assign P[19] = in1[83] ^ in2[83];
    assign G[20] = in1[82] & in2[82];
    assign P[20] = in1[82] ^ in2[82];
    assign G[21] = in1[81] & in2[81];
    assign P[21] = in1[81] ^ in2[81];
    assign G[22] = in1[80] & in2[80];
    assign P[22] = in1[80] ^ in2[80];
    assign G[23] = in1[79] & in2[79];
    assign P[23] = in1[79] ^ in2[79];
    assign G[24] = in1[78] & in2[78];
    assign P[24] = in1[78] ^ in2[78];
    assign G[25] = in1[77] & in2[77];
    assign P[25] = in1[77] ^ in2[77];
    assign G[26] = in1[76] & in2[76];
    assign P[26] = in1[76] ^ in2[76];
    assign G[27] = in1[75] & in2[75];
    assign P[27] = in1[75] ^ in2[75];
    assign G[28] = in1[74] & in2[74];
    assign P[28] = in1[74] ^ in2[74];
    assign G[29] = in1[73] & in2[73];
    assign P[29] = in1[73] ^ in2[73];
    assign G[30] = in1[72] & in2[72];
    assign P[30] = in1[72] ^ in2[72];
    assign G[31] = in1[71] & in2[71];
    assign P[31] = in1[71] ^ in2[71];
    assign G[32] = in1[70] & in2[70];
    assign P[32] = in1[70] ^ in2[70];
    assign G[33] = in1[69] & in2[69];
    assign P[33] = in1[69] ^ in2[69];
    assign G[34] = in1[68] & in2[68];
    assign P[34] = in1[68] ^ in2[68];
    assign G[35] = in1[67] & in2[67];
    assign P[35] = in1[67] ^ in2[67];
    assign G[36] = in1[66] & in2[66];
    assign P[36] = in1[66] ^ in2[66];
    assign G[37] = in1[65] & in2[65];
    assign P[37] = in1[65] ^ in2[65];
    assign G[38] = in1[64] & in2[64];
    assign P[38] = in1[64] ^ in2[64];
    assign G[39] = in1[63] & in2[63];
    assign P[39] = in1[63] ^ in2[63];
    assign G[40] = in1[62] & in2[62];
    assign P[40] = in1[62] ^ in2[62];
    assign G[41] = in1[61] & in2[61];
    assign P[41] = in1[61] ^ in2[61];
    assign G[42] = in1[60] & in2[60];
    assign P[42] = in1[60] ^ in2[60];
    assign G[43] = in1[59] & in2[59];
    assign P[43] = in1[59] ^ in2[59];
    assign G[44] = in1[58] & in2[58];
    assign P[44] = in1[58] ^ in2[58];
    assign G[45] = in1[57] & in2[57];
    assign P[45] = in1[57] ^ in2[57];
    assign G[46] = in1[56] & in2[56];
    assign P[46] = in1[56] ^ in2[56];
    assign G[47] = in1[55] & in2[55];
    assign P[47] = in1[55] ^ in2[55];
    assign G[48] = in1[54] & in2[54];
    assign P[48] = in1[54] ^ in2[54];
    assign G[49] = in1[53] & in2[53];
    assign P[49] = in1[53] ^ in2[53];
    assign G[50] = in1[52] & in2[52];
    assign P[50] = in1[52] ^ in2[52];
    assign G[51] = in1[51] & in2[51];
    assign P[51] = in1[51] ^ in2[51];
    assign G[52] = in1[50] & in2[50];
    assign P[52] = in1[50] ^ in2[50];
    assign G[53] = in1[49] & in2[49];
    assign P[53] = in1[49] ^ in2[49];
    assign G[54] = in1[48] & in2[48];
    assign P[54] = in1[48] ^ in2[48];
    assign G[55] = in1[47] & in2[47];
    assign P[55] = in1[47] ^ in2[47];
    assign G[56] = in1[46] & in2[46];
    assign P[56] = in1[46] ^ in2[46];
    assign G[57] = in1[45] & in2[45];
    assign P[57] = in1[45] ^ in2[45];
    assign G[58] = in1[44] & in2[44];
    assign P[58] = in1[44] ^ in2[44];
    assign G[59] = in1[43] & in2[43];
    assign P[59] = in1[43] ^ in2[43];
    assign G[60] = in1[42] & in2[42];
    assign P[60] = in1[42] ^ in2[42];
    assign G[61] = in1[41] & in2[41];
    assign P[61] = in1[41] ^ in2[41];
    assign G[62] = in1[40] & in2[40];
    assign P[62] = in1[40] ^ in2[40];
    assign G[63] = in1[39] & in2[39];
    assign P[63] = in1[39] ^ in2[39];
    assign G[64] = in1[38] & in2[38];
    assign P[64] = in1[38] ^ in2[38];
    assign G[65] = in1[37] & in2[37];
    assign P[65] = in1[37] ^ in2[37];
    assign G[66] = in1[36] & in2[36];
    assign P[66] = in1[36] ^ in2[36];
    assign G[67] = in1[35] & in2[35];
    assign P[67] = in1[35] ^ in2[35];
    assign G[68] = in1[34] & in2[34];
    assign P[68] = in1[34] ^ in2[34];
    assign G[69] = in1[33] & in2[33];
    assign P[69] = in1[33] ^ in2[33];
    assign G[70] = in1[32] & in2[32];
    assign P[70] = in1[32] ^ in2[32];
    assign G[71] = in1[31] & in2[31];
    assign P[71] = in1[31] ^ in2[31];
    assign G[72] = in1[30] & in2[30];
    assign P[72] = in1[30] ^ in2[30];
    assign G[73] = in1[29] & in2[29];
    assign P[73] = in1[29] ^ in2[29];
    assign G[74] = in1[28] & in2[28];
    assign P[74] = in1[28] ^ in2[28];
    assign G[75] = in1[27] & in2[27];
    assign P[75] = in1[27] ^ in2[27];
    assign G[76] = in1[26] & in2[26];
    assign P[76] = in1[26] ^ in2[26];
    assign G[77] = in1[25] & in2[25];
    assign P[77] = in1[25] ^ in2[25];
    assign G[78] = in1[24] & in2[24];
    assign P[78] = in1[24] ^ in2[24];
    assign G[79] = in1[23] & in2[23];
    assign P[79] = in1[23] ^ in2[23];
    assign G[80] = in1[22] & in2[22];
    assign P[80] = in1[22] ^ in2[22];
    assign G[81] = in1[21] & in2[21];
    assign P[81] = in1[21] ^ in2[21];
    assign G[82] = in1[20] & in2[20];
    assign P[82] = in1[20] ^ in2[20];
    assign G[83] = in1[19] & in2[19];
    assign P[83] = in1[19] ^ in2[19];
    assign G[84] = in1[18] & in2[18];
    assign P[84] = in1[18] ^ in2[18];
    assign G[85] = in1[17] & in2[17];
    assign P[85] = in1[17] ^ in2[17];
    assign G[86] = in1[16] & in2[16];
    assign P[86] = in1[16] ^ in2[16];
    assign G[87] = in1[15] & in2[15];
    assign P[87] = in1[15] ^ in2[15];
    assign G[88] = in1[14] & in2[14];
    assign P[88] = in1[14] ^ in2[14];
    assign G[89] = in1[13] & in2[13];
    assign P[89] = in1[13] ^ in2[13];
    assign G[90] = in1[12] & in2[12];
    assign P[90] = in1[12] ^ in2[12];
    assign G[91] = in1[11] & in2[11];
    assign P[91] = in1[11] ^ in2[11];
    assign G[92] = in1[10] & in2[10];
    assign P[92] = in1[10] ^ in2[10];
    assign G[93] = in1[9] & in2[9];
    assign P[93] = in1[9] ^ in2[9];
    assign G[94] = in1[8] & in2[8];
    assign P[94] = in1[8] ^ in2[8];
    assign G[95] = in1[7] & in2[7];
    assign P[95] = in1[7] ^ in2[7];
    assign G[96] = in1[6] & in2[6];
    assign P[96] = in1[6] ^ in2[6];
    assign G[97] = in1[5] & in2[5];
    assign P[97] = in1[5] ^ in2[5];
    assign G[98] = in1[4] & in2[4];
    assign P[98] = in1[4] ^ in2[4];
    assign G[99] = in1[3] & in2[3];
    assign P[99] = in1[3] ^ in2[3];
    assign G[100] = in1[2] & in2[2];
    assign P[100] = in1[2] ^ in2[2];
    assign G[101] = in1[1] & in2[1];
    assign P[101] = in1[1] ^ in2[1];
    assign G[102] = in1[0] & in2[0];
    assign P[102] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign cout = G[102] | (P[102] & C[102]);
    assign sum = P ^ C;
endmodule

module CLA_102(output [101:0] sum, output cout, input [101:0] in1, input [101:0] in2);

    wire[101:0] G;
    wire[101:0] C;
    wire[101:0] P;

    assign G[0] = in1[101] & in2[101];
    assign P[0] = in1[101] ^ in2[101];
    assign G[1] = in1[100] & in2[100];
    assign P[1] = in1[100] ^ in2[100];
    assign G[2] = in1[99] & in2[99];
    assign P[2] = in1[99] ^ in2[99];
    assign G[3] = in1[98] & in2[98];
    assign P[3] = in1[98] ^ in2[98];
    assign G[4] = in1[97] & in2[97];
    assign P[4] = in1[97] ^ in2[97];
    assign G[5] = in1[96] & in2[96];
    assign P[5] = in1[96] ^ in2[96];
    assign G[6] = in1[95] & in2[95];
    assign P[6] = in1[95] ^ in2[95];
    assign G[7] = in1[94] & in2[94];
    assign P[7] = in1[94] ^ in2[94];
    assign G[8] = in1[93] & in2[93];
    assign P[8] = in1[93] ^ in2[93];
    assign G[9] = in1[92] & in2[92];
    assign P[9] = in1[92] ^ in2[92];
    assign G[10] = in1[91] & in2[91];
    assign P[10] = in1[91] ^ in2[91];
    assign G[11] = in1[90] & in2[90];
    assign P[11] = in1[90] ^ in2[90];
    assign G[12] = in1[89] & in2[89];
    assign P[12] = in1[89] ^ in2[89];
    assign G[13] = in1[88] & in2[88];
    assign P[13] = in1[88] ^ in2[88];
    assign G[14] = in1[87] & in2[87];
    assign P[14] = in1[87] ^ in2[87];
    assign G[15] = in1[86] & in2[86];
    assign P[15] = in1[86] ^ in2[86];
    assign G[16] = in1[85] & in2[85];
    assign P[16] = in1[85] ^ in2[85];
    assign G[17] = in1[84] & in2[84];
    assign P[17] = in1[84] ^ in2[84];
    assign G[18] = in1[83] & in2[83];
    assign P[18] = in1[83] ^ in2[83];
    assign G[19] = in1[82] & in2[82];
    assign P[19] = in1[82] ^ in2[82];
    assign G[20] = in1[81] & in2[81];
    assign P[20] = in1[81] ^ in2[81];
    assign G[21] = in1[80] & in2[80];
    assign P[21] = in1[80] ^ in2[80];
    assign G[22] = in1[79] & in2[79];
    assign P[22] = in1[79] ^ in2[79];
    assign G[23] = in1[78] & in2[78];
    assign P[23] = in1[78] ^ in2[78];
    assign G[24] = in1[77] & in2[77];
    assign P[24] = in1[77] ^ in2[77];
    assign G[25] = in1[76] & in2[76];
    assign P[25] = in1[76] ^ in2[76];
    assign G[26] = in1[75] & in2[75];
    assign P[26] = in1[75] ^ in2[75];
    assign G[27] = in1[74] & in2[74];
    assign P[27] = in1[74] ^ in2[74];
    assign G[28] = in1[73] & in2[73];
    assign P[28] = in1[73] ^ in2[73];
    assign G[29] = in1[72] & in2[72];
    assign P[29] = in1[72] ^ in2[72];
    assign G[30] = in1[71] & in2[71];
    assign P[30] = in1[71] ^ in2[71];
    assign G[31] = in1[70] & in2[70];
    assign P[31] = in1[70] ^ in2[70];
    assign G[32] = in1[69] & in2[69];
    assign P[32] = in1[69] ^ in2[69];
    assign G[33] = in1[68] & in2[68];
    assign P[33] = in1[68] ^ in2[68];
    assign G[34] = in1[67] & in2[67];
    assign P[34] = in1[67] ^ in2[67];
    assign G[35] = in1[66] & in2[66];
    assign P[35] = in1[66] ^ in2[66];
    assign G[36] = in1[65] & in2[65];
    assign P[36] = in1[65] ^ in2[65];
    assign G[37] = in1[64] & in2[64];
    assign P[37] = in1[64] ^ in2[64];
    assign G[38] = in1[63] & in2[63];
    assign P[38] = in1[63] ^ in2[63];
    assign G[39] = in1[62] & in2[62];
    assign P[39] = in1[62] ^ in2[62];
    assign G[40] = in1[61] & in2[61];
    assign P[40] = in1[61] ^ in2[61];
    assign G[41] = in1[60] & in2[60];
    assign P[41] = in1[60] ^ in2[60];
    assign G[42] = in1[59] & in2[59];
    assign P[42] = in1[59] ^ in2[59];
    assign G[43] = in1[58] & in2[58];
    assign P[43] = in1[58] ^ in2[58];
    assign G[44] = in1[57] & in2[57];
    assign P[44] = in1[57] ^ in2[57];
    assign G[45] = in1[56] & in2[56];
    assign P[45] = in1[56] ^ in2[56];
    assign G[46] = in1[55] & in2[55];
    assign P[46] = in1[55] ^ in2[55];
    assign G[47] = in1[54] & in2[54];
    assign P[47] = in1[54] ^ in2[54];
    assign G[48] = in1[53] & in2[53];
    assign P[48] = in1[53] ^ in2[53];
    assign G[49] = in1[52] & in2[52];
    assign P[49] = in1[52] ^ in2[52];
    assign G[50] = in1[51] & in2[51];
    assign P[50] = in1[51] ^ in2[51];
    assign G[51] = in1[50] & in2[50];
    assign P[51] = in1[50] ^ in2[50];
    assign G[52] = in1[49] & in2[49];
    assign P[52] = in1[49] ^ in2[49];
    assign G[53] = in1[48] & in2[48];
    assign P[53] = in1[48] ^ in2[48];
    assign G[54] = in1[47] & in2[47];
    assign P[54] = in1[47] ^ in2[47];
    assign G[55] = in1[46] & in2[46];
    assign P[55] = in1[46] ^ in2[46];
    assign G[56] = in1[45] & in2[45];
    assign P[56] = in1[45] ^ in2[45];
    assign G[57] = in1[44] & in2[44];
    assign P[57] = in1[44] ^ in2[44];
    assign G[58] = in1[43] & in2[43];
    assign P[58] = in1[43] ^ in2[43];
    assign G[59] = in1[42] & in2[42];
    assign P[59] = in1[42] ^ in2[42];
    assign G[60] = in1[41] & in2[41];
    assign P[60] = in1[41] ^ in2[41];
    assign G[61] = in1[40] & in2[40];
    assign P[61] = in1[40] ^ in2[40];
    assign G[62] = in1[39] & in2[39];
    assign P[62] = in1[39] ^ in2[39];
    assign G[63] = in1[38] & in2[38];
    assign P[63] = in1[38] ^ in2[38];
    assign G[64] = in1[37] & in2[37];
    assign P[64] = in1[37] ^ in2[37];
    assign G[65] = in1[36] & in2[36];
    assign P[65] = in1[36] ^ in2[36];
    assign G[66] = in1[35] & in2[35];
    assign P[66] = in1[35] ^ in2[35];
    assign G[67] = in1[34] & in2[34];
    assign P[67] = in1[34] ^ in2[34];
    assign G[68] = in1[33] & in2[33];
    assign P[68] = in1[33] ^ in2[33];
    assign G[69] = in1[32] & in2[32];
    assign P[69] = in1[32] ^ in2[32];
    assign G[70] = in1[31] & in2[31];
    assign P[70] = in1[31] ^ in2[31];
    assign G[71] = in1[30] & in2[30];
    assign P[71] = in1[30] ^ in2[30];
    assign G[72] = in1[29] & in2[29];
    assign P[72] = in1[29] ^ in2[29];
    assign G[73] = in1[28] & in2[28];
    assign P[73] = in1[28] ^ in2[28];
    assign G[74] = in1[27] & in2[27];
    assign P[74] = in1[27] ^ in2[27];
    assign G[75] = in1[26] & in2[26];
    assign P[75] = in1[26] ^ in2[26];
    assign G[76] = in1[25] & in2[25];
    assign P[76] = in1[25] ^ in2[25];
    assign G[77] = in1[24] & in2[24];
    assign P[77] = in1[24] ^ in2[24];
    assign G[78] = in1[23] & in2[23];
    assign P[78] = in1[23] ^ in2[23];
    assign G[79] = in1[22] & in2[22];
    assign P[79] = in1[22] ^ in2[22];
    assign G[80] = in1[21] & in2[21];
    assign P[80] = in1[21] ^ in2[21];
    assign G[81] = in1[20] & in2[20];
    assign P[81] = in1[20] ^ in2[20];
    assign G[82] = in1[19] & in2[19];
    assign P[82] = in1[19] ^ in2[19];
    assign G[83] = in1[18] & in2[18];
    assign P[83] = in1[18] ^ in2[18];
    assign G[84] = in1[17] & in2[17];
    assign P[84] = in1[17] ^ in2[17];
    assign G[85] = in1[16] & in2[16];
    assign P[85] = in1[16] ^ in2[16];
    assign G[86] = in1[15] & in2[15];
    assign P[86] = in1[15] ^ in2[15];
    assign G[87] = in1[14] & in2[14];
    assign P[87] = in1[14] ^ in2[14];
    assign G[88] = in1[13] & in2[13];
    assign P[88] = in1[13] ^ in2[13];
    assign G[89] = in1[12] & in2[12];
    assign P[89] = in1[12] ^ in2[12];
    assign G[90] = in1[11] & in2[11];
    assign P[90] = in1[11] ^ in2[11];
    assign G[91] = in1[10] & in2[10];
    assign P[91] = in1[10] ^ in2[10];
    assign G[92] = in1[9] & in2[9];
    assign P[92] = in1[9] ^ in2[9];
    assign G[93] = in1[8] & in2[8];
    assign P[93] = in1[8] ^ in2[8];
    assign G[94] = in1[7] & in2[7];
    assign P[94] = in1[7] ^ in2[7];
    assign G[95] = in1[6] & in2[6];
    assign P[95] = in1[6] ^ in2[6];
    assign G[96] = in1[5] & in2[5];
    assign P[96] = in1[5] ^ in2[5];
    assign G[97] = in1[4] & in2[4];
    assign P[97] = in1[4] ^ in2[4];
    assign G[98] = in1[3] & in2[3];
    assign P[98] = in1[3] ^ in2[3];
    assign G[99] = in1[2] & in2[2];
    assign P[99] = in1[2] ^ in2[2];
    assign G[100] = in1[1] & in2[1];
    assign P[100] = in1[1] ^ in2[1];
    assign G[101] = in1[0] & in2[0];
    assign P[101] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign cout = G[101] | (P[101] & C[101]);
    assign sum = P ^ C;
endmodule

module CLA_101(output [100:0] sum, output cout, input [100:0] in1, input [100:0] in2);

    wire[100:0] G;
    wire[100:0] C;
    wire[100:0] P;

    assign G[0] = in1[100] & in2[100];
    assign P[0] = in1[100] ^ in2[100];
    assign G[1] = in1[99] & in2[99];
    assign P[1] = in1[99] ^ in2[99];
    assign G[2] = in1[98] & in2[98];
    assign P[2] = in1[98] ^ in2[98];
    assign G[3] = in1[97] & in2[97];
    assign P[3] = in1[97] ^ in2[97];
    assign G[4] = in1[96] & in2[96];
    assign P[4] = in1[96] ^ in2[96];
    assign G[5] = in1[95] & in2[95];
    assign P[5] = in1[95] ^ in2[95];
    assign G[6] = in1[94] & in2[94];
    assign P[6] = in1[94] ^ in2[94];
    assign G[7] = in1[93] & in2[93];
    assign P[7] = in1[93] ^ in2[93];
    assign G[8] = in1[92] & in2[92];
    assign P[8] = in1[92] ^ in2[92];
    assign G[9] = in1[91] & in2[91];
    assign P[9] = in1[91] ^ in2[91];
    assign G[10] = in1[90] & in2[90];
    assign P[10] = in1[90] ^ in2[90];
    assign G[11] = in1[89] & in2[89];
    assign P[11] = in1[89] ^ in2[89];
    assign G[12] = in1[88] & in2[88];
    assign P[12] = in1[88] ^ in2[88];
    assign G[13] = in1[87] & in2[87];
    assign P[13] = in1[87] ^ in2[87];
    assign G[14] = in1[86] & in2[86];
    assign P[14] = in1[86] ^ in2[86];
    assign G[15] = in1[85] & in2[85];
    assign P[15] = in1[85] ^ in2[85];
    assign G[16] = in1[84] & in2[84];
    assign P[16] = in1[84] ^ in2[84];
    assign G[17] = in1[83] & in2[83];
    assign P[17] = in1[83] ^ in2[83];
    assign G[18] = in1[82] & in2[82];
    assign P[18] = in1[82] ^ in2[82];
    assign G[19] = in1[81] & in2[81];
    assign P[19] = in1[81] ^ in2[81];
    assign G[20] = in1[80] & in2[80];
    assign P[20] = in1[80] ^ in2[80];
    assign G[21] = in1[79] & in2[79];
    assign P[21] = in1[79] ^ in2[79];
    assign G[22] = in1[78] & in2[78];
    assign P[22] = in1[78] ^ in2[78];
    assign G[23] = in1[77] & in2[77];
    assign P[23] = in1[77] ^ in2[77];
    assign G[24] = in1[76] & in2[76];
    assign P[24] = in1[76] ^ in2[76];
    assign G[25] = in1[75] & in2[75];
    assign P[25] = in1[75] ^ in2[75];
    assign G[26] = in1[74] & in2[74];
    assign P[26] = in1[74] ^ in2[74];
    assign G[27] = in1[73] & in2[73];
    assign P[27] = in1[73] ^ in2[73];
    assign G[28] = in1[72] & in2[72];
    assign P[28] = in1[72] ^ in2[72];
    assign G[29] = in1[71] & in2[71];
    assign P[29] = in1[71] ^ in2[71];
    assign G[30] = in1[70] & in2[70];
    assign P[30] = in1[70] ^ in2[70];
    assign G[31] = in1[69] & in2[69];
    assign P[31] = in1[69] ^ in2[69];
    assign G[32] = in1[68] & in2[68];
    assign P[32] = in1[68] ^ in2[68];
    assign G[33] = in1[67] & in2[67];
    assign P[33] = in1[67] ^ in2[67];
    assign G[34] = in1[66] & in2[66];
    assign P[34] = in1[66] ^ in2[66];
    assign G[35] = in1[65] & in2[65];
    assign P[35] = in1[65] ^ in2[65];
    assign G[36] = in1[64] & in2[64];
    assign P[36] = in1[64] ^ in2[64];
    assign G[37] = in1[63] & in2[63];
    assign P[37] = in1[63] ^ in2[63];
    assign G[38] = in1[62] & in2[62];
    assign P[38] = in1[62] ^ in2[62];
    assign G[39] = in1[61] & in2[61];
    assign P[39] = in1[61] ^ in2[61];
    assign G[40] = in1[60] & in2[60];
    assign P[40] = in1[60] ^ in2[60];
    assign G[41] = in1[59] & in2[59];
    assign P[41] = in1[59] ^ in2[59];
    assign G[42] = in1[58] & in2[58];
    assign P[42] = in1[58] ^ in2[58];
    assign G[43] = in1[57] & in2[57];
    assign P[43] = in1[57] ^ in2[57];
    assign G[44] = in1[56] & in2[56];
    assign P[44] = in1[56] ^ in2[56];
    assign G[45] = in1[55] & in2[55];
    assign P[45] = in1[55] ^ in2[55];
    assign G[46] = in1[54] & in2[54];
    assign P[46] = in1[54] ^ in2[54];
    assign G[47] = in1[53] & in2[53];
    assign P[47] = in1[53] ^ in2[53];
    assign G[48] = in1[52] & in2[52];
    assign P[48] = in1[52] ^ in2[52];
    assign G[49] = in1[51] & in2[51];
    assign P[49] = in1[51] ^ in2[51];
    assign G[50] = in1[50] & in2[50];
    assign P[50] = in1[50] ^ in2[50];
    assign G[51] = in1[49] & in2[49];
    assign P[51] = in1[49] ^ in2[49];
    assign G[52] = in1[48] & in2[48];
    assign P[52] = in1[48] ^ in2[48];
    assign G[53] = in1[47] & in2[47];
    assign P[53] = in1[47] ^ in2[47];
    assign G[54] = in1[46] & in2[46];
    assign P[54] = in1[46] ^ in2[46];
    assign G[55] = in1[45] & in2[45];
    assign P[55] = in1[45] ^ in2[45];
    assign G[56] = in1[44] & in2[44];
    assign P[56] = in1[44] ^ in2[44];
    assign G[57] = in1[43] & in2[43];
    assign P[57] = in1[43] ^ in2[43];
    assign G[58] = in1[42] & in2[42];
    assign P[58] = in1[42] ^ in2[42];
    assign G[59] = in1[41] & in2[41];
    assign P[59] = in1[41] ^ in2[41];
    assign G[60] = in1[40] & in2[40];
    assign P[60] = in1[40] ^ in2[40];
    assign G[61] = in1[39] & in2[39];
    assign P[61] = in1[39] ^ in2[39];
    assign G[62] = in1[38] & in2[38];
    assign P[62] = in1[38] ^ in2[38];
    assign G[63] = in1[37] & in2[37];
    assign P[63] = in1[37] ^ in2[37];
    assign G[64] = in1[36] & in2[36];
    assign P[64] = in1[36] ^ in2[36];
    assign G[65] = in1[35] & in2[35];
    assign P[65] = in1[35] ^ in2[35];
    assign G[66] = in1[34] & in2[34];
    assign P[66] = in1[34] ^ in2[34];
    assign G[67] = in1[33] & in2[33];
    assign P[67] = in1[33] ^ in2[33];
    assign G[68] = in1[32] & in2[32];
    assign P[68] = in1[32] ^ in2[32];
    assign G[69] = in1[31] & in2[31];
    assign P[69] = in1[31] ^ in2[31];
    assign G[70] = in1[30] & in2[30];
    assign P[70] = in1[30] ^ in2[30];
    assign G[71] = in1[29] & in2[29];
    assign P[71] = in1[29] ^ in2[29];
    assign G[72] = in1[28] & in2[28];
    assign P[72] = in1[28] ^ in2[28];
    assign G[73] = in1[27] & in2[27];
    assign P[73] = in1[27] ^ in2[27];
    assign G[74] = in1[26] & in2[26];
    assign P[74] = in1[26] ^ in2[26];
    assign G[75] = in1[25] & in2[25];
    assign P[75] = in1[25] ^ in2[25];
    assign G[76] = in1[24] & in2[24];
    assign P[76] = in1[24] ^ in2[24];
    assign G[77] = in1[23] & in2[23];
    assign P[77] = in1[23] ^ in2[23];
    assign G[78] = in1[22] & in2[22];
    assign P[78] = in1[22] ^ in2[22];
    assign G[79] = in1[21] & in2[21];
    assign P[79] = in1[21] ^ in2[21];
    assign G[80] = in1[20] & in2[20];
    assign P[80] = in1[20] ^ in2[20];
    assign G[81] = in1[19] & in2[19];
    assign P[81] = in1[19] ^ in2[19];
    assign G[82] = in1[18] & in2[18];
    assign P[82] = in1[18] ^ in2[18];
    assign G[83] = in1[17] & in2[17];
    assign P[83] = in1[17] ^ in2[17];
    assign G[84] = in1[16] & in2[16];
    assign P[84] = in1[16] ^ in2[16];
    assign G[85] = in1[15] & in2[15];
    assign P[85] = in1[15] ^ in2[15];
    assign G[86] = in1[14] & in2[14];
    assign P[86] = in1[14] ^ in2[14];
    assign G[87] = in1[13] & in2[13];
    assign P[87] = in1[13] ^ in2[13];
    assign G[88] = in1[12] & in2[12];
    assign P[88] = in1[12] ^ in2[12];
    assign G[89] = in1[11] & in2[11];
    assign P[89] = in1[11] ^ in2[11];
    assign G[90] = in1[10] & in2[10];
    assign P[90] = in1[10] ^ in2[10];
    assign G[91] = in1[9] & in2[9];
    assign P[91] = in1[9] ^ in2[9];
    assign G[92] = in1[8] & in2[8];
    assign P[92] = in1[8] ^ in2[8];
    assign G[93] = in1[7] & in2[7];
    assign P[93] = in1[7] ^ in2[7];
    assign G[94] = in1[6] & in2[6];
    assign P[94] = in1[6] ^ in2[6];
    assign G[95] = in1[5] & in2[5];
    assign P[95] = in1[5] ^ in2[5];
    assign G[96] = in1[4] & in2[4];
    assign P[96] = in1[4] ^ in2[4];
    assign G[97] = in1[3] & in2[3];
    assign P[97] = in1[3] ^ in2[3];
    assign G[98] = in1[2] & in2[2];
    assign P[98] = in1[2] ^ in2[2];
    assign G[99] = in1[1] & in2[1];
    assign P[99] = in1[1] ^ in2[1];
    assign G[100] = in1[0] & in2[0];
    assign P[100] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign cout = G[100] | (P[100] & C[100]);
    assign sum = P ^ C;
endmodule

module CLA_100(output [99:0] sum, output cout, input [99:0] in1, input [99:0] in2);

    wire[99:0] G;
    wire[99:0] C;
    wire[99:0] P;

    assign G[0] = in1[99] & in2[99];
    assign P[0] = in1[99] ^ in2[99];
    assign G[1] = in1[98] & in2[98];
    assign P[1] = in1[98] ^ in2[98];
    assign G[2] = in1[97] & in2[97];
    assign P[2] = in1[97] ^ in2[97];
    assign G[3] = in1[96] & in2[96];
    assign P[3] = in1[96] ^ in2[96];
    assign G[4] = in1[95] & in2[95];
    assign P[4] = in1[95] ^ in2[95];
    assign G[5] = in1[94] & in2[94];
    assign P[5] = in1[94] ^ in2[94];
    assign G[6] = in1[93] & in2[93];
    assign P[6] = in1[93] ^ in2[93];
    assign G[7] = in1[92] & in2[92];
    assign P[7] = in1[92] ^ in2[92];
    assign G[8] = in1[91] & in2[91];
    assign P[8] = in1[91] ^ in2[91];
    assign G[9] = in1[90] & in2[90];
    assign P[9] = in1[90] ^ in2[90];
    assign G[10] = in1[89] & in2[89];
    assign P[10] = in1[89] ^ in2[89];
    assign G[11] = in1[88] & in2[88];
    assign P[11] = in1[88] ^ in2[88];
    assign G[12] = in1[87] & in2[87];
    assign P[12] = in1[87] ^ in2[87];
    assign G[13] = in1[86] & in2[86];
    assign P[13] = in1[86] ^ in2[86];
    assign G[14] = in1[85] & in2[85];
    assign P[14] = in1[85] ^ in2[85];
    assign G[15] = in1[84] & in2[84];
    assign P[15] = in1[84] ^ in2[84];
    assign G[16] = in1[83] & in2[83];
    assign P[16] = in1[83] ^ in2[83];
    assign G[17] = in1[82] & in2[82];
    assign P[17] = in1[82] ^ in2[82];
    assign G[18] = in1[81] & in2[81];
    assign P[18] = in1[81] ^ in2[81];
    assign G[19] = in1[80] & in2[80];
    assign P[19] = in1[80] ^ in2[80];
    assign G[20] = in1[79] & in2[79];
    assign P[20] = in1[79] ^ in2[79];
    assign G[21] = in1[78] & in2[78];
    assign P[21] = in1[78] ^ in2[78];
    assign G[22] = in1[77] & in2[77];
    assign P[22] = in1[77] ^ in2[77];
    assign G[23] = in1[76] & in2[76];
    assign P[23] = in1[76] ^ in2[76];
    assign G[24] = in1[75] & in2[75];
    assign P[24] = in1[75] ^ in2[75];
    assign G[25] = in1[74] & in2[74];
    assign P[25] = in1[74] ^ in2[74];
    assign G[26] = in1[73] & in2[73];
    assign P[26] = in1[73] ^ in2[73];
    assign G[27] = in1[72] & in2[72];
    assign P[27] = in1[72] ^ in2[72];
    assign G[28] = in1[71] & in2[71];
    assign P[28] = in1[71] ^ in2[71];
    assign G[29] = in1[70] & in2[70];
    assign P[29] = in1[70] ^ in2[70];
    assign G[30] = in1[69] & in2[69];
    assign P[30] = in1[69] ^ in2[69];
    assign G[31] = in1[68] & in2[68];
    assign P[31] = in1[68] ^ in2[68];
    assign G[32] = in1[67] & in2[67];
    assign P[32] = in1[67] ^ in2[67];
    assign G[33] = in1[66] & in2[66];
    assign P[33] = in1[66] ^ in2[66];
    assign G[34] = in1[65] & in2[65];
    assign P[34] = in1[65] ^ in2[65];
    assign G[35] = in1[64] & in2[64];
    assign P[35] = in1[64] ^ in2[64];
    assign G[36] = in1[63] & in2[63];
    assign P[36] = in1[63] ^ in2[63];
    assign G[37] = in1[62] & in2[62];
    assign P[37] = in1[62] ^ in2[62];
    assign G[38] = in1[61] & in2[61];
    assign P[38] = in1[61] ^ in2[61];
    assign G[39] = in1[60] & in2[60];
    assign P[39] = in1[60] ^ in2[60];
    assign G[40] = in1[59] & in2[59];
    assign P[40] = in1[59] ^ in2[59];
    assign G[41] = in1[58] & in2[58];
    assign P[41] = in1[58] ^ in2[58];
    assign G[42] = in1[57] & in2[57];
    assign P[42] = in1[57] ^ in2[57];
    assign G[43] = in1[56] & in2[56];
    assign P[43] = in1[56] ^ in2[56];
    assign G[44] = in1[55] & in2[55];
    assign P[44] = in1[55] ^ in2[55];
    assign G[45] = in1[54] & in2[54];
    assign P[45] = in1[54] ^ in2[54];
    assign G[46] = in1[53] & in2[53];
    assign P[46] = in1[53] ^ in2[53];
    assign G[47] = in1[52] & in2[52];
    assign P[47] = in1[52] ^ in2[52];
    assign G[48] = in1[51] & in2[51];
    assign P[48] = in1[51] ^ in2[51];
    assign G[49] = in1[50] & in2[50];
    assign P[49] = in1[50] ^ in2[50];
    assign G[50] = in1[49] & in2[49];
    assign P[50] = in1[49] ^ in2[49];
    assign G[51] = in1[48] & in2[48];
    assign P[51] = in1[48] ^ in2[48];
    assign G[52] = in1[47] & in2[47];
    assign P[52] = in1[47] ^ in2[47];
    assign G[53] = in1[46] & in2[46];
    assign P[53] = in1[46] ^ in2[46];
    assign G[54] = in1[45] & in2[45];
    assign P[54] = in1[45] ^ in2[45];
    assign G[55] = in1[44] & in2[44];
    assign P[55] = in1[44] ^ in2[44];
    assign G[56] = in1[43] & in2[43];
    assign P[56] = in1[43] ^ in2[43];
    assign G[57] = in1[42] & in2[42];
    assign P[57] = in1[42] ^ in2[42];
    assign G[58] = in1[41] & in2[41];
    assign P[58] = in1[41] ^ in2[41];
    assign G[59] = in1[40] & in2[40];
    assign P[59] = in1[40] ^ in2[40];
    assign G[60] = in1[39] & in2[39];
    assign P[60] = in1[39] ^ in2[39];
    assign G[61] = in1[38] & in2[38];
    assign P[61] = in1[38] ^ in2[38];
    assign G[62] = in1[37] & in2[37];
    assign P[62] = in1[37] ^ in2[37];
    assign G[63] = in1[36] & in2[36];
    assign P[63] = in1[36] ^ in2[36];
    assign G[64] = in1[35] & in2[35];
    assign P[64] = in1[35] ^ in2[35];
    assign G[65] = in1[34] & in2[34];
    assign P[65] = in1[34] ^ in2[34];
    assign G[66] = in1[33] & in2[33];
    assign P[66] = in1[33] ^ in2[33];
    assign G[67] = in1[32] & in2[32];
    assign P[67] = in1[32] ^ in2[32];
    assign G[68] = in1[31] & in2[31];
    assign P[68] = in1[31] ^ in2[31];
    assign G[69] = in1[30] & in2[30];
    assign P[69] = in1[30] ^ in2[30];
    assign G[70] = in1[29] & in2[29];
    assign P[70] = in1[29] ^ in2[29];
    assign G[71] = in1[28] & in2[28];
    assign P[71] = in1[28] ^ in2[28];
    assign G[72] = in1[27] & in2[27];
    assign P[72] = in1[27] ^ in2[27];
    assign G[73] = in1[26] & in2[26];
    assign P[73] = in1[26] ^ in2[26];
    assign G[74] = in1[25] & in2[25];
    assign P[74] = in1[25] ^ in2[25];
    assign G[75] = in1[24] & in2[24];
    assign P[75] = in1[24] ^ in2[24];
    assign G[76] = in1[23] & in2[23];
    assign P[76] = in1[23] ^ in2[23];
    assign G[77] = in1[22] & in2[22];
    assign P[77] = in1[22] ^ in2[22];
    assign G[78] = in1[21] & in2[21];
    assign P[78] = in1[21] ^ in2[21];
    assign G[79] = in1[20] & in2[20];
    assign P[79] = in1[20] ^ in2[20];
    assign G[80] = in1[19] & in2[19];
    assign P[80] = in1[19] ^ in2[19];
    assign G[81] = in1[18] & in2[18];
    assign P[81] = in1[18] ^ in2[18];
    assign G[82] = in1[17] & in2[17];
    assign P[82] = in1[17] ^ in2[17];
    assign G[83] = in1[16] & in2[16];
    assign P[83] = in1[16] ^ in2[16];
    assign G[84] = in1[15] & in2[15];
    assign P[84] = in1[15] ^ in2[15];
    assign G[85] = in1[14] & in2[14];
    assign P[85] = in1[14] ^ in2[14];
    assign G[86] = in1[13] & in2[13];
    assign P[86] = in1[13] ^ in2[13];
    assign G[87] = in1[12] & in2[12];
    assign P[87] = in1[12] ^ in2[12];
    assign G[88] = in1[11] & in2[11];
    assign P[88] = in1[11] ^ in2[11];
    assign G[89] = in1[10] & in2[10];
    assign P[89] = in1[10] ^ in2[10];
    assign G[90] = in1[9] & in2[9];
    assign P[90] = in1[9] ^ in2[9];
    assign G[91] = in1[8] & in2[8];
    assign P[91] = in1[8] ^ in2[8];
    assign G[92] = in1[7] & in2[7];
    assign P[92] = in1[7] ^ in2[7];
    assign G[93] = in1[6] & in2[6];
    assign P[93] = in1[6] ^ in2[6];
    assign G[94] = in1[5] & in2[5];
    assign P[94] = in1[5] ^ in2[5];
    assign G[95] = in1[4] & in2[4];
    assign P[95] = in1[4] ^ in2[4];
    assign G[96] = in1[3] & in2[3];
    assign P[96] = in1[3] ^ in2[3];
    assign G[97] = in1[2] & in2[2];
    assign P[97] = in1[2] ^ in2[2];
    assign G[98] = in1[1] & in2[1];
    assign P[98] = in1[1] ^ in2[1];
    assign G[99] = in1[0] & in2[0];
    assign P[99] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign cout = G[99] | (P[99] & C[99]);
    assign sum = P ^ C;
endmodule

module CLA_99(output [98:0] sum, output cout, input [98:0] in1, input [98:0] in2);

    wire[98:0] G;
    wire[98:0] C;
    wire[98:0] P;

    assign G[0] = in1[98] & in2[98];
    assign P[0] = in1[98] ^ in2[98];
    assign G[1] = in1[97] & in2[97];
    assign P[1] = in1[97] ^ in2[97];
    assign G[2] = in1[96] & in2[96];
    assign P[2] = in1[96] ^ in2[96];
    assign G[3] = in1[95] & in2[95];
    assign P[3] = in1[95] ^ in2[95];
    assign G[4] = in1[94] & in2[94];
    assign P[4] = in1[94] ^ in2[94];
    assign G[5] = in1[93] & in2[93];
    assign P[5] = in1[93] ^ in2[93];
    assign G[6] = in1[92] & in2[92];
    assign P[6] = in1[92] ^ in2[92];
    assign G[7] = in1[91] & in2[91];
    assign P[7] = in1[91] ^ in2[91];
    assign G[8] = in1[90] & in2[90];
    assign P[8] = in1[90] ^ in2[90];
    assign G[9] = in1[89] & in2[89];
    assign P[9] = in1[89] ^ in2[89];
    assign G[10] = in1[88] & in2[88];
    assign P[10] = in1[88] ^ in2[88];
    assign G[11] = in1[87] & in2[87];
    assign P[11] = in1[87] ^ in2[87];
    assign G[12] = in1[86] & in2[86];
    assign P[12] = in1[86] ^ in2[86];
    assign G[13] = in1[85] & in2[85];
    assign P[13] = in1[85] ^ in2[85];
    assign G[14] = in1[84] & in2[84];
    assign P[14] = in1[84] ^ in2[84];
    assign G[15] = in1[83] & in2[83];
    assign P[15] = in1[83] ^ in2[83];
    assign G[16] = in1[82] & in2[82];
    assign P[16] = in1[82] ^ in2[82];
    assign G[17] = in1[81] & in2[81];
    assign P[17] = in1[81] ^ in2[81];
    assign G[18] = in1[80] & in2[80];
    assign P[18] = in1[80] ^ in2[80];
    assign G[19] = in1[79] & in2[79];
    assign P[19] = in1[79] ^ in2[79];
    assign G[20] = in1[78] & in2[78];
    assign P[20] = in1[78] ^ in2[78];
    assign G[21] = in1[77] & in2[77];
    assign P[21] = in1[77] ^ in2[77];
    assign G[22] = in1[76] & in2[76];
    assign P[22] = in1[76] ^ in2[76];
    assign G[23] = in1[75] & in2[75];
    assign P[23] = in1[75] ^ in2[75];
    assign G[24] = in1[74] & in2[74];
    assign P[24] = in1[74] ^ in2[74];
    assign G[25] = in1[73] & in2[73];
    assign P[25] = in1[73] ^ in2[73];
    assign G[26] = in1[72] & in2[72];
    assign P[26] = in1[72] ^ in2[72];
    assign G[27] = in1[71] & in2[71];
    assign P[27] = in1[71] ^ in2[71];
    assign G[28] = in1[70] & in2[70];
    assign P[28] = in1[70] ^ in2[70];
    assign G[29] = in1[69] & in2[69];
    assign P[29] = in1[69] ^ in2[69];
    assign G[30] = in1[68] & in2[68];
    assign P[30] = in1[68] ^ in2[68];
    assign G[31] = in1[67] & in2[67];
    assign P[31] = in1[67] ^ in2[67];
    assign G[32] = in1[66] & in2[66];
    assign P[32] = in1[66] ^ in2[66];
    assign G[33] = in1[65] & in2[65];
    assign P[33] = in1[65] ^ in2[65];
    assign G[34] = in1[64] & in2[64];
    assign P[34] = in1[64] ^ in2[64];
    assign G[35] = in1[63] & in2[63];
    assign P[35] = in1[63] ^ in2[63];
    assign G[36] = in1[62] & in2[62];
    assign P[36] = in1[62] ^ in2[62];
    assign G[37] = in1[61] & in2[61];
    assign P[37] = in1[61] ^ in2[61];
    assign G[38] = in1[60] & in2[60];
    assign P[38] = in1[60] ^ in2[60];
    assign G[39] = in1[59] & in2[59];
    assign P[39] = in1[59] ^ in2[59];
    assign G[40] = in1[58] & in2[58];
    assign P[40] = in1[58] ^ in2[58];
    assign G[41] = in1[57] & in2[57];
    assign P[41] = in1[57] ^ in2[57];
    assign G[42] = in1[56] & in2[56];
    assign P[42] = in1[56] ^ in2[56];
    assign G[43] = in1[55] & in2[55];
    assign P[43] = in1[55] ^ in2[55];
    assign G[44] = in1[54] & in2[54];
    assign P[44] = in1[54] ^ in2[54];
    assign G[45] = in1[53] & in2[53];
    assign P[45] = in1[53] ^ in2[53];
    assign G[46] = in1[52] & in2[52];
    assign P[46] = in1[52] ^ in2[52];
    assign G[47] = in1[51] & in2[51];
    assign P[47] = in1[51] ^ in2[51];
    assign G[48] = in1[50] & in2[50];
    assign P[48] = in1[50] ^ in2[50];
    assign G[49] = in1[49] & in2[49];
    assign P[49] = in1[49] ^ in2[49];
    assign G[50] = in1[48] & in2[48];
    assign P[50] = in1[48] ^ in2[48];
    assign G[51] = in1[47] & in2[47];
    assign P[51] = in1[47] ^ in2[47];
    assign G[52] = in1[46] & in2[46];
    assign P[52] = in1[46] ^ in2[46];
    assign G[53] = in1[45] & in2[45];
    assign P[53] = in1[45] ^ in2[45];
    assign G[54] = in1[44] & in2[44];
    assign P[54] = in1[44] ^ in2[44];
    assign G[55] = in1[43] & in2[43];
    assign P[55] = in1[43] ^ in2[43];
    assign G[56] = in1[42] & in2[42];
    assign P[56] = in1[42] ^ in2[42];
    assign G[57] = in1[41] & in2[41];
    assign P[57] = in1[41] ^ in2[41];
    assign G[58] = in1[40] & in2[40];
    assign P[58] = in1[40] ^ in2[40];
    assign G[59] = in1[39] & in2[39];
    assign P[59] = in1[39] ^ in2[39];
    assign G[60] = in1[38] & in2[38];
    assign P[60] = in1[38] ^ in2[38];
    assign G[61] = in1[37] & in2[37];
    assign P[61] = in1[37] ^ in2[37];
    assign G[62] = in1[36] & in2[36];
    assign P[62] = in1[36] ^ in2[36];
    assign G[63] = in1[35] & in2[35];
    assign P[63] = in1[35] ^ in2[35];
    assign G[64] = in1[34] & in2[34];
    assign P[64] = in1[34] ^ in2[34];
    assign G[65] = in1[33] & in2[33];
    assign P[65] = in1[33] ^ in2[33];
    assign G[66] = in1[32] & in2[32];
    assign P[66] = in1[32] ^ in2[32];
    assign G[67] = in1[31] & in2[31];
    assign P[67] = in1[31] ^ in2[31];
    assign G[68] = in1[30] & in2[30];
    assign P[68] = in1[30] ^ in2[30];
    assign G[69] = in1[29] & in2[29];
    assign P[69] = in1[29] ^ in2[29];
    assign G[70] = in1[28] & in2[28];
    assign P[70] = in1[28] ^ in2[28];
    assign G[71] = in1[27] & in2[27];
    assign P[71] = in1[27] ^ in2[27];
    assign G[72] = in1[26] & in2[26];
    assign P[72] = in1[26] ^ in2[26];
    assign G[73] = in1[25] & in2[25];
    assign P[73] = in1[25] ^ in2[25];
    assign G[74] = in1[24] & in2[24];
    assign P[74] = in1[24] ^ in2[24];
    assign G[75] = in1[23] & in2[23];
    assign P[75] = in1[23] ^ in2[23];
    assign G[76] = in1[22] & in2[22];
    assign P[76] = in1[22] ^ in2[22];
    assign G[77] = in1[21] & in2[21];
    assign P[77] = in1[21] ^ in2[21];
    assign G[78] = in1[20] & in2[20];
    assign P[78] = in1[20] ^ in2[20];
    assign G[79] = in1[19] & in2[19];
    assign P[79] = in1[19] ^ in2[19];
    assign G[80] = in1[18] & in2[18];
    assign P[80] = in1[18] ^ in2[18];
    assign G[81] = in1[17] & in2[17];
    assign P[81] = in1[17] ^ in2[17];
    assign G[82] = in1[16] & in2[16];
    assign P[82] = in1[16] ^ in2[16];
    assign G[83] = in1[15] & in2[15];
    assign P[83] = in1[15] ^ in2[15];
    assign G[84] = in1[14] & in2[14];
    assign P[84] = in1[14] ^ in2[14];
    assign G[85] = in1[13] & in2[13];
    assign P[85] = in1[13] ^ in2[13];
    assign G[86] = in1[12] & in2[12];
    assign P[86] = in1[12] ^ in2[12];
    assign G[87] = in1[11] & in2[11];
    assign P[87] = in1[11] ^ in2[11];
    assign G[88] = in1[10] & in2[10];
    assign P[88] = in1[10] ^ in2[10];
    assign G[89] = in1[9] & in2[9];
    assign P[89] = in1[9] ^ in2[9];
    assign G[90] = in1[8] & in2[8];
    assign P[90] = in1[8] ^ in2[8];
    assign G[91] = in1[7] & in2[7];
    assign P[91] = in1[7] ^ in2[7];
    assign G[92] = in1[6] & in2[6];
    assign P[92] = in1[6] ^ in2[6];
    assign G[93] = in1[5] & in2[5];
    assign P[93] = in1[5] ^ in2[5];
    assign G[94] = in1[4] & in2[4];
    assign P[94] = in1[4] ^ in2[4];
    assign G[95] = in1[3] & in2[3];
    assign P[95] = in1[3] ^ in2[3];
    assign G[96] = in1[2] & in2[2];
    assign P[96] = in1[2] ^ in2[2];
    assign G[97] = in1[1] & in2[1];
    assign P[97] = in1[1] ^ in2[1];
    assign G[98] = in1[0] & in2[0];
    assign P[98] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign cout = G[98] | (P[98] & C[98]);
    assign sum = P ^ C;
endmodule

module CLA_98(output [97:0] sum, output cout, input [97:0] in1, input [97:0] in2);

    wire[97:0] G;
    wire[97:0] C;
    wire[97:0] P;

    assign G[0] = in1[97] & in2[97];
    assign P[0] = in1[97] ^ in2[97];
    assign G[1] = in1[96] & in2[96];
    assign P[1] = in1[96] ^ in2[96];
    assign G[2] = in1[95] & in2[95];
    assign P[2] = in1[95] ^ in2[95];
    assign G[3] = in1[94] & in2[94];
    assign P[3] = in1[94] ^ in2[94];
    assign G[4] = in1[93] & in2[93];
    assign P[4] = in1[93] ^ in2[93];
    assign G[5] = in1[92] & in2[92];
    assign P[5] = in1[92] ^ in2[92];
    assign G[6] = in1[91] & in2[91];
    assign P[6] = in1[91] ^ in2[91];
    assign G[7] = in1[90] & in2[90];
    assign P[7] = in1[90] ^ in2[90];
    assign G[8] = in1[89] & in2[89];
    assign P[8] = in1[89] ^ in2[89];
    assign G[9] = in1[88] & in2[88];
    assign P[9] = in1[88] ^ in2[88];
    assign G[10] = in1[87] & in2[87];
    assign P[10] = in1[87] ^ in2[87];
    assign G[11] = in1[86] & in2[86];
    assign P[11] = in1[86] ^ in2[86];
    assign G[12] = in1[85] & in2[85];
    assign P[12] = in1[85] ^ in2[85];
    assign G[13] = in1[84] & in2[84];
    assign P[13] = in1[84] ^ in2[84];
    assign G[14] = in1[83] & in2[83];
    assign P[14] = in1[83] ^ in2[83];
    assign G[15] = in1[82] & in2[82];
    assign P[15] = in1[82] ^ in2[82];
    assign G[16] = in1[81] & in2[81];
    assign P[16] = in1[81] ^ in2[81];
    assign G[17] = in1[80] & in2[80];
    assign P[17] = in1[80] ^ in2[80];
    assign G[18] = in1[79] & in2[79];
    assign P[18] = in1[79] ^ in2[79];
    assign G[19] = in1[78] & in2[78];
    assign P[19] = in1[78] ^ in2[78];
    assign G[20] = in1[77] & in2[77];
    assign P[20] = in1[77] ^ in2[77];
    assign G[21] = in1[76] & in2[76];
    assign P[21] = in1[76] ^ in2[76];
    assign G[22] = in1[75] & in2[75];
    assign P[22] = in1[75] ^ in2[75];
    assign G[23] = in1[74] & in2[74];
    assign P[23] = in1[74] ^ in2[74];
    assign G[24] = in1[73] & in2[73];
    assign P[24] = in1[73] ^ in2[73];
    assign G[25] = in1[72] & in2[72];
    assign P[25] = in1[72] ^ in2[72];
    assign G[26] = in1[71] & in2[71];
    assign P[26] = in1[71] ^ in2[71];
    assign G[27] = in1[70] & in2[70];
    assign P[27] = in1[70] ^ in2[70];
    assign G[28] = in1[69] & in2[69];
    assign P[28] = in1[69] ^ in2[69];
    assign G[29] = in1[68] & in2[68];
    assign P[29] = in1[68] ^ in2[68];
    assign G[30] = in1[67] & in2[67];
    assign P[30] = in1[67] ^ in2[67];
    assign G[31] = in1[66] & in2[66];
    assign P[31] = in1[66] ^ in2[66];
    assign G[32] = in1[65] & in2[65];
    assign P[32] = in1[65] ^ in2[65];
    assign G[33] = in1[64] & in2[64];
    assign P[33] = in1[64] ^ in2[64];
    assign G[34] = in1[63] & in2[63];
    assign P[34] = in1[63] ^ in2[63];
    assign G[35] = in1[62] & in2[62];
    assign P[35] = in1[62] ^ in2[62];
    assign G[36] = in1[61] & in2[61];
    assign P[36] = in1[61] ^ in2[61];
    assign G[37] = in1[60] & in2[60];
    assign P[37] = in1[60] ^ in2[60];
    assign G[38] = in1[59] & in2[59];
    assign P[38] = in1[59] ^ in2[59];
    assign G[39] = in1[58] & in2[58];
    assign P[39] = in1[58] ^ in2[58];
    assign G[40] = in1[57] & in2[57];
    assign P[40] = in1[57] ^ in2[57];
    assign G[41] = in1[56] & in2[56];
    assign P[41] = in1[56] ^ in2[56];
    assign G[42] = in1[55] & in2[55];
    assign P[42] = in1[55] ^ in2[55];
    assign G[43] = in1[54] & in2[54];
    assign P[43] = in1[54] ^ in2[54];
    assign G[44] = in1[53] & in2[53];
    assign P[44] = in1[53] ^ in2[53];
    assign G[45] = in1[52] & in2[52];
    assign P[45] = in1[52] ^ in2[52];
    assign G[46] = in1[51] & in2[51];
    assign P[46] = in1[51] ^ in2[51];
    assign G[47] = in1[50] & in2[50];
    assign P[47] = in1[50] ^ in2[50];
    assign G[48] = in1[49] & in2[49];
    assign P[48] = in1[49] ^ in2[49];
    assign G[49] = in1[48] & in2[48];
    assign P[49] = in1[48] ^ in2[48];
    assign G[50] = in1[47] & in2[47];
    assign P[50] = in1[47] ^ in2[47];
    assign G[51] = in1[46] & in2[46];
    assign P[51] = in1[46] ^ in2[46];
    assign G[52] = in1[45] & in2[45];
    assign P[52] = in1[45] ^ in2[45];
    assign G[53] = in1[44] & in2[44];
    assign P[53] = in1[44] ^ in2[44];
    assign G[54] = in1[43] & in2[43];
    assign P[54] = in1[43] ^ in2[43];
    assign G[55] = in1[42] & in2[42];
    assign P[55] = in1[42] ^ in2[42];
    assign G[56] = in1[41] & in2[41];
    assign P[56] = in1[41] ^ in2[41];
    assign G[57] = in1[40] & in2[40];
    assign P[57] = in1[40] ^ in2[40];
    assign G[58] = in1[39] & in2[39];
    assign P[58] = in1[39] ^ in2[39];
    assign G[59] = in1[38] & in2[38];
    assign P[59] = in1[38] ^ in2[38];
    assign G[60] = in1[37] & in2[37];
    assign P[60] = in1[37] ^ in2[37];
    assign G[61] = in1[36] & in2[36];
    assign P[61] = in1[36] ^ in2[36];
    assign G[62] = in1[35] & in2[35];
    assign P[62] = in1[35] ^ in2[35];
    assign G[63] = in1[34] & in2[34];
    assign P[63] = in1[34] ^ in2[34];
    assign G[64] = in1[33] & in2[33];
    assign P[64] = in1[33] ^ in2[33];
    assign G[65] = in1[32] & in2[32];
    assign P[65] = in1[32] ^ in2[32];
    assign G[66] = in1[31] & in2[31];
    assign P[66] = in1[31] ^ in2[31];
    assign G[67] = in1[30] & in2[30];
    assign P[67] = in1[30] ^ in2[30];
    assign G[68] = in1[29] & in2[29];
    assign P[68] = in1[29] ^ in2[29];
    assign G[69] = in1[28] & in2[28];
    assign P[69] = in1[28] ^ in2[28];
    assign G[70] = in1[27] & in2[27];
    assign P[70] = in1[27] ^ in2[27];
    assign G[71] = in1[26] & in2[26];
    assign P[71] = in1[26] ^ in2[26];
    assign G[72] = in1[25] & in2[25];
    assign P[72] = in1[25] ^ in2[25];
    assign G[73] = in1[24] & in2[24];
    assign P[73] = in1[24] ^ in2[24];
    assign G[74] = in1[23] & in2[23];
    assign P[74] = in1[23] ^ in2[23];
    assign G[75] = in1[22] & in2[22];
    assign P[75] = in1[22] ^ in2[22];
    assign G[76] = in1[21] & in2[21];
    assign P[76] = in1[21] ^ in2[21];
    assign G[77] = in1[20] & in2[20];
    assign P[77] = in1[20] ^ in2[20];
    assign G[78] = in1[19] & in2[19];
    assign P[78] = in1[19] ^ in2[19];
    assign G[79] = in1[18] & in2[18];
    assign P[79] = in1[18] ^ in2[18];
    assign G[80] = in1[17] & in2[17];
    assign P[80] = in1[17] ^ in2[17];
    assign G[81] = in1[16] & in2[16];
    assign P[81] = in1[16] ^ in2[16];
    assign G[82] = in1[15] & in2[15];
    assign P[82] = in1[15] ^ in2[15];
    assign G[83] = in1[14] & in2[14];
    assign P[83] = in1[14] ^ in2[14];
    assign G[84] = in1[13] & in2[13];
    assign P[84] = in1[13] ^ in2[13];
    assign G[85] = in1[12] & in2[12];
    assign P[85] = in1[12] ^ in2[12];
    assign G[86] = in1[11] & in2[11];
    assign P[86] = in1[11] ^ in2[11];
    assign G[87] = in1[10] & in2[10];
    assign P[87] = in1[10] ^ in2[10];
    assign G[88] = in1[9] & in2[9];
    assign P[88] = in1[9] ^ in2[9];
    assign G[89] = in1[8] & in2[8];
    assign P[89] = in1[8] ^ in2[8];
    assign G[90] = in1[7] & in2[7];
    assign P[90] = in1[7] ^ in2[7];
    assign G[91] = in1[6] & in2[6];
    assign P[91] = in1[6] ^ in2[6];
    assign G[92] = in1[5] & in2[5];
    assign P[92] = in1[5] ^ in2[5];
    assign G[93] = in1[4] & in2[4];
    assign P[93] = in1[4] ^ in2[4];
    assign G[94] = in1[3] & in2[3];
    assign P[94] = in1[3] ^ in2[3];
    assign G[95] = in1[2] & in2[2];
    assign P[95] = in1[2] ^ in2[2];
    assign G[96] = in1[1] & in2[1];
    assign P[96] = in1[1] ^ in2[1];
    assign G[97] = in1[0] & in2[0];
    assign P[97] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign cout = G[97] | (P[97] & C[97]);
    assign sum = P ^ C;
endmodule

module CLA_97(output [96:0] sum, output cout, input [96:0] in1, input [96:0] in2);

    wire[96:0] G;
    wire[96:0] C;
    wire[96:0] P;

    assign G[0] = in1[96] & in2[96];
    assign P[0] = in1[96] ^ in2[96];
    assign G[1] = in1[95] & in2[95];
    assign P[1] = in1[95] ^ in2[95];
    assign G[2] = in1[94] & in2[94];
    assign P[2] = in1[94] ^ in2[94];
    assign G[3] = in1[93] & in2[93];
    assign P[3] = in1[93] ^ in2[93];
    assign G[4] = in1[92] & in2[92];
    assign P[4] = in1[92] ^ in2[92];
    assign G[5] = in1[91] & in2[91];
    assign P[5] = in1[91] ^ in2[91];
    assign G[6] = in1[90] & in2[90];
    assign P[6] = in1[90] ^ in2[90];
    assign G[7] = in1[89] & in2[89];
    assign P[7] = in1[89] ^ in2[89];
    assign G[8] = in1[88] & in2[88];
    assign P[8] = in1[88] ^ in2[88];
    assign G[9] = in1[87] & in2[87];
    assign P[9] = in1[87] ^ in2[87];
    assign G[10] = in1[86] & in2[86];
    assign P[10] = in1[86] ^ in2[86];
    assign G[11] = in1[85] & in2[85];
    assign P[11] = in1[85] ^ in2[85];
    assign G[12] = in1[84] & in2[84];
    assign P[12] = in1[84] ^ in2[84];
    assign G[13] = in1[83] & in2[83];
    assign P[13] = in1[83] ^ in2[83];
    assign G[14] = in1[82] & in2[82];
    assign P[14] = in1[82] ^ in2[82];
    assign G[15] = in1[81] & in2[81];
    assign P[15] = in1[81] ^ in2[81];
    assign G[16] = in1[80] & in2[80];
    assign P[16] = in1[80] ^ in2[80];
    assign G[17] = in1[79] & in2[79];
    assign P[17] = in1[79] ^ in2[79];
    assign G[18] = in1[78] & in2[78];
    assign P[18] = in1[78] ^ in2[78];
    assign G[19] = in1[77] & in2[77];
    assign P[19] = in1[77] ^ in2[77];
    assign G[20] = in1[76] & in2[76];
    assign P[20] = in1[76] ^ in2[76];
    assign G[21] = in1[75] & in2[75];
    assign P[21] = in1[75] ^ in2[75];
    assign G[22] = in1[74] & in2[74];
    assign P[22] = in1[74] ^ in2[74];
    assign G[23] = in1[73] & in2[73];
    assign P[23] = in1[73] ^ in2[73];
    assign G[24] = in1[72] & in2[72];
    assign P[24] = in1[72] ^ in2[72];
    assign G[25] = in1[71] & in2[71];
    assign P[25] = in1[71] ^ in2[71];
    assign G[26] = in1[70] & in2[70];
    assign P[26] = in1[70] ^ in2[70];
    assign G[27] = in1[69] & in2[69];
    assign P[27] = in1[69] ^ in2[69];
    assign G[28] = in1[68] & in2[68];
    assign P[28] = in1[68] ^ in2[68];
    assign G[29] = in1[67] & in2[67];
    assign P[29] = in1[67] ^ in2[67];
    assign G[30] = in1[66] & in2[66];
    assign P[30] = in1[66] ^ in2[66];
    assign G[31] = in1[65] & in2[65];
    assign P[31] = in1[65] ^ in2[65];
    assign G[32] = in1[64] & in2[64];
    assign P[32] = in1[64] ^ in2[64];
    assign G[33] = in1[63] & in2[63];
    assign P[33] = in1[63] ^ in2[63];
    assign G[34] = in1[62] & in2[62];
    assign P[34] = in1[62] ^ in2[62];
    assign G[35] = in1[61] & in2[61];
    assign P[35] = in1[61] ^ in2[61];
    assign G[36] = in1[60] & in2[60];
    assign P[36] = in1[60] ^ in2[60];
    assign G[37] = in1[59] & in2[59];
    assign P[37] = in1[59] ^ in2[59];
    assign G[38] = in1[58] & in2[58];
    assign P[38] = in1[58] ^ in2[58];
    assign G[39] = in1[57] & in2[57];
    assign P[39] = in1[57] ^ in2[57];
    assign G[40] = in1[56] & in2[56];
    assign P[40] = in1[56] ^ in2[56];
    assign G[41] = in1[55] & in2[55];
    assign P[41] = in1[55] ^ in2[55];
    assign G[42] = in1[54] & in2[54];
    assign P[42] = in1[54] ^ in2[54];
    assign G[43] = in1[53] & in2[53];
    assign P[43] = in1[53] ^ in2[53];
    assign G[44] = in1[52] & in2[52];
    assign P[44] = in1[52] ^ in2[52];
    assign G[45] = in1[51] & in2[51];
    assign P[45] = in1[51] ^ in2[51];
    assign G[46] = in1[50] & in2[50];
    assign P[46] = in1[50] ^ in2[50];
    assign G[47] = in1[49] & in2[49];
    assign P[47] = in1[49] ^ in2[49];
    assign G[48] = in1[48] & in2[48];
    assign P[48] = in1[48] ^ in2[48];
    assign G[49] = in1[47] & in2[47];
    assign P[49] = in1[47] ^ in2[47];
    assign G[50] = in1[46] & in2[46];
    assign P[50] = in1[46] ^ in2[46];
    assign G[51] = in1[45] & in2[45];
    assign P[51] = in1[45] ^ in2[45];
    assign G[52] = in1[44] & in2[44];
    assign P[52] = in1[44] ^ in2[44];
    assign G[53] = in1[43] & in2[43];
    assign P[53] = in1[43] ^ in2[43];
    assign G[54] = in1[42] & in2[42];
    assign P[54] = in1[42] ^ in2[42];
    assign G[55] = in1[41] & in2[41];
    assign P[55] = in1[41] ^ in2[41];
    assign G[56] = in1[40] & in2[40];
    assign P[56] = in1[40] ^ in2[40];
    assign G[57] = in1[39] & in2[39];
    assign P[57] = in1[39] ^ in2[39];
    assign G[58] = in1[38] & in2[38];
    assign P[58] = in1[38] ^ in2[38];
    assign G[59] = in1[37] & in2[37];
    assign P[59] = in1[37] ^ in2[37];
    assign G[60] = in1[36] & in2[36];
    assign P[60] = in1[36] ^ in2[36];
    assign G[61] = in1[35] & in2[35];
    assign P[61] = in1[35] ^ in2[35];
    assign G[62] = in1[34] & in2[34];
    assign P[62] = in1[34] ^ in2[34];
    assign G[63] = in1[33] & in2[33];
    assign P[63] = in1[33] ^ in2[33];
    assign G[64] = in1[32] & in2[32];
    assign P[64] = in1[32] ^ in2[32];
    assign G[65] = in1[31] & in2[31];
    assign P[65] = in1[31] ^ in2[31];
    assign G[66] = in1[30] & in2[30];
    assign P[66] = in1[30] ^ in2[30];
    assign G[67] = in1[29] & in2[29];
    assign P[67] = in1[29] ^ in2[29];
    assign G[68] = in1[28] & in2[28];
    assign P[68] = in1[28] ^ in2[28];
    assign G[69] = in1[27] & in2[27];
    assign P[69] = in1[27] ^ in2[27];
    assign G[70] = in1[26] & in2[26];
    assign P[70] = in1[26] ^ in2[26];
    assign G[71] = in1[25] & in2[25];
    assign P[71] = in1[25] ^ in2[25];
    assign G[72] = in1[24] & in2[24];
    assign P[72] = in1[24] ^ in2[24];
    assign G[73] = in1[23] & in2[23];
    assign P[73] = in1[23] ^ in2[23];
    assign G[74] = in1[22] & in2[22];
    assign P[74] = in1[22] ^ in2[22];
    assign G[75] = in1[21] & in2[21];
    assign P[75] = in1[21] ^ in2[21];
    assign G[76] = in1[20] & in2[20];
    assign P[76] = in1[20] ^ in2[20];
    assign G[77] = in1[19] & in2[19];
    assign P[77] = in1[19] ^ in2[19];
    assign G[78] = in1[18] & in2[18];
    assign P[78] = in1[18] ^ in2[18];
    assign G[79] = in1[17] & in2[17];
    assign P[79] = in1[17] ^ in2[17];
    assign G[80] = in1[16] & in2[16];
    assign P[80] = in1[16] ^ in2[16];
    assign G[81] = in1[15] & in2[15];
    assign P[81] = in1[15] ^ in2[15];
    assign G[82] = in1[14] & in2[14];
    assign P[82] = in1[14] ^ in2[14];
    assign G[83] = in1[13] & in2[13];
    assign P[83] = in1[13] ^ in2[13];
    assign G[84] = in1[12] & in2[12];
    assign P[84] = in1[12] ^ in2[12];
    assign G[85] = in1[11] & in2[11];
    assign P[85] = in1[11] ^ in2[11];
    assign G[86] = in1[10] & in2[10];
    assign P[86] = in1[10] ^ in2[10];
    assign G[87] = in1[9] & in2[9];
    assign P[87] = in1[9] ^ in2[9];
    assign G[88] = in1[8] & in2[8];
    assign P[88] = in1[8] ^ in2[8];
    assign G[89] = in1[7] & in2[7];
    assign P[89] = in1[7] ^ in2[7];
    assign G[90] = in1[6] & in2[6];
    assign P[90] = in1[6] ^ in2[6];
    assign G[91] = in1[5] & in2[5];
    assign P[91] = in1[5] ^ in2[5];
    assign G[92] = in1[4] & in2[4];
    assign P[92] = in1[4] ^ in2[4];
    assign G[93] = in1[3] & in2[3];
    assign P[93] = in1[3] ^ in2[3];
    assign G[94] = in1[2] & in2[2];
    assign P[94] = in1[2] ^ in2[2];
    assign G[95] = in1[1] & in2[1];
    assign P[95] = in1[1] ^ in2[1];
    assign G[96] = in1[0] & in2[0];
    assign P[96] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign cout = G[96] | (P[96] & C[96]);
    assign sum = P ^ C;
endmodule

module CLA_96(output [95:0] sum, output cout, input [95:0] in1, input [95:0] in2);

    wire[95:0] G;
    wire[95:0] C;
    wire[95:0] P;

    assign G[0] = in1[95] & in2[95];
    assign P[0] = in1[95] ^ in2[95];
    assign G[1] = in1[94] & in2[94];
    assign P[1] = in1[94] ^ in2[94];
    assign G[2] = in1[93] & in2[93];
    assign P[2] = in1[93] ^ in2[93];
    assign G[3] = in1[92] & in2[92];
    assign P[3] = in1[92] ^ in2[92];
    assign G[4] = in1[91] & in2[91];
    assign P[4] = in1[91] ^ in2[91];
    assign G[5] = in1[90] & in2[90];
    assign P[5] = in1[90] ^ in2[90];
    assign G[6] = in1[89] & in2[89];
    assign P[6] = in1[89] ^ in2[89];
    assign G[7] = in1[88] & in2[88];
    assign P[7] = in1[88] ^ in2[88];
    assign G[8] = in1[87] & in2[87];
    assign P[8] = in1[87] ^ in2[87];
    assign G[9] = in1[86] & in2[86];
    assign P[9] = in1[86] ^ in2[86];
    assign G[10] = in1[85] & in2[85];
    assign P[10] = in1[85] ^ in2[85];
    assign G[11] = in1[84] & in2[84];
    assign P[11] = in1[84] ^ in2[84];
    assign G[12] = in1[83] & in2[83];
    assign P[12] = in1[83] ^ in2[83];
    assign G[13] = in1[82] & in2[82];
    assign P[13] = in1[82] ^ in2[82];
    assign G[14] = in1[81] & in2[81];
    assign P[14] = in1[81] ^ in2[81];
    assign G[15] = in1[80] & in2[80];
    assign P[15] = in1[80] ^ in2[80];
    assign G[16] = in1[79] & in2[79];
    assign P[16] = in1[79] ^ in2[79];
    assign G[17] = in1[78] & in2[78];
    assign P[17] = in1[78] ^ in2[78];
    assign G[18] = in1[77] & in2[77];
    assign P[18] = in1[77] ^ in2[77];
    assign G[19] = in1[76] & in2[76];
    assign P[19] = in1[76] ^ in2[76];
    assign G[20] = in1[75] & in2[75];
    assign P[20] = in1[75] ^ in2[75];
    assign G[21] = in1[74] & in2[74];
    assign P[21] = in1[74] ^ in2[74];
    assign G[22] = in1[73] & in2[73];
    assign P[22] = in1[73] ^ in2[73];
    assign G[23] = in1[72] & in2[72];
    assign P[23] = in1[72] ^ in2[72];
    assign G[24] = in1[71] & in2[71];
    assign P[24] = in1[71] ^ in2[71];
    assign G[25] = in1[70] & in2[70];
    assign P[25] = in1[70] ^ in2[70];
    assign G[26] = in1[69] & in2[69];
    assign P[26] = in1[69] ^ in2[69];
    assign G[27] = in1[68] & in2[68];
    assign P[27] = in1[68] ^ in2[68];
    assign G[28] = in1[67] & in2[67];
    assign P[28] = in1[67] ^ in2[67];
    assign G[29] = in1[66] & in2[66];
    assign P[29] = in1[66] ^ in2[66];
    assign G[30] = in1[65] & in2[65];
    assign P[30] = in1[65] ^ in2[65];
    assign G[31] = in1[64] & in2[64];
    assign P[31] = in1[64] ^ in2[64];
    assign G[32] = in1[63] & in2[63];
    assign P[32] = in1[63] ^ in2[63];
    assign G[33] = in1[62] & in2[62];
    assign P[33] = in1[62] ^ in2[62];
    assign G[34] = in1[61] & in2[61];
    assign P[34] = in1[61] ^ in2[61];
    assign G[35] = in1[60] & in2[60];
    assign P[35] = in1[60] ^ in2[60];
    assign G[36] = in1[59] & in2[59];
    assign P[36] = in1[59] ^ in2[59];
    assign G[37] = in1[58] & in2[58];
    assign P[37] = in1[58] ^ in2[58];
    assign G[38] = in1[57] & in2[57];
    assign P[38] = in1[57] ^ in2[57];
    assign G[39] = in1[56] & in2[56];
    assign P[39] = in1[56] ^ in2[56];
    assign G[40] = in1[55] & in2[55];
    assign P[40] = in1[55] ^ in2[55];
    assign G[41] = in1[54] & in2[54];
    assign P[41] = in1[54] ^ in2[54];
    assign G[42] = in1[53] & in2[53];
    assign P[42] = in1[53] ^ in2[53];
    assign G[43] = in1[52] & in2[52];
    assign P[43] = in1[52] ^ in2[52];
    assign G[44] = in1[51] & in2[51];
    assign P[44] = in1[51] ^ in2[51];
    assign G[45] = in1[50] & in2[50];
    assign P[45] = in1[50] ^ in2[50];
    assign G[46] = in1[49] & in2[49];
    assign P[46] = in1[49] ^ in2[49];
    assign G[47] = in1[48] & in2[48];
    assign P[47] = in1[48] ^ in2[48];
    assign G[48] = in1[47] & in2[47];
    assign P[48] = in1[47] ^ in2[47];
    assign G[49] = in1[46] & in2[46];
    assign P[49] = in1[46] ^ in2[46];
    assign G[50] = in1[45] & in2[45];
    assign P[50] = in1[45] ^ in2[45];
    assign G[51] = in1[44] & in2[44];
    assign P[51] = in1[44] ^ in2[44];
    assign G[52] = in1[43] & in2[43];
    assign P[52] = in1[43] ^ in2[43];
    assign G[53] = in1[42] & in2[42];
    assign P[53] = in1[42] ^ in2[42];
    assign G[54] = in1[41] & in2[41];
    assign P[54] = in1[41] ^ in2[41];
    assign G[55] = in1[40] & in2[40];
    assign P[55] = in1[40] ^ in2[40];
    assign G[56] = in1[39] & in2[39];
    assign P[56] = in1[39] ^ in2[39];
    assign G[57] = in1[38] & in2[38];
    assign P[57] = in1[38] ^ in2[38];
    assign G[58] = in1[37] & in2[37];
    assign P[58] = in1[37] ^ in2[37];
    assign G[59] = in1[36] & in2[36];
    assign P[59] = in1[36] ^ in2[36];
    assign G[60] = in1[35] & in2[35];
    assign P[60] = in1[35] ^ in2[35];
    assign G[61] = in1[34] & in2[34];
    assign P[61] = in1[34] ^ in2[34];
    assign G[62] = in1[33] & in2[33];
    assign P[62] = in1[33] ^ in2[33];
    assign G[63] = in1[32] & in2[32];
    assign P[63] = in1[32] ^ in2[32];
    assign G[64] = in1[31] & in2[31];
    assign P[64] = in1[31] ^ in2[31];
    assign G[65] = in1[30] & in2[30];
    assign P[65] = in1[30] ^ in2[30];
    assign G[66] = in1[29] & in2[29];
    assign P[66] = in1[29] ^ in2[29];
    assign G[67] = in1[28] & in2[28];
    assign P[67] = in1[28] ^ in2[28];
    assign G[68] = in1[27] & in2[27];
    assign P[68] = in1[27] ^ in2[27];
    assign G[69] = in1[26] & in2[26];
    assign P[69] = in1[26] ^ in2[26];
    assign G[70] = in1[25] & in2[25];
    assign P[70] = in1[25] ^ in2[25];
    assign G[71] = in1[24] & in2[24];
    assign P[71] = in1[24] ^ in2[24];
    assign G[72] = in1[23] & in2[23];
    assign P[72] = in1[23] ^ in2[23];
    assign G[73] = in1[22] & in2[22];
    assign P[73] = in1[22] ^ in2[22];
    assign G[74] = in1[21] & in2[21];
    assign P[74] = in1[21] ^ in2[21];
    assign G[75] = in1[20] & in2[20];
    assign P[75] = in1[20] ^ in2[20];
    assign G[76] = in1[19] & in2[19];
    assign P[76] = in1[19] ^ in2[19];
    assign G[77] = in1[18] & in2[18];
    assign P[77] = in1[18] ^ in2[18];
    assign G[78] = in1[17] & in2[17];
    assign P[78] = in1[17] ^ in2[17];
    assign G[79] = in1[16] & in2[16];
    assign P[79] = in1[16] ^ in2[16];
    assign G[80] = in1[15] & in2[15];
    assign P[80] = in1[15] ^ in2[15];
    assign G[81] = in1[14] & in2[14];
    assign P[81] = in1[14] ^ in2[14];
    assign G[82] = in1[13] & in2[13];
    assign P[82] = in1[13] ^ in2[13];
    assign G[83] = in1[12] & in2[12];
    assign P[83] = in1[12] ^ in2[12];
    assign G[84] = in1[11] & in2[11];
    assign P[84] = in1[11] ^ in2[11];
    assign G[85] = in1[10] & in2[10];
    assign P[85] = in1[10] ^ in2[10];
    assign G[86] = in1[9] & in2[9];
    assign P[86] = in1[9] ^ in2[9];
    assign G[87] = in1[8] & in2[8];
    assign P[87] = in1[8] ^ in2[8];
    assign G[88] = in1[7] & in2[7];
    assign P[88] = in1[7] ^ in2[7];
    assign G[89] = in1[6] & in2[6];
    assign P[89] = in1[6] ^ in2[6];
    assign G[90] = in1[5] & in2[5];
    assign P[90] = in1[5] ^ in2[5];
    assign G[91] = in1[4] & in2[4];
    assign P[91] = in1[4] ^ in2[4];
    assign G[92] = in1[3] & in2[3];
    assign P[92] = in1[3] ^ in2[3];
    assign G[93] = in1[2] & in2[2];
    assign P[93] = in1[2] ^ in2[2];
    assign G[94] = in1[1] & in2[1];
    assign P[94] = in1[1] ^ in2[1];
    assign G[95] = in1[0] & in2[0];
    assign P[95] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign cout = G[95] | (P[95] & C[95]);
    assign sum = P ^ C;
endmodule

module CLA_95(output [94:0] sum, output cout, input [94:0] in1, input [94:0] in2);

    wire[94:0] G;
    wire[94:0] C;
    wire[94:0] P;

    assign G[0] = in1[94] & in2[94];
    assign P[0] = in1[94] ^ in2[94];
    assign G[1] = in1[93] & in2[93];
    assign P[1] = in1[93] ^ in2[93];
    assign G[2] = in1[92] & in2[92];
    assign P[2] = in1[92] ^ in2[92];
    assign G[3] = in1[91] & in2[91];
    assign P[3] = in1[91] ^ in2[91];
    assign G[4] = in1[90] & in2[90];
    assign P[4] = in1[90] ^ in2[90];
    assign G[5] = in1[89] & in2[89];
    assign P[5] = in1[89] ^ in2[89];
    assign G[6] = in1[88] & in2[88];
    assign P[6] = in1[88] ^ in2[88];
    assign G[7] = in1[87] & in2[87];
    assign P[7] = in1[87] ^ in2[87];
    assign G[8] = in1[86] & in2[86];
    assign P[8] = in1[86] ^ in2[86];
    assign G[9] = in1[85] & in2[85];
    assign P[9] = in1[85] ^ in2[85];
    assign G[10] = in1[84] & in2[84];
    assign P[10] = in1[84] ^ in2[84];
    assign G[11] = in1[83] & in2[83];
    assign P[11] = in1[83] ^ in2[83];
    assign G[12] = in1[82] & in2[82];
    assign P[12] = in1[82] ^ in2[82];
    assign G[13] = in1[81] & in2[81];
    assign P[13] = in1[81] ^ in2[81];
    assign G[14] = in1[80] & in2[80];
    assign P[14] = in1[80] ^ in2[80];
    assign G[15] = in1[79] & in2[79];
    assign P[15] = in1[79] ^ in2[79];
    assign G[16] = in1[78] & in2[78];
    assign P[16] = in1[78] ^ in2[78];
    assign G[17] = in1[77] & in2[77];
    assign P[17] = in1[77] ^ in2[77];
    assign G[18] = in1[76] & in2[76];
    assign P[18] = in1[76] ^ in2[76];
    assign G[19] = in1[75] & in2[75];
    assign P[19] = in1[75] ^ in2[75];
    assign G[20] = in1[74] & in2[74];
    assign P[20] = in1[74] ^ in2[74];
    assign G[21] = in1[73] & in2[73];
    assign P[21] = in1[73] ^ in2[73];
    assign G[22] = in1[72] & in2[72];
    assign P[22] = in1[72] ^ in2[72];
    assign G[23] = in1[71] & in2[71];
    assign P[23] = in1[71] ^ in2[71];
    assign G[24] = in1[70] & in2[70];
    assign P[24] = in1[70] ^ in2[70];
    assign G[25] = in1[69] & in2[69];
    assign P[25] = in1[69] ^ in2[69];
    assign G[26] = in1[68] & in2[68];
    assign P[26] = in1[68] ^ in2[68];
    assign G[27] = in1[67] & in2[67];
    assign P[27] = in1[67] ^ in2[67];
    assign G[28] = in1[66] & in2[66];
    assign P[28] = in1[66] ^ in2[66];
    assign G[29] = in1[65] & in2[65];
    assign P[29] = in1[65] ^ in2[65];
    assign G[30] = in1[64] & in2[64];
    assign P[30] = in1[64] ^ in2[64];
    assign G[31] = in1[63] & in2[63];
    assign P[31] = in1[63] ^ in2[63];
    assign G[32] = in1[62] & in2[62];
    assign P[32] = in1[62] ^ in2[62];
    assign G[33] = in1[61] & in2[61];
    assign P[33] = in1[61] ^ in2[61];
    assign G[34] = in1[60] & in2[60];
    assign P[34] = in1[60] ^ in2[60];
    assign G[35] = in1[59] & in2[59];
    assign P[35] = in1[59] ^ in2[59];
    assign G[36] = in1[58] & in2[58];
    assign P[36] = in1[58] ^ in2[58];
    assign G[37] = in1[57] & in2[57];
    assign P[37] = in1[57] ^ in2[57];
    assign G[38] = in1[56] & in2[56];
    assign P[38] = in1[56] ^ in2[56];
    assign G[39] = in1[55] & in2[55];
    assign P[39] = in1[55] ^ in2[55];
    assign G[40] = in1[54] & in2[54];
    assign P[40] = in1[54] ^ in2[54];
    assign G[41] = in1[53] & in2[53];
    assign P[41] = in1[53] ^ in2[53];
    assign G[42] = in1[52] & in2[52];
    assign P[42] = in1[52] ^ in2[52];
    assign G[43] = in1[51] & in2[51];
    assign P[43] = in1[51] ^ in2[51];
    assign G[44] = in1[50] & in2[50];
    assign P[44] = in1[50] ^ in2[50];
    assign G[45] = in1[49] & in2[49];
    assign P[45] = in1[49] ^ in2[49];
    assign G[46] = in1[48] & in2[48];
    assign P[46] = in1[48] ^ in2[48];
    assign G[47] = in1[47] & in2[47];
    assign P[47] = in1[47] ^ in2[47];
    assign G[48] = in1[46] & in2[46];
    assign P[48] = in1[46] ^ in2[46];
    assign G[49] = in1[45] & in2[45];
    assign P[49] = in1[45] ^ in2[45];
    assign G[50] = in1[44] & in2[44];
    assign P[50] = in1[44] ^ in2[44];
    assign G[51] = in1[43] & in2[43];
    assign P[51] = in1[43] ^ in2[43];
    assign G[52] = in1[42] & in2[42];
    assign P[52] = in1[42] ^ in2[42];
    assign G[53] = in1[41] & in2[41];
    assign P[53] = in1[41] ^ in2[41];
    assign G[54] = in1[40] & in2[40];
    assign P[54] = in1[40] ^ in2[40];
    assign G[55] = in1[39] & in2[39];
    assign P[55] = in1[39] ^ in2[39];
    assign G[56] = in1[38] & in2[38];
    assign P[56] = in1[38] ^ in2[38];
    assign G[57] = in1[37] & in2[37];
    assign P[57] = in1[37] ^ in2[37];
    assign G[58] = in1[36] & in2[36];
    assign P[58] = in1[36] ^ in2[36];
    assign G[59] = in1[35] & in2[35];
    assign P[59] = in1[35] ^ in2[35];
    assign G[60] = in1[34] & in2[34];
    assign P[60] = in1[34] ^ in2[34];
    assign G[61] = in1[33] & in2[33];
    assign P[61] = in1[33] ^ in2[33];
    assign G[62] = in1[32] & in2[32];
    assign P[62] = in1[32] ^ in2[32];
    assign G[63] = in1[31] & in2[31];
    assign P[63] = in1[31] ^ in2[31];
    assign G[64] = in1[30] & in2[30];
    assign P[64] = in1[30] ^ in2[30];
    assign G[65] = in1[29] & in2[29];
    assign P[65] = in1[29] ^ in2[29];
    assign G[66] = in1[28] & in2[28];
    assign P[66] = in1[28] ^ in2[28];
    assign G[67] = in1[27] & in2[27];
    assign P[67] = in1[27] ^ in2[27];
    assign G[68] = in1[26] & in2[26];
    assign P[68] = in1[26] ^ in2[26];
    assign G[69] = in1[25] & in2[25];
    assign P[69] = in1[25] ^ in2[25];
    assign G[70] = in1[24] & in2[24];
    assign P[70] = in1[24] ^ in2[24];
    assign G[71] = in1[23] & in2[23];
    assign P[71] = in1[23] ^ in2[23];
    assign G[72] = in1[22] & in2[22];
    assign P[72] = in1[22] ^ in2[22];
    assign G[73] = in1[21] & in2[21];
    assign P[73] = in1[21] ^ in2[21];
    assign G[74] = in1[20] & in2[20];
    assign P[74] = in1[20] ^ in2[20];
    assign G[75] = in1[19] & in2[19];
    assign P[75] = in1[19] ^ in2[19];
    assign G[76] = in1[18] & in2[18];
    assign P[76] = in1[18] ^ in2[18];
    assign G[77] = in1[17] & in2[17];
    assign P[77] = in1[17] ^ in2[17];
    assign G[78] = in1[16] & in2[16];
    assign P[78] = in1[16] ^ in2[16];
    assign G[79] = in1[15] & in2[15];
    assign P[79] = in1[15] ^ in2[15];
    assign G[80] = in1[14] & in2[14];
    assign P[80] = in1[14] ^ in2[14];
    assign G[81] = in1[13] & in2[13];
    assign P[81] = in1[13] ^ in2[13];
    assign G[82] = in1[12] & in2[12];
    assign P[82] = in1[12] ^ in2[12];
    assign G[83] = in1[11] & in2[11];
    assign P[83] = in1[11] ^ in2[11];
    assign G[84] = in1[10] & in2[10];
    assign P[84] = in1[10] ^ in2[10];
    assign G[85] = in1[9] & in2[9];
    assign P[85] = in1[9] ^ in2[9];
    assign G[86] = in1[8] & in2[8];
    assign P[86] = in1[8] ^ in2[8];
    assign G[87] = in1[7] & in2[7];
    assign P[87] = in1[7] ^ in2[7];
    assign G[88] = in1[6] & in2[6];
    assign P[88] = in1[6] ^ in2[6];
    assign G[89] = in1[5] & in2[5];
    assign P[89] = in1[5] ^ in2[5];
    assign G[90] = in1[4] & in2[4];
    assign P[90] = in1[4] ^ in2[4];
    assign G[91] = in1[3] & in2[3];
    assign P[91] = in1[3] ^ in2[3];
    assign G[92] = in1[2] & in2[2];
    assign P[92] = in1[2] ^ in2[2];
    assign G[93] = in1[1] & in2[1];
    assign P[93] = in1[1] ^ in2[1];
    assign G[94] = in1[0] & in2[0];
    assign P[94] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign cout = G[94] | (P[94] & C[94]);
    assign sum = P ^ C;
endmodule

module CLA_94(output [93:0] sum, output cout, input [93:0] in1, input [93:0] in2);

    wire[93:0] G;
    wire[93:0] C;
    wire[93:0] P;

    assign G[0] = in1[93] & in2[93];
    assign P[0] = in1[93] ^ in2[93];
    assign G[1] = in1[92] & in2[92];
    assign P[1] = in1[92] ^ in2[92];
    assign G[2] = in1[91] & in2[91];
    assign P[2] = in1[91] ^ in2[91];
    assign G[3] = in1[90] & in2[90];
    assign P[3] = in1[90] ^ in2[90];
    assign G[4] = in1[89] & in2[89];
    assign P[4] = in1[89] ^ in2[89];
    assign G[5] = in1[88] & in2[88];
    assign P[5] = in1[88] ^ in2[88];
    assign G[6] = in1[87] & in2[87];
    assign P[6] = in1[87] ^ in2[87];
    assign G[7] = in1[86] & in2[86];
    assign P[7] = in1[86] ^ in2[86];
    assign G[8] = in1[85] & in2[85];
    assign P[8] = in1[85] ^ in2[85];
    assign G[9] = in1[84] & in2[84];
    assign P[9] = in1[84] ^ in2[84];
    assign G[10] = in1[83] & in2[83];
    assign P[10] = in1[83] ^ in2[83];
    assign G[11] = in1[82] & in2[82];
    assign P[11] = in1[82] ^ in2[82];
    assign G[12] = in1[81] & in2[81];
    assign P[12] = in1[81] ^ in2[81];
    assign G[13] = in1[80] & in2[80];
    assign P[13] = in1[80] ^ in2[80];
    assign G[14] = in1[79] & in2[79];
    assign P[14] = in1[79] ^ in2[79];
    assign G[15] = in1[78] & in2[78];
    assign P[15] = in1[78] ^ in2[78];
    assign G[16] = in1[77] & in2[77];
    assign P[16] = in1[77] ^ in2[77];
    assign G[17] = in1[76] & in2[76];
    assign P[17] = in1[76] ^ in2[76];
    assign G[18] = in1[75] & in2[75];
    assign P[18] = in1[75] ^ in2[75];
    assign G[19] = in1[74] & in2[74];
    assign P[19] = in1[74] ^ in2[74];
    assign G[20] = in1[73] & in2[73];
    assign P[20] = in1[73] ^ in2[73];
    assign G[21] = in1[72] & in2[72];
    assign P[21] = in1[72] ^ in2[72];
    assign G[22] = in1[71] & in2[71];
    assign P[22] = in1[71] ^ in2[71];
    assign G[23] = in1[70] & in2[70];
    assign P[23] = in1[70] ^ in2[70];
    assign G[24] = in1[69] & in2[69];
    assign P[24] = in1[69] ^ in2[69];
    assign G[25] = in1[68] & in2[68];
    assign P[25] = in1[68] ^ in2[68];
    assign G[26] = in1[67] & in2[67];
    assign P[26] = in1[67] ^ in2[67];
    assign G[27] = in1[66] & in2[66];
    assign P[27] = in1[66] ^ in2[66];
    assign G[28] = in1[65] & in2[65];
    assign P[28] = in1[65] ^ in2[65];
    assign G[29] = in1[64] & in2[64];
    assign P[29] = in1[64] ^ in2[64];
    assign G[30] = in1[63] & in2[63];
    assign P[30] = in1[63] ^ in2[63];
    assign G[31] = in1[62] & in2[62];
    assign P[31] = in1[62] ^ in2[62];
    assign G[32] = in1[61] & in2[61];
    assign P[32] = in1[61] ^ in2[61];
    assign G[33] = in1[60] & in2[60];
    assign P[33] = in1[60] ^ in2[60];
    assign G[34] = in1[59] & in2[59];
    assign P[34] = in1[59] ^ in2[59];
    assign G[35] = in1[58] & in2[58];
    assign P[35] = in1[58] ^ in2[58];
    assign G[36] = in1[57] & in2[57];
    assign P[36] = in1[57] ^ in2[57];
    assign G[37] = in1[56] & in2[56];
    assign P[37] = in1[56] ^ in2[56];
    assign G[38] = in1[55] & in2[55];
    assign P[38] = in1[55] ^ in2[55];
    assign G[39] = in1[54] & in2[54];
    assign P[39] = in1[54] ^ in2[54];
    assign G[40] = in1[53] & in2[53];
    assign P[40] = in1[53] ^ in2[53];
    assign G[41] = in1[52] & in2[52];
    assign P[41] = in1[52] ^ in2[52];
    assign G[42] = in1[51] & in2[51];
    assign P[42] = in1[51] ^ in2[51];
    assign G[43] = in1[50] & in2[50];
    assign P[43] = in1[50] ^ in2[50];
    assign G[44] = in1[49] & in2[49];
    assign P[44] = in1[49] ^ in2[49];
    assign G[45] = in1[48] & in2[48];
    assign P[45] = in1[48] ^ in2[48];
    assign G[46] = in1[47] & in2[47];
    assign P[46] = in1[47] ^ in2[47];
    assign G[47] = in1[46] & in2[46];
    assign P[47] = in1[46] ^ in2[46];
    assign G[48] = in1[45] & in2[45];
    assign P[48] = in1[45] ^ in2[45];
    assign G[49] = in1[44] & in2[44];
    assign P[49] = in1[44] ^ in2[44];
    assign G[50] = in1[43] & in2[43];
    assign P[50] = in1[43] ^ in2[43];
    assign G[51] = in1[42] & in2[42];
    assign P[51] = in1[42] ^ in2[42];
    assign G[52] = in1[41] & in2[41];
    assign P[52] = in1[41] ^ in2[41];
    assign G[53] = in1[40] & in2[40];
    assign P[53] = in1[40] ^ in2[40];
    assign G[54] = in1[39] & in2[39];
    assign P[54] = in1[39] ^ in2[39];
    assign G[55] = in1[38] & in2[38];
    assign P[55] = in1[38] ^ in2[38];
    assign G[56] = in1[37] & in2[37];
    assign P[56] = in1[37] ^ in2[37];
    assign G[57] = in1[36] & in2[36];
    assign P[57] = in1[36] ^ in2[36];
    assign G[58] = in1[35] & in2[35];
    assign P[58] = in1[35] ^ in2[35];
    assign G[59] = in1[34] & in2[34];
    assign P[59] = in1[34] ^ in2[34];
    assign G[60] = in1[33] & in2[33];
    assign P[60] = in1[33] ^ in2[33];
    assign G[61] = in1[32] & in2[32];
    assign P[61] = in1[32] ^ in2[32];
    assign G[62] = in1[31] & in2[31];
    assign P[62] = in1[31] ^ in2[31];
    assign G[63] = in1[30] & in2[30];
    assign P[63] = in1[30] ^ in2[30];
    assign G[64] = in1[29] & in2[29];
    assign P[64] = in1[29] ^ in2[29];
    assign G[65] = in1[28] & in2[28];
    assign P[65] = in1[28] ^ in2[28];
    assign G[66] = in1[27] & in2[27];
    assign P[66] = in1[27] ^ in2[27];
    assign G[67] = in1[26] & in2[26];
    assign P[67] = in1[26] ^ in2[26];
    assign G[68] = in1[25] & in2[25];
    assign P[68] = in1[25] ^ in2[25];
    assign G[69] = in1[24] & in2[24];
    assign P[69] = in1[24] ^ in2[24];
    assign G[70] = in1[23] & in2[23];
    assign P[70] = in1[23] ^ in2[23];
    assign G[71] = in1[22] & in2[22];
    assign P[71] = in1[22] ^ in2[22];
    assign G[72] = in1[21] & in2[21];
    assign P[72] = in1[21] ^ in2[21];
    assign G[73] = in1[20] & in2[20];
    assign P[73] = in1[20] ^ in2[20];
    assign G[74] = in1[19] & in2[19];
    assign P[74] = in1[19] ^ in2[19];
    assign G[75] = in1[18] & in2[18];
    assign P[75] = in1[18] ^ in2[18];
    assign G[76] = in1[17] & in2[17];
    assign P[76] = in1[17] ^ in2[17];
    assign G[77] = in1[16] & in2[16];
    assign P[77] = in1[16] ^ in2[16];
    assign G[78] = in1[15] & in2[15];
    assign P[78] = in1[15] ^ in2[15];
    assign G[79] = in1[14] & in2[14];
    assign P[79] = in1[14] ^ in2[14];
    assign G[80] = in1[13] & in2[13];
    assign P[80] = in1[13] ^ in2[13];
    assign G[81] = in1[12] & in2[12];
    assign P[81] = in1[12] ^ in2[12];
    assign G[82] = in1[11] & in2[11];
    assign P[82] = in1[11] ^ in2[11];
    assign G[83] = in1[10] & in2[10];
    assign P[83] = in1[10] ^ in2[10];
    assign G[84] = in1[9] & in2[9];
    assign P[84] = in1[9] ^ in2[9];
    assign G[85] = in1[8] & in2[8];
    assign P[85] = in1[8] ^ in2[8];
    assign G[86] = in1[7] & in2[7];
    assign P[86] = in1[7] ^ in2[7];
    assign G[87] = in1[6] & in2[6];
    assign P[87] = in1[6] ^ in2[6];
    assign G[88] = in1[5] & in2[5];
    assign P[88] = in1[5] ^ in2[5];
    assign G[89] = in1[4] & in2[4];
    assign P[89] = in1[4] ^ in2[4];
    assign G[90] = in1[3] & in2[3];
    assign P[90] = in1[3] ^ in2[3];
    assign G[91] = in1[2] & in2[2];
    assign P[91] = in1[2] ^ in2[2];
    assign G[92] = in1[1] & in2[1];
    assign P[92] = in1[1] ^ in2[1];
    assign G[93] = in1[0] & in2[0];
    assign P[93] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign cout = G[93] | (P[93] & C[93]);
    assign sum = P ^ C;
endmodule

module CLA_93(output [92:0] sum, output cout, input [92:0] in1, input [92:0] in2);

    wire[92:0] G;
    wire[92:0] C;
    wire[92:0] P;

    assign G[0] = in1[92] & in2[92];
    assign P[0] = in1[92] ^ in2[92];
    assign G[1] = in1[91] & in2[91];
    assign P[1] = in1[91] ^ in2[91];
    assign G[2] = in1[90] & in2[90];
    assign P[2] = in1[90] ^ in2[90];
    assign G[3] = in1[89] & in2[89];
    assign P[3] = in1[89] ^ in2[89];
    assign G[4] = in1[88] & in2[88];
    assign P[4] = in1[88] ^ in2[88];
    assign G[5] = in1[87] & in2[87];
    assign P[5] = in1[87] ^ in2[87];
    assign G[6] = in1[86] & in2[86];
    assign P[6] = in1[86] ^ in2[86];
    assign G[7] = in1[85] & in2[85];
    assign P[7] = in1[85] ^ in2[85];
    assign G[8] = in1[84] & in2[84];
    assign P[8] = in1[84] ^ in2[84];
    assign G[9] = in1[83] & in2[83];
    assign P[9] = in1[83] ^ in2[83];
    assign G[10] = in1[82] & in2[82];
    assign P[10] = in1[82] ^ in2[82];
    assign G[11] = in1[81] & in2[81];
    assign P[11] = in1[81] ^ in2[81];
    assign G[12] = in1[80] & in2[80];
    assign P[12] = in1[80] ^ in2[80];
    assign G[13] = in1[79] & in2[79];
    assign P[13] = in1[79] ^ in2[79];
    assign G[14] = in1[78] & in2[78];
    assign P[14] = in1[78] ^ in2[78];
    assign G[15] = in1[77] & in2[77];
    assign P[15] = in1[77] ^ in2[77];
    assign G[16] = in1[76] & in2[76];
    assign P[16] = in1[76] ^ in2[76];
    assign G[17] = in1[75] & in2[75];
    assign P[17] = in1[75] ^ in2[75];
    assign G[18] = in1[74] & in2[74];
    assign P[18] = in1[74] ^ in2[74];
    assign G[19] = in1[73] & in2[73];
    assign P[19] = in1[73] ^ in2[73];
    assign G[20] = in1[72] & in2[72];
    assign P[20] = in1[72] ^ in2[72];
    assign G[21] = in1[71] & in2[71];
    assign P[21] = in1[71] ^ in2[71];
    assign G[22] = in1[70] & in2[70];
    assign P[22] = in1[70] ^ in2[70];
    assign G[23] = in1[69] & in2[69];
    assign P[23] = in1[69] ^ in2[69];
    assign G[24] = in1[68] & in2[68];
    assign P[24] = in1[68] ^ in2[68];
    assign G[25] = in1[67] & in2[67];
    assign P[25] = in1[67] ^ in2[67];
    assign G[26] = in1[66] & in2[66];
    assign P[26] = in1[66] ^ in2[66];
    assign G[27] = in1[65] & in2[65];
    assign P[27] = in1[65] ^ in2[65];
    assign G[28] = in1[64] & in2[64];
    assign P[28] = in1[64] ^ in2[64];
    assign G[29] = in1[63] & in2[63];
    assign P[29] = in1[63] ^ in2[63];
    assign G[30] = in1[62] & in2[62];
    assign P[30] = in1[62] ^ in2[62];
    assign G[31] = in1[61] & in2[61];
    assign P[31] = in1[61] ^ in2[61];
    assign G[32] = in1[60] & in2[60];
    assign P[32] = in1[60] ^ in2[60];
    assign G[33] = in1[59] & in2[59];
    assign P[33] = in1[59] ^ in2[59];
    assign G[34] = in1[58] & in2[58];
    assign P[34] = in1[58] ^ in2[58];
    assign G[35] = in1[57] & in2[57];
    assign P[35] = in1[57] ^ in2[57];
    assign G[36] = in1[56] & in2[56];
    assign P[36] = in1[56] ^ in2[56];
    assign G[37] = in1[55] & in2[55];
    assign P[37] = in1[55] ^ in2[55];
    assign G[38] = in1[54] & in2[54];
    assign P[38] = in1[54] ^ in2[54];
    assign G[39] = in1[53] & in2[53];
    assign P[39] = in1[53] ^ in2[53];
    assign G[40] = in1[52] & in2[52];
    assign P[40] = in1[52] ^ in2[52];
    assign G[41] = in1[51] & in2[51];
    assign P[41] = in1[51] ^ in2[51];
    assign G[42] = in1[50] & in2[50];
    assign P[42] = in1[50] ^ in2[50];
    assign G[43] = in1[49] & in2[49];
    assign P[43] = in1[49] ^ in2[49];
    assign G[44] = in1[48] & in2[48];
    assign P[44] = in1[48] ^ in2[48];
    assign G[45] = in1[47] & in2[47];
    assign P[45] = in1[47] ^ in2[47];
    assign G[46] = in1[46] & in2[46];
    assign P[46] = in1[46] ^ in2[46];
    assign G[47] = in1[45] & in2[45];
    assign P[47] = in1[45] ^ in2[45];
    assign G[48] = in1[44] & in2[44];
    assign P[48] = in1[44] ^ in2[44];
    assign G[49] = in1[43] & in2[43];
    assign P[49] = in1[43] ^ in2[43];
    assign G[50] = in1[42] & in2[42];
    assign P[50] = in1[42] ^ in2[42];
    assign G[51] = in1[41] & in2[41];
    assign P[51] = in1[41] ^ in2[41];
    assign G[52] = in1[40] & in2[40];
    assign P[52] = in1[40] ^ in2[40];
    assign G[53] = in1[39] & in2[39];
    assign P[53] = in1[39] ^ in2[39];
    assign G[54] = in1[38] & in2[38];
    assign P[54] = in1[38] ^ in2[38];
    assign G[55] = in1[37] & in2[37];
    assign P[55] = in1[37] ^ in2[37];
    assign G[56] = in1[36] & in2[36];
    assign P[56] = in1[36] ^ in2[36];
    assign G[57] = in1[35] & in2[35];
    assign P[57] = in1[35] ^ in2[35];
    assign G[58] = in1[34] & in2[34];
    assign P[58] = in1[34] ^ in2[34];
    assign G[59] = in1[33] & in2[33];
    assign P[59] = in1[33] ^ in2[33];
    assign G[60] = in1[32] & in2[32];
    assign P[60] = in1[32] ^ in2[32];
    assign G[61] = in1[31] & in2[31];
    assign P[61] = in1[31] ^ in2[31];
    assign G[62] = in1[30] & in2[30];
    assign P[62] = in1[30] ^ in2[30];
    assign G[63] = in1[29] & in2[29];
    assign P[63] = in1[29] ^ in2[29];
    assign G[64] = in1[28] & in2[28];
    assign P[64] = in1[28] ^ in2[28];
    assign G[65] = in1[27] & in2[27];
    assign P[65] = in1[27] ^ in2[27];
    assign G[66] = in1[26] & in2[26];
    assign P[66] = in1[26] ^ in2[26];
    assign G[67] = in1[25] & in2[25];
    assign P[67] = in1[25] ^ in2[25];
    assign G[68] = in1[24] & in2[24];
    assign P[68] = in1[24] ^ in2[24];
    assign G[69] = in1[23] & in2[23];
    assign P[69] = in1[23] ^ in2[23];
    assign G[70] = in1[22] & in2[22];
    assign P[70] = in1[22] ^ in2[22];
    assign G[71] = in1[21] & in2[21];
    assign P[71] = in1[21] ^ in2[21];
    assign G[72] = in1[20] & in2[20];
    assign P[72] = in1[20] ^ in2[20];
    assign G[73] = in1[19] & in2[19];
    assign P[73] = in1[19] ^ in2[19];
    assign G[74] = in1[18] & in2[18];
    assign P[74] = in1[18] ^ in2[18];
    assign G[75] = in1[17] & in2[17];
    assign P[75] = in1[17] ^ in2[17];
    assign G[76] = in1[16] & in2[16];
    assign P[76] = in1[16] ^ in2[16];
    assign G[77] = in1[15] & in2[15];
    assign P[77] = in1[15] ^ in2[15];
    assign G[78] = in1[14] & in2[14];
    assign P[78] = in1[14] ^ in2[14];
    assign G[79] = in1[13] & in2[13];
    assign P[79] = in1[13] ^ in2[13];
    assign G[80] = in1[12] & in2[12];
    assign P[80] = in1[12] ^ in2[12];
    assign G[81] = in1[11] & in2[11];
    assign P[81] = in1[11] ^ in2[11];
    assign G[82] = in1[10] & in2[10];
    assign P[82] = in1[10] ^ in2[10];
    assign G[83] = in1[9] & in2[9];
    assign P[83] = in1[9] ^ in2[9];
    assign G[84] = in1[8] & in2[8];
    assign P[84] = in1[8] ^ in2[8];
    assign G[85] = in1[7] & in2[7];
    assign P[85] = in1[7] ^ in2[7];
    assign G[86] = in1[6] & in2[6];
    assign P[86] = in1[6] ^ in2[6];
    assign G[87] = in1[5] & in2[5];
    assign P[87] = in1[5] ^ in2[5];
    assign G[88] = in1[4] & in2[4];
    assign P[88] = in1[4] ^ in2[4];
    assign G[89] = in1[3] & in2[3];
    assign P[89] = in1[3] ^ in2[3];
    assign G[90] = in1[2] & in2[2];
    assign P[90] = in1[2] ^ in2[2];
    assign G[91] = in1[1] & in2[1];
    assign P[91] = in1[1] ^ in2[1];
    assign G[92] = in1[0] & in2[0];
    assign P[92] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign cout = G[92] | (P[92] & C[92]);
    assign sum = P ^ C;
endmodule

module CLA_92(output [91:0] sum, output cout, input [91:0] in1, input [91:0] in2);

    wire[91:0] G;
    wire[91:0] C;
    wire[91:0] P;

    assign G[0] = in1[91] & in2[91];
    assign P[0] = in1[91] ^ in2[91];
    assign G[1] = in1[90] & in2[90];
    assign P[1] = in1[90] ^ in2[90];
    assign G[2] = in1[89] & in2[89];
    assign P[2] = in1[89] ^ in2[89];
    assign G[3] = in1[88] & in2[88];
    assign P[3] = in1[88] ^ in2[88];
    assign G[4] = in1[87] & in2[87];
    assign P[4] = in1[87] ^ in2[87];
    assign G[5] = in1[86] & in2[86];
    assign P[5] = in1[86] ^ in2[86];
    assign G[6] = in1[85] & in2[85];
    assign P[6] = in1[85] ^ in2[85];
    assign G[7] = in1[84] & in2[84];
    assign P[7] = in1[84] ^ in2[84];
    assign G[8] = in1[83] & in2[83];
    assign P[8] = in1[83] ^ in2[83];
    assign G[9] = in1[82] & in2[82];
    assign P[9] = in1[82] ^ in2[82];
    assign G[10] = in1[81] & in2[81];
    assign P[10] = in1[81] ^ in2[81];
    assign G[11] = in1[80] & in2[80];
    assign P[11] = in1[80] ^ in2[80];
    assign G[12] = in1[79] & in2[79];
    assign P[12] = in1[79] ^ in2[79];
    assign G[13] = in1[78] & in2[78];
    assign P[13] = in1[78] ^ in2[78];
    assign G[14] = in1[77] & in2[77];
    assign P[14] = in1[77] ^ in2[77];
    assign G[15] = in1[76] & in2[76];
    assign P[15] = in1[76] ^ in2[76];
    assign G[16] = in1[75] & in2[75];
    assign P[16] = in1[75] ^ in2[75];
    assign G[17] = in1[74] & in2[74];
    assign P[17] = in1[74] ^ in2[74];
    assign G[18] = in1[73] & in2[73];
    assign P[18] = in1[73] ^ in2[73];
    assign G[19] = in1[72] & in2[72];
    assign P[19] = in1[72] ^ in2[72];
    assign G[20] = in1[71] & in2[71];
    assign P[20] = in1[71] ^ in2[71];
    assign G[21] = in1[70] & in2[70];
    assign P[21] = in1[70] ^ in2[70];
    assign G[22] = in1[69] & in2[69];
    assign P[22] = in1[69] ^ in2[69];
    assign G[23] = in1[68] & in2[68];
    assign P[23] = in1[68] ^ in2[68];
    assign G[24] = in1[67] & in2[67];
    assign P[24] = in1[67] ^ in2[67];
    assign G[25] = in1[66] & in2[66];
    assign P[25] = in1[66] ^ in2[66];
    assign G[26] = in1[65] & in2[65];
    assign P[26] = in1[65] ^ in2[65];
    assign G[27] = in1[64] & in2[64];
    assign P[27] = in1[64] ^ in2[64];
    assign G[28] = in1[63] & in2[63];
    assign P[28] = in1[63] ^ in2[63];
    assign G[29] = in1[62] & in2[62];
    assign P[29] = in1[62] ^ in2[62];
    assign G[30] = in1[61] & in2[61];
    assign P[30] = in1[61] ^ in2[61];
    assign G[31] = in1[60] & in2[60];
    assign P[31] = in1[60] ^ in2[60];
    assign G[32] = in1[59] & in2[59];
    assign P[32] = in1[59] ^ in2[59];
    assign G[33] = in1[58] & in2[58];
    assign P[33] = in1[58] ^ in2[58];
    assign G[34] = in1[57] & in2[57];
    assign P[34] = in1[57] ^ in2[57];
    assign G[35] = in1[56] & in2[56];
    assign P[35] = in1[56] ^ in2[56];
    assign G[36] = in1[55] & in2[55];
    assign P[36] = in1[55] ^ in2[55];
    assign G[37] = in1[54] & in2[54];
    assign P[37] = in1[54] ^ in2[54];
    assign G[38] = in1[53] & in2[53];
    assign P[38] = in1[53] ^ in2[53];
    assign G[39] = in1[52] & in2[52];
    assign P[39] = in1[52] ^ in2[52];
    assign G[40] = in1[51] & in2[51];
    assign P[40] = in1[51] ^ in2[51];
    assign G[41] = in1[50] & in2[50];
    assign P[41] = in1[50] ^ in2[50];
    assign G[42] = in1[49] & in2[49];
    assign P[42] = in1[49] ^ in2[49];
    assign G[43] = in1[48] & in2[48];
    assign P[43] = in1[48] ^ in2[48];
    assign G[44] = in1[47] & in2[47];
    assign P[44] = in1[47] ^ in2[47];
    assign G[45] = in1[46] & in2[46];
    assign P[45] = in1[46] ^ in2[46];
    assign G[46] = in1[45] & in2[45];
    assign P[46] = in1[45] ^ in2[45];
    assign G[47] = in1[44] & in2[44];
    assign P[47] = in1[44] ^ in2[44];
    assign G[48] = in1[43] & in2[43];
    assign P[48] = in1[43] ^ in2[43];
    assign G[49] = in1[42] & in2[42];
    assign P[49] = in1[42] ^ in2[42];
    assign G[50] = in1[41] & in2[41];
    assign P[50] = in1[41] ^ in2[41];
    assign G[51] = in1[40] & in2[40];
    assign P[51] = in1[40] ^ in2[40];
    assign G[52] = in1[39] & in2[39];
    assign P[52] = in1[39] ^ in2[39];
    assign G[53] = in1[38] & in2[38];
    assign P[53] = in1[38] ^ in2[38];
    assign G[54] = in1[37] & in2[37];
    assign P[54] = in1[37] ^ in2[37];
    assign G[55] = in1[36] & in2[36];
    assign P[55] = in1[36] ^ in2[36];
    assign G[56] = in1[35] & in2[35];
    assign P[56] = in1[35] ^ in2[35];
    assign G[57] = in1[34] & in2[34];
    assign P[57] = in1[34] ^ in2[34];
    assign G[58] = in1[33] & in2[33];
    assign P[58] = in1[33] ^ in2[33];
    assign G[59] = in1[32] & in2[32];
    assign P[59] = in1[32] ^ in2[32];
    assign G[60] = in1[31] & in2[31];
    assign P[60] = in1[31] ^ in2[31];
    assign G[61] = in1[30] & in2[30];
    assign P[61] = in1[30] ^ in2[30];
    assign G[62] = in1[29] & in2[29];
    assign P[62] = in1[29] ^ in2[29];
    assign G[63] = in1[28] & in2[28];
    assign P[63] = in1[28] ^ in2[28];
    assign G[64] = in1[27] & in2[27];
    assign P[64] = in1[27] ^ in2[27];
    assign G[65] = in1[26] & in2[26];
    assign P[65] = in1[26] ^ in2[26];
    assign G[66] = in1[25] & in2[25];
    assign P[66] = in1[25] ^ in2[25];
    assign G[67] = in1[24] & in2[24];
    assign P[67] = in1[24] ^ in2[24];
    assign G[68] = in1[23] & in2[23];
    assign P[68] = in1[23] ^ in2[23];
    assign G[69] = in1[22] & in2[22];
    assign P[69] = in1[22] ^ in2[22];
    assign G[70] = in1[21] & in2[21];
    assign P[70] = in1[21] ^ in2[21];
    assign G[71] = in1[20] & in2[20];
    assign P[71] = in1[20] ^ in2[20];
    assign G[72] = in1[19] & in2[19];
    assign P[72] = in1[19] ^ in2[19];
    assign G[73] = in1[18] & in2[18];
    assign P[73] = in1[18] ^ in2[18];
    assign G[74] = in1[17] & in2[17];
    assign P[74] = in1[17] ^ in2[17];
    assign G[75] = in1[16] & in2[16];
    assign P[75] = in1[16] ^ in2[16];
    assign G[76] = in1[15] & in2[15];
    assign P[76] = in1[15] ^ in2[15];
    assign G[77] = in1[14] & in2[14];
    assign P[77] = in1[14] ^ in2[14];
    assign G[78] = in1[13] & in2[13];
    assign P[78] = in1[13] ^ in2[13];
    assign G[79] = in1[12] & in2[12];
    assign P[79] = in1[12] ^ in2[12];
    assign G[80] = in1[11] & in2[11];
    assign P[80] = in1[11] ^ in2[11];
    assign G[81] = in1[10] & in2[10];
    assign P[81] = in1[10] ^ in2[10];
    assign G[82] = in1[9] & in2[9];
    assign P[82] = in1[9] ^ in2[9];
    assign G[83] = in1[8] & in2[8];
    assign P[83] = in1[8] ^ in2[8];
    assign G[84] = in1[7] & in2[7];
    assign P[84] = in1[7] ^ in2[7];
    assign G[85] = in1[6] & in2[6];
    assign P[85] = in1[6] ^ in2[6];
    assign G[86] = in1[5] & in2[5];
    assign P[86] = in1[5] ^ in2[5];
    assign G[87] = in1[4] & in2[4];
    assign P[87] = in1[4] ^ in2[4];
    assign G[88] = in1[3] & in2[3];
    assign P[88] = in1[3] ^ in2[3];
    assign G[89] = in1[2] & in2[2];
    assign P[89] = in1[2] ^ in2[2];
    assign G[90] = in1[1] & in2[1];
    assign P[90] = in1[1] ^ in2[1];
    assign G[91] = in1[0] & in2[0];
    assign P[91] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign cout = G[91] | (P[91] & C[91]);
    assign sum = P ^ C;
endmodule

module CLA_91(output [90:0] sum, output cout, input [90:0] in1, input [90:0] in2);

    wire[90:0] G;
    wire[90:0] C;
    wire[90:0] P;

    assign G[0] = in1[90] & in2[90];
    assign P[0] = in1[90] ^ in2[90];
    assign G[1] = in1[89] & in2[89];
    assign P[1] = in1[89] ^ in2[89];
    assign G[2] = in1[88] & in2[88];
    assign P[2] = in1[88] ^ in2[88];
    assign G[3] = in1[87] & in2[87];
    assign P[3] = in1[87] ^ in2[87];
    assign G[4] = in1[86] & in2[86];
    assign P[4] = in1[86] ^ in2[86];
    assign G[5] = in1[85] & in2[85];
    assign P[5] = in1[85] ^ in2[85];
    assign G[6] = in1[84] & in2[84];
    assign P[6] = in1[84] ^ in2[84];
    assign G[7] = in1[83] & in2[83];
    assign P[7] = in1[83] ^ in2[83];
    assign G[8] = in1[82] & in2[82];
    assign P[8] = in1[82] ^ in2[82];
    assign G[9] = in1[81] & in2[81];
    assign P[9] = in1[81] ^ in2[81];
    assign G[10] = in1[80] & in2[80];
    assign P[10] = in1[80] ^ in2[80];
    assign G[11] = in1[79] & in2[79];
    assign P[11] = in1[79] ^ in2[79];
    assign G[12] = in1[78] & in2[78];
    assign P[12] = in1[78] ^ in2[78];
    assign G[13] = in1[77] & in2[77];
    assign P[13] = in1[77] ^ in2[77];
    assign G[14] = in1[76] & in2[76];
    assign P[14] = in1[76] ^ in2[76];
    assign G[15] = in1[75] & in2[75];
    assign P[15] = in1[75] ^ in2[75];
    assign G[16] = in1[74] & in2[74];
    assign P[16] = in1[74] ^ in2[74];
    assign G[17] = in1[73] & in2[73];
    assign P[17] = in1[73] ^ in2[73];
    assign G[18] = in1[72] & in2[72];
    assign P[18] = in1[72] ^ in2[72];
    assign G[19] = in1[71] & in2[71];
    assign P[19] = in1[71] ^ in2[71];
    assign G[20] = in1[70] & in2[70];
    assign P[20] = in1[70] ^ in2[70];
    assign G[21] = in1[69] & in2[69];
    assign P[21] = in1[69] ^ in2[69];
    assign G[22] = in1[68] & in2[68];
    assign P[22] = in1[68] ^ in2[68];
    assign G[23] = in1[67] & in2[67];
    assign P[23] = in1[67] ^ in2[67];
    assign G[24] = in1[66] & in2[66];
    assign P[24] = in1[66] ^ in2[66];
    assign G[25] = in1[65] & in2[65];
    assign P[25] = in1[65] ^ in2[65];
    assign G[26] = in1[64] & in2[64];
    assign P[26] = in1[64] ^ in2[64];
    assign G[27] = in1[63] & in2[63];
    assign P[27] = in1[63] ^ in2[63];
    assign G[28] = in1[62] & in2[62];
    assign P[28] = in1[62] ^ in2[62];
    assign G[29] = in1[61] & in2[61];
    assign P[29] = in1[61] ^ in2[61];
    assign G[30] = in1[60] & in2[60];
    assign P[30] = in1[60] ^ in2[60];
    assign G[31] = in1[59] & in2[59];
    assign P[31] = in1[59] ^ in2[59];
    assign G[32] = in1[58] & in2[58];
    assign P[32] = in1[58] ^ in2[58];
    assign G[33] = in1[57] & in2[57];
    assign P[33] = in1[57] ^ in2[57];
    assign G[34] = in1[56] & in2[56];
    assign P[34] = in1[56] ^ in2[56];
    assign G[35] = in1[55] & in2[55];
    assign P[35] = in1[55] ^ in2[55];
    assign G[36] = in1[54] & in2[54];
    assign P[36] = in1[54] ^ in2[54];
    assign G[37] = in1[53] & in2[53];
    assign P[37] = in1[53] ^ in2[53];
    assign G[38] = in1[52] & in2[52];
    assign P[38] = in1[52] ^ in2[52];
    assign G[39] = in1[51] & in2[51];
    assign P[39] = in1[51] ^ in2[51];
    assign G[40] = in1[50] & in2[50];
    assign P[40] = in1[50] ^ in2[50];
    assign G[41] = in1[49] & in2[49];
    assign P[41] = in1[49] ^ in2[49];
    assign G[42] = in1[48] & in2[48];
    assign P[42] = in1[48] ^ in2[48];
    assign G[43] = in1[47] & in2[47];
    assign P[43] = in1[47] ^ in2[47];
    assign G[44] = in1[46] & in2[46];
    assign P[44] = in1[46] ^ in2[46];
    assign G[45] = in1[45] & in2[45];
    assign P[45] = in1[45] ^ in2[45];
    assign G[46] = in1[44] & in2[44];
    assign P[46] = in1[44] ^ in2[44];
    assign G[47] = in1[43] & in2[43];
    assign P[47] = in1[43] ^ in2[43];
    assign G[48] = in1[42] & in2[42];
    assign P[48] = in1[42] ^ in2[42];
    assign G[49] = in1[41] & in2[41];
    assign P[49] = in1[41] ^ in2[41];
    assign G[50] = in1[40] & in2[40];
    assign P[50] = in1[40] ^ in2[40];
    assign G[51] = in1[39] & in2[39];
    assign P[51] = in1[39] ^ in2[39];
    assign G[52] = in1[38] & in2[38];
    assign P[52] = in1[38] ^ in2[38];
    assign G[53] = in1[37] & in2[37];
    assign P[53] = in1[37] ^ in2[37];
    assign G[54] = in1[36] & in2[36];
    assign P[54] = in1[36] ^ in2[36];
    assign G[55] = in1[35] & in2[35];
    assign P[55] = in1[35] ^ in2[35];
    assign G[56] = in1[34] & in2[34];
    assign P[56] = in1[34] ^ in2[34];
    assign G[57] = in1[33] & in2[33];
    assign P[57] = in1[33] ^ in2[33];
    assign G[58] = in1[32] & in2[32];
    assign P[58] = in1[32] ^ in2[32];
    assign G[59] = in1[31] & in2[31];
    assign P[59] = in1[31] ^ in2[31];
    assign G[60] = in1[30] & in2[30];
    assign P[60] = in1[30] ^ in2[30];
    assign G[61] = in1[29] & in2[29];
    assign P[61] = in1[29] ^ in2[29];
    assign G[62] = in1[28] & in2[28];
    assign P[62] = in1[28] ^ in2[28];
    assign G[63] = in1[27] & in2[27];
    assign P[63] = in1[27] ^ in2[27];
    assign G[64] = in1[26] & in2[26];
    assign P[64] = in1[26] ^ in2[26];
    assign G[65] = in1[25] & in2[25];
    assign P[65] = in1[25] ^ in2[25];
    assign G[66] = in1[24] & in2[24];
    assign P[66] = in1[24] ^ in2[24];
    assign G[67] = in1[23] & in2[23];
    assign P[67] = in1[23] ^ in2[23];
    assign G[68] = in1[22] & in2[22];
    assign P[68] = in1[22] ^ in2[22];
    assign G[69] = in1[21] & in2[21];
    assign P[69] = in1[21] ^ in2[21];
    assign G[70] = in1[20] & in2[20];
    assign P[70] = in1[20] ^ in2[20];
    assign G[71] = in1[19] & in2[19];
    assign P[71] = in1[19] ^ in2[19];
    assign G[72] = in1[18] & in2[18];
    assign P[72] = in1[18] ^ in2[18];
    assign G[73] = in1[17] & in2[17];
    assign P[73] = in1[17] ^ in2[17];
    assign G[74] = in1[16] & in2[16];
    assign P[74] = in1[16] ^ in2[16];
    assign G[75] = in1[15] & in2[15];
    assign P[75] = in1[15] ^ in2[15];
    assign G[76] = in1[14] & in2[14];
    assign P[76] = in1[14] ^ in2[14];
    assign G[77] = in1[13] & in2[13];
    assign P[77] = in1[13] ^ in2[13];
    assign G[78] = in1[12] & in2[12];
    assign P[78] = in1[12] ^ in2[12];
    assign G[79] = in1[11] & in2[11];
    assign P[79] = in1[11] ^ in2[11];
    assign G[80] = in1[10] & in2[10];
    assign P[80] = in1[10] ^ in2[10];
    assign G[81] = in1[9] & in2[9];
    assign P[81] = in1[9] ^ in2[9];
    assign G[82] = in1[8] & in2[8];
    assign P[82] = in1[8] ^ in2[8];
    assign G[83] = in1[7] & in2[7];
    assign P[83] = in1[7] ^ in2[7];
    assign G[84] = in1[6] & in2[6];
    assign P[84] = in1[6] ^ in2[6];
    assign G[85] = in1[5] & in2[5];
    assign P[85] = in1[5] ^ in2[5];
    assign G[86] = in1[4] & in2[4];
    assign P[86] = in1[4] ^ in2[4];
    assign G[87] = in1[3] & in2[3];
    assign P[87] = in1[3] ^ in2[3];
    assign G[88] = in1[2] & in2[2];
    assign P[88] = in1[2] ^ in2[2];
    assign G[89] = in1[1] & in2[1];
    assign P[89] = in1[1] ^ in2[1];
    assign G[90] = in1[0] & in2[0];
    assign P[90] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign cout = G[90] | (P[90] & C[90]);
    assign sum = P ^ C;
endmodule

module CLA_90(output [89:0] sum, output cout, input [89:0] in1, input [89:0] in2);

    wire[89:0] G;
    wire[89:0] C;
    wire[89:0] P;

    assign G[0] = in1[89] & in2[89];
    assign P[0] = in1[89] ^ in2[89];
    assign G[1] = in1[88] & in2[88];
    assign P[1] = in1[88] ^ in2[88];
    assign G[2] = in1[87] & in2[87];
    assign P[2] = in1[87] ^ in2[87];
    assign G[3] = in1[86] & in2[86];
    assign P[3] = in1[86] ^ in2[86];
    assign G[4] = in1[85] & in2[85];
    assign P[4] = in1[85] ^ in2[85];
    assign G[5] = in1[84] & in2[84];
    assign P[5] = in1[84] ^ in2[84];
    assign G[6] = in1[83] & in2[83];
    assign P[6] = in1[83] ^ in2[83];
    assign G[7] = in1[82] & in2[82];
    assign P[7] = in1[82] ^ in2[82];
    assign G[8] = in1[81] & in2[81];
    assign P[8] = in1[81] ^ in2[81];
    assign G[9] = in1[80] & in2[80];
    assign P[9] = in1[80] ^ in2[80];
    assign G[10] = in1[79] & in2[79];
    assign P[10] = in1[79] ^ in2[79];
    assign G[11] = in1[78] & in2[78];
    assign P[11] = in1[78] ^ in2[78];
    assign G[12] = in1[77] & in2[77];
    assign P[12] = in1[77] ^ in2[77];
    assign G[13] = in1[76] & in2[76];
    assign P[13] = in1[76] ^ in2[76];
    assign G[14] = in1[75] & in2[75];
    assign P[14] = in1[75] ^ in2[75];
    assign G[15] = in1[74] & in2[74];
    assign P[15] = in1[74] ^ in2[74];
    assign G[16] = in1[73] & in2[73];
    assign P[16] = in1[73] ^ in2[73];
    assign G[17] = in1[72] & in2[72];
    assign P[17] = in1[72] ^ in2[72];
    assign G[18] = in1[71] & in2[71];
    assign P[18] = in1[71] ^ in2[71];
    assign G[19] = in1[70] & in2[70];
    assign P[19] = in1[70] ^ in2[70];
    assign G[20] = in1[69] & in2[69];
    assign P[20] = in1[69] ^ in2[69];
    assign G[21] = in1[68] & in2[68];
    assign P[21] = in1[68] ^ in2[68];
    assign G[22] = in1[67] & in2[67];
    assign P[22] = in1[67] ^ in2[67];
    assign G[23] = in1[66] & in2[66];
    assign P[23] = in1[66] ^ in2[66];
    assign G[24] = in1[65] & in2[65];
    assign P[24] = in1[65] ^ in2[65];
    assign G[25] = in1[64] & in2[64];
    assign P[25] = in1[64] ^ in2[64];
    assign G[26] = in1[63] & in2[63];
    assign P[26] = in1[63] ^ in2[63];
    assign G[27] = in1[62] & in2[62];
    assign P[27] = in1[62] ^ in2[62];
    assign G[28] = in1[61] & in2[61];
    assign P[28] = in1[61] ^ in2[61];
    assign G[29] = in1[60] & in2[60];
    assign P[29] = in1[60] ^ in2[60];
    assign G[30] = in1[59] & in2[59];
    assign P[30] = in1[59] ^ in2[59];
    assign G[31] = in1[58] & in2[58];
    assign P[31] = in1[58] ^ in2[58];
    assign G[32] = in1[57] & in2[57];
    assign P[32] = in1[57] ^ in2[57];
    assign G[33] = in1[56] & in2[56];
    assign P[33] = in1[56] ^ in2[56];
    assign G[34] = in1[55] & in2[55];
    assign P[34] = in1[55] ^ in2[55];
    assign G[35] = in1[54] & in2[54];
    assign P[35] = in1[54] ^ in2[54];
    assign G[36] = in1[53] & in2[53];
    assign P[36] = in1[53] ^ in2[53];
    assign G[37] = in1[52] & in2[52];
    assign P[37] = in1[52] ^ in2[52];
    assign G[38] = in1[51] & in2[51];
    assign P[38] = in1[51] ^ in2[51];
    assign G[39] = in1[50] & in2[50];
    assign P[39] = in1[50] ^ in2[50];
    assign G[40] = in1[49] & in2[49];
    assign P[40] = in1[49] ^ in2[49];
    assign G[41] = in1[48] & in2[48];
    assign P[41] = in1[48] ^ in2[48];
    assign G[42] = in1[47] & in2[47];
    assign P[42] = in1[47] ^ in2[47];
    assign G[43] = in1[46] & in2[46];
    assign P[43] = in1[46] ^ in2[46];
    assign G[44] = in1[45] & in2[45];
    assign P[44] = in1[45] ^ in2[45];
    assign G[45] = in1[44] & in2[44];
    assign P[45] = in1[44] ^ in2[44];
    assign G[46] = in1[43] & in2[43];
    assign P[46] = in1[43] ^ in2[43];
    assign G[47] = in1[42] & in2[42];
    assign P[47] = in1[42] ^ in2[42];
    assign G[48] = in1[41] & in2[41];
    assign P[48] = in1[41] ^ in2[41];
    assign G[49] = in1[40] & in2[40];
    assign P[49] = in1[40] ^ in2[40];
    assign G[50] = in1[39] & in2[39];
    assign P[50] = in1[39] ^ in2[39];
    assign G[51] = in1[38] & in2[38];
    assign P[51] = in1[38] ^ in2[38];
    assign G[52] = in1[37] & in2[37];
    assign P[52] = in1[37] ^ in2[37];
    assign G[53] = in1[36] & in2[36];
    assign P[53] = in1[36] ^ in2[36];
    assign G[54] = in1[35] & in2[35];
    assign P[54] = in1[35] ^ in2[35];
    assign G[55] = in1[34] & in2[34];
    assign P[55] = in1[34] ^ in2[34];
    assign G[56] = in1[33] & in2[33];
    assign P[56] = in1[33] ^ in2[33];
    assign G[57] = in1[32] & in2[32];
    assign P[57] = in1[32] ^ in2[32];
    assign G[58] = in1[31] & in2[31];
    assign P[58] = in1[31] ^ in2[31];
    assign G[59] = in1[30] & in2[30];
    assign P[59] = in1[30] ^ in2[30];
    assign G[60] = in1[29] & in2[29];
    assign P[60] = in1[29] ^ in2[29];
    assign G[61] = in1[28] & in2[28];
    assign P[61] = in1[28] ^ in2[28];
    assign G[62] = in1[27] & in2[27];
    assign P[62] = in1[27] ^ in2[27];
    assign G[63] = in1[26] & in2[26];
    assign P[63] = in1[26] ^ in2[26];
    assign G[64] = in1[25] & in2[25];
    assign P[64] = in1[25] ^ in2[25];
    assign G[65] = in1[24] & in2[24];
    assign P[65] = in1[24] ^ in2[24];
    assign G[66] = in1[23] & in2[23];
    assign P[66] = in1[23] ^ in2[23];
    assign G[67] = in1[22] & in2[22];
    assign P[67] = in1[22] ^ in2[22];
    assign G[68] = in1[21] & in2[21];
    assign P[68] = in1[21] ^ in2[21];
    assign G[69] = in1[20] & in2[20];
    assign P[69] = in1[20] ^ in2[20];
    assign G[70] = in1[19] & in2[19];
    assign P[70] = in1[19] ^ in2[19];
    assign G[71] = in1[18] & in2[18];
    assign P[71] = in1[18] ^ in2[18];
    assign G[72] = in1[17] & in2[17];
    assign P[72] = in1[17] ^ in2[17];
    assign G[73] = in1[16] & in2[16];
    assign P[73] = in1[16] ^ in2[16];
    assign G[74] = in1[15] & in2[15];
    assign P[74] = in1[15] ^ in2[15];
    assign G[75] = in1[14] & in2[14];
    assign P[75] = in1[14] ^ in2[14];
    assign G[76] = in1[13] & in2[13];
    assign P[76] = in1[13] ^ in2[13];
    assign G[77] = in1[12] & in2[12];
    assign P[77] = in1[12] ^ in2[12];
    assign G[78] = in1[11] & in2[11];
    assign P[78] = in1[11] ^ in2[11];
    assign G[79] = in1[10] & in2[10];
    assign P[79] = in1[10] ^ in2[10];
    assign G[80] = in1[9] & in2[9];
    assign P[80] = in1[9] ^ in2[9];
    assign G[81] = in1[8] & in2[8];
    assign P[81] = in1[8] ^ in2[8];
    assign G[82] = in1[7] & in2[7];
    assign P[82] = in1[7] ^ in2[7];
    assign G[83] = in1[6] & in2[6];
    assign P[83] = in1[6] ^ in2[6];
    assign G[84] = in1[5] & in2[5];
    assign P[84] = in1[5] ^ in2[5];
    assign G[85] = in1[4] & in2[4];
    assign P[85] = in1[4] ^ in2[4];
    assign G[86] = in1[3] & in2[3];
    assign P[86] = in1[3] ^ in2[3];
    assign G[87] = in1[2] & in2[2];
    assign P[87] = in1[2] ^ in2[2];
    assign G[88] = in1[1] & in2[1];
    assign P[88] = in1[1] ^ in2[1];
    assign G[89] = in1[0] & in2[0];
    assign P[89] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign cout = G[89] | (P[89] & C[89]);
    assign sum = P ^ C;
endmodule

module CLA_89(output [88:0] sum, output cout, input [88:0] in1, input [88:0] in2);

    wire[88:0] G;
    wire[88:0] C;
    wire[88:0] P;

    assign G[0] = in1[88] & in2[88];
    assign P[0] = in1[88] ^ in2[88];
    assign G[1] = in1[87] & in2[87];
    assign P[1] = in1[87] ^ in2[87];
    assign G[2] = in1[86] & in2[86];
    assign P[2] = in1[86] ^ in2[86];
    assign G[3] = in1[85] & in2[85];
    assign P[3] = in1[85] ^ in2[85];
    assign G[4] = in1[84] & in2[84];
    assign P[4] = in1[84] ^ in2[84];
    assign G[5] = in1[83] & in2[83];
    assign P[5] = in1[83] ^ in2[83];
    assign G[6] = in1[82] & in2[82];
    assign P[6] = in1[82] ^ in2[82];
    assign G[7] = in1[81] & in2[81];
    assign P[7] = in1[81] ^ in2[81];
    assign G[8] = in1[80] & in2[80];
    assign P[8] = in1[80] ^ in2[80];
    assign G[9] = in1[79] & in2[79];
    assign P[9] = in1[79] ^ in2[79];
    assign G[10] = in1[78] & in2[78];
    assign P[10] = in1[78] ^ in2[78];
    assign G[11] = in1[77] & in2[77];
    assign P[11] = in1[77] ^ in2[77];
    assign G[12] = in1[76] & in2[76];
    assign P[12] = in1[76] ^ in2[76];
    assign G[13] = in1[75] & in2[75];
    assign P[13] = in1[75] ^ in2[75];
    assign G[14] = in1[74] & in2[74];
    assign P[14] = in1[74] ^ in2[74];
    assign G[15] = in1[73] & in2[73];
    assign P[15] = in1[73] ^ in2[73];
    assign G[16] = in1[72] & in2[72];
    assign P[16] = in1[72] ^ in2[72];
    assign G[17] = in1[71] & in2[71];
    assign P[17] = in1[71] ^ in2[71];
    assign G[18] = in1[70] & in2[70];
    assign P[18] = in1[70] ^ in2[70];
    assign G[19] = in1[69] & in2[69];
    assign P[19] = in1[69] ^ in2[69];
    assign G[20] = in1[68] & in2[68];
    assign P[20] = in1[68] ^ in2[68];
    assign G[21] = in1[67] & in2[67];
    assign P[21] = in1[67] ^ in2[67];
    assign G[22] = in1[66] & in2[66];
    assign P[22] = in1[66] ^ in2[66];
    assign G[23] = in1[65] & in2[65];
    assign P[23] = in1[65] ^ in2[65];
    assign G[24] = in1[64] & in2[64];
    assign P[24] = in1[64] ^ in2[64];
    assign G[25] = in1[63] & in2[63];
    assign P[25] = in1[63] ^ in2[63];
    assign G[26] = in1[62] & in2[62];
    assign P[26] = in1[62] ^ in2[62];
    assign G[27] = in1[61] & in2[61];
    assign P[27] = in1[61] ^ in2[61];
    assign G[28] = in1[60] & in2[60];
    assign P[28] = in1[60] ^ in2[60];
    assign G[29] = in1[59] & in2[59];
    assign P[29] = in1[59] ^ in2[59];
    assign G[30] = in1[58] & in2[58];
    assign P[30] = in1[58] ^ in2[58];
    assign G[31] = in1[57] & in2[57];
    assign P[31] = in1[57] ^ in2[57];
    assign G[32] = in1[56] & in2[56];
    assign P[32] = in1[56] ^ in2[56];
    assign G[33] = in1[55] & in2[55];
    assign P[33] = in1[55] ^ in2[55];
    assign G[34] = in1[54] & in2[54];
    assign P[34] = in1[54] ^ in2[54];
    assign G[35] = in1[53] & in2[53];
    assign P[35] = in1[53] ^ in2[53];
    assign G[36] = in1[52] & in2[52];
    assign P[36] = in1[52] ^ in2[52];
    assign G[37] = in1[51] & in2[51];
    assign P[37] = in1[51] ^ in2[51];
    assign G[38] = in1[50] & in2[50];
    assign P[38] = in1[50] ^ in2[50];
    assign G[39] = in1[49] & in2[49];
    assign P[39] = in1[49] ^ in2[49];
    assign G[40] = in1[48] & in2[48];
    assign P[40] = in1[48] ^ in2[48];
    assign G[41] = in1[47] & in2[47];
    assign P[41] = in1[47] ^ in2[47];
    assign G[42] = in1[46] & in2[46];
    assign P[42] = in1[46] ^ in2[46];
    assign G[43] = in1[45] & in2[45];
    assign P[43] = in1[45] ^ in2[45];
    assign G[44] = in1[44] & in2[44];
    assign P[44] = in1[44] ^ in2[44];
    assign G[45] = in1[43] & in2[43];
    assign P[45] = in1[43] ^ in2[43];
    assign G[46] = in1[42] & in2[42];
    assign P[46] = in1[42] ^ in2[42];
    assign G[47] = in1[41] & in2[41];
    assign P[47] = in1[41] ^ in2[41];
    assign G[48] = in1[40] & in2[40];
    assign P[48] = in1[40] ^ in2[40];
    assign G[49] = in1[39] & in2[39];
    assign P[49] = in1[39] ^ in2[39];
    assign G[50] = in1[38] & in2[38];
    assign P[50] = in1[38] ^ in2[38];
    assign G[51] = in1[37] & in2[37];
    assign P[51] = in1[37] ^ in2[37];
    assign G[52] = in1[36] & in2[36];
    assign P[52] = in1[36] ^ in2[36];
    assign G[53] = in1[35] & in2[35];
    assign P[53] = in1[35] ^ in2[35];
    assign G[54] = in1[34] & in2[34];
    assign P[54] = in1[34] ^ in2[34];
    assign G[55] = in1[33] & in2[33];
    assign P[55] = in1[33] ^ in2[33];
    assign G[56] = in1[32] & in2[32];
    assign P[56] = in1[32] ^ in2[32];
    assign G[57] = in1[31] & in2[31];
    assign P[57] = in1[31] ^ in2[31];
    assign G[58] = in1[30] & in2[30];
    assign P[58] = in1[30] ^ in2[30];
    assign G[59] = in1[29] & in2[29];
    assign P[59] = in1[29] ^ in2[29];
    assign G[60] = in1[28] & in2[28];
    assign P[60] = in1[28] ^ in2[28];
    assign G[61] = in1[27] & in2[27];
    assign P[61] = in1[27] ^ in2[27];
    assign G[62] = in1[26] & in2[26];
    assign P[62] = in1[26] ^ in2[26];
    assign G[63] = in1[25] & in2[25];
    assign P[63] = in1[25] ^ in2[25];
    assign G[64] = in1[24] & in2[24];
    assign P[64] = in1[24] ^ in2[24];
    assign G[65] = in1[23] & in2[23];
    assign P[65] = in1[23] ^ in2[23];
    assign G[66] = in1[22] & in2[22];
    assign P[66] = in1[22] ^ in2[22];
    assign G[67] = in1[21] & in2[21];
    assign P[67] = in1[21] ^ in2[21];
    assign G[68] = in1[20] & in2[20];
    assign P[68] = in1[20] ^ in2[20];
    assign G[69] = in1[19] & in2[19];
    assign P[69] = in1[19] ^ in2[19];
    assign G[70] = in1[18] & in2[18];
    assign P[70] = in1[18] ^ in2[18];
    assign G[71] = in1[17] & in2[17];
    assign P[71] = in1[17] ^ in2[17];
    assign G[72] = in1[16] & in2[16];
    assign P[72] = in1[16] ^ in2[16];
    assign G[73] = in1[15] & in2[15];
    assign P[73] = in1[15] ^ in2[15];
    assign G[74] = in1[14] & in2[14];
    assign P[74] = in1[14] ^ in2[14];
    assign G[75] = in1[13] & in2[13];
    assign P[75] = in1[13] ^ in2[13];
    assign G[76] = in1[12] & in2[12];
    assign P[76] = in1[12] ^ in2[12];
    assign G[77] = in1[11] & in2[11];
    assign P[77] = in1[11] ^ in2[11];
    assign G[78] = in1[10] & in2[10];
    assign P[78] = in1[10] ^ in2[10];
    assign G[79] = in1[9] & in2[9];
    assign P[79] = in1[9] ^ in2[9];
    assign G[80] = in1[8] & in2[8];
    assign P[80] = in1[8] ^ in2[8];
    assign G[81] = in1[7] & in2[7];
    assign P[81] = in1[7] ^ in2[7];
    assign G[82] = in1[6] & in2[6];
    assign P[82] = in1[6] ^ in2[6];
    assign G[83] = in1[5] & in2[5];
    assign P[83] = in1[5] ^ in2[5];
    assign G[84] = in1[4] & in2[4];
    assign P[84] = in1[4] ^ in2[4];
    assign G[85] = in1[3] & in2[3];
    assign P[85] = in1[3] ^ in2[3];
    assign G[86] = in1[2] & in2[2];
    assign P[86] = in1[2] ^ in2[2];
    assign G[87] = in1[1] & in2[1];
    assign P[87] = in1[1] ^ in2[1];
    assign G[88] = in1[0] & in2[0];
    assign P[88] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign cout = G[88] | (P[88] & C[88]);
    assign sum = P ^ C;
endmodule

module CLA_88(output [87:0] sum, output cout, input [87:0] in1, input [87:0] in2);

    wire[87:0] G;
    wire[87:0] C;
    wire[87:0] P;

    assign G[0] = in1[87] & in2[87];
    assign P[0] = in1[87] ^ in2[87];
    assign G[1] = in1[86] & in2[86];
    assign P[1] = in1[86] ^ in2[86];
    assign G[2] = in1[85] & in2[85];
    assign P[2] = in1[85] ^ in2[85];
    assign G[3] = in1[84] & in2[84];
    assign P[3] = in1[84] ^ in2[84];
    assign G[4] = in1[83] & in2[83];
    assign P[4] = in1[83] ^ in2[83];
    assign G[5] = in1[82] & in2[82];
    assign P[5] = in1[82] ^ in2[82];
    assign G[6] = in1[81] & in2[81];
    assign P[6] = in1[81] ^ in2[81];
    assign G[7] = in1[80] & in2[80];
    assign P[7] = in1[80] ^ in2[80];
    assign G[8] = in1[79] & in2[79];
    assign P[8] = in1[79] ^ in2[79];
    assign G[9] = in1[78] & in2[78];
    assign P[9] = in1[78] ^ in2[78];
    assign G[10] = in1[77] & in2[77];
    assign P[10] = in1[77] ^ in2[77];
    assign G[11] = in1[76] & in2[76];
    assign P[11] = in1[76] ^ in2[76];
    assign G[12] = in1[75] & in2[75];
    assign P[12] = in1[75] ^ in2[75];
    assign G[13] = in1[74] & in2[74];
    assign P[13] = in1[74] ^ in2[74];
    assign G[14] = in1[73] & in2[73];
    assign P[14] = in1[73] ^ in2[73];
    assign G[15] = in1[72] & in2[72];
    assign P[15] = in1[72] ^ in2[72];
    assign G[16] = in1[71] & in2[71];
    assign P[16] = in1[71] ^ in2[71];
    assign G[17] = in1[70] & in2[70];
    assign P[17] = in1[70] ^ in2[70];
    assign G[18] = in1[69] & in2[69];
    assign P[18] = in1[69] ^ in2[69];
    assign G[19] = in1[68] & in2[68];
    assign P[19] = in1[68] ^ in2[68];
    assign G[20] = in1[67] & in2[67];
    assign P[20] = in1[67] ^ in2[67];
    assign G[21] = in1[66] & in2[66];
    assign P[21] = in1[66] ^ in2[66];
    assign G[22] = in1[65] & in2[65];
    assign P[22] = in1[65] ^ in2[65];
    assign G[23] = in1[64] & in2[64];
    assign P[23] = in1[64] ^ in2[64];
    assign G[24] = in1[63] & in2[63];
    assign P[24] = in1[63] ^ in2[63];
    assign G[25] = in1[62] & in2[62];
    assign P[25] = in1[62] ^ in2[62];
    assign G[26] = in1[61] & in2[61];
    assign P[26] = in1[61] ^ in2[61];
    assign G[27] = in1[60] & in2[60];
    assign P[27] = in1[60] ^ in2[60];
    assign G[28] = in1[59] & in2[59];
    assign P[28] = in1[59] ^ in2[59];
    assign G[29] = in1[58] & in2[58];
    assign P[29] = in1[58] ^ in2[58];
    assign G[30] = in1[57] & in2[57];
    assign P[30] = in1[57] ^ in2[57];
    assign G[31] = in1[56] & in2[56];
    assign P[31] = in1[56] ^ in2[56];
    assign G[32] = in1[55] & in2[55];
    assign P[32] = in1[55] ^ in2[55];
    assign G[33] = in1[54] & in2[54];
    assign P[33] = in1[54] ^ in2[54];
    assign G[34] = in1[53] & in2[53];
    assign P[34] = in1[53] ^ in2[53];
    assign G[35] = in1[52] & in2[52];
    assign P[35] = in1[52] ^ in2[52];
    assign G[36] = in1[51] & in2[51];
    assign P[36] = in1[51] ^ in2[51];
    assign G[37] = in1[50] & in2[50];
    assign P[37] = in1[50] ^ in2[50];
    assign G[38] = in1[49] & in2[49];
    assign P[38] = in1[49] ^ in2[49];
    assign G[39] = in1[48] & in2[48];
    assign P[39] = in1[48] ^ in2[48];
    assign G[40] = in1[47] & in2[47];
    assign P[40] = in1[47] ^ in2[47];
    assign G[41] = in1[46] & in2[46];
    assign P[41] = in1[46] ^ in2[46];
    assign G[42] = in1[45] & in2[45];
    assign P[42] = in1[45] ^ in2[45];
    assign G[43] = in1[44] & in2[44];
    assign P[43] = in1[44] ^ in2[44];
    assign G[44] = in1[43] & in2[43];
    assign P[44] = in1[43] ^ in2[43];
    assign G[45] = in1[42] & in2[42];
    assign P[45] = in1[42] ^ in2[42];
    assign G[46] = in1[41] & in2[41];
    assign P[46] = in1[41] ^ in2[41];
    assign G[47] = in1[40] & in2[40];
    assign P[47] = in1[40] ^ in2[40];
    assign G[48] = in1[39] & in2[39];
    assign P[48] = in1[39] ^ in2[39];
    assign G[49] = in1[38] & in2[38];
    assign P[49] = in1[38] ^ in2[38];
    assign G[50] = in1[37] & in2[37];
    assign P[50] = in1[37] ^ in2[37];
    assign G[51] = in1[36] & in2[36];
    assign P[51] = in1[36] ^ in2[36];
    assign G[52] = in1[35] & in2[35];
    assign P[52] = in1[35] ^ in2[35];
    assign G[53] = in1[34] & in2[34];
    assign P[53] = in1[34] ^ in2[34];
    assign G[54] = in1[33] & in2[33];
    assign P[54] = in1[33] ^ in2[33];
    assign G[55] = in1[32] & in2[32];
    assign P[55] = in1[32] ^ in2[32];
    assign G[56] = in1[31] & in2[31];
    assign P[56] = in1[31] ^ in2[31];
    assign G[57] = in1[30] & in2[30];
    assign P[57] = in1[30] ^ in2[30];
    assign G[58] = in1[29] & in2[29];
    assign P[58] = in1[29] ^ in2[29];
    assign G[59] = in1[28] & in2[28];
    assign P[59] = in1[28] ^ in2[28];
    assign G[60] = in1[27] & in2[27];
    assign P[60] = in1[27] ^ in2[27];
    assign G[61] = in1[26] & in2[26];
    assign P[61] = in1[26] ^ in2[26];
    assign G[62] = in1[25] & in2[25];
    assign P[62] = in1[25] ^ in2[25];
    assign G[63] = in1[24] & in2[24];
    assign P[63] = in1[24] ^ in2[24];
    assign G[64] = in1[23] & in2[23];
    assign P[64] = in1[23] ^ in2[23];
    assign G[65] = in1[22] & in2[22];
    assign P[65] = in1[22] ^ in2[22];
    assign G[66] = in1[21] & in2[21];
    assign P[66] = in1[21] ^ in2[21];
    assign G[67] = in1[20] & in2[20];
    assign P[67] = in1[20] ^ in2[20];
    assign G[68] = in1[19] & in2[19];
    assign P[68] = in1[19] ^ in2[19];
    assign G[69] = in1[18] & in2[18];
    assign P[69] = in1[18] ^ in2[18];
    assign G[70] = in1[17] & in2[17];
    assign P[70] = in1[17] ^ in2[17];
    assign G[71] = in1[16] & in2[16];
    assign P[71] = in1[16] ^ in2[16];
    assign G[72] = in1[15] & in2[15];
    assign P[72] = in1[15] ^ in2[15];
    assign G[73] = in1[14] & in2[14];
    assign P[73] = in1[14] ^ in2[14];
    assign G[74] = in1[13] & in2[13];
    assign P[74] = in1[13] ^ in2[13];
    assign G[75] = in1[12] & in2[12];
    assign P[75] = in1[12] ^ in2[12];
    assign G[76] = in1[11] & in2[11];
    assign P[76] = in1[11] ^ in2[11];
    assign G[77] = in1[10] & in2[10];
    assign P[77] = in1[10] ^ in2[10];
    assign G[78] = in1[9] & in2[9];
    assign P[78] = in1[9] ^ in2[9];
    assign G[79] = in1[8] & in2[8];
    assign P[79] = in1[8] ^ in2[8];
    assign G[80] = in1[7] & in2[7];
    assign P[80] = in1[7] ^ in2[7];
    assign G[81] = in1[6] & in2[6];
    assign P[81] = in1[6] ^ in2[6];
    assign G[82] = in1[5] & in2[5];
    assign P[82] = in1[5] ^ in2[5];
    assign G[83] = in1[4] & in2[4];
    assign P[83] = in1[4] ^ in2[4];
    assign G[84] = in1[3] & in2[3];
    assign P[84] = in1[3] ^ in2[3];
    assign G[85] = in1[2] & in2[2];
    assign P[85] = in1[2] ^ in2[2];
    assign G[86] = in1[1] & in2[1];
    assign P[86] = in1[1] ^ in2[1];
    assign G[87] = in1[0] & in2[0];
    assign P[87] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign cout = G[87] | (P[87] & C[87]);
    assign sum = P ^ C;
endmodule

module CLA_87(output [86:0] sum, output cout, input [86:0] in1, input [86:0] in2);

    wire[86:0] G;
    wire[86:0] C;
    wire[86:0] P;

    assign G[0] = in1[86] & in2[86];
    assign P[0] = in1[86] ^ in2[86];
    assign G[1] = in1[85] & in2[85];
    assign P[1] = in1[85] ^ in2[85];
    assign G[2] = in1[84] & in2[84];
    assign P[2] = in1[84] ^ in2[84];
    assign G[3] = in1[83] & in2[83];
    assign P[3] = in1[83] ^ in2[83];
    assign G[4] = in1[82] & in2[82];
    assign P[4] = in1[82] ^ in2[82];
    assign G[5] = in1[81] & in2[81];
    assign P[5] = in1[81] ^ in2[81];
    assign G[6] = in1[80] & in2[80];
    assign P[6] = in1[80] ^ in2[80];
    assign G[7] = in1[79] & in2[79];
    assign P[7] = in1[79] ^ in2[79];
    assign G[8] = in1[78] & in2[78];
    assign P[8] = in1[78] ^ in2[78];
    assign G[9] = in1[77] & in2[77];
    assign P[9] = in1[77] ^ in2[77];
    assign G[10] = in1[76] & in2[76];
    assign P[10] = in1[76] ^ in2[76];
    assign G[11] = in1[75] & in2[75];
    assign P[11] = in1[75] ^ in2[75];
    assign G[12] = in1[74] & in2[74];
    assign P[12] = in1[74] ^ in2[74];
    assign G[13] = in1[73] & in2[73];
    assign P[13] = in1[73] ^ in2[73];
    assign G[14] = in1[72] & in2[72];
    assign P[14] = in1[72] ^ in2[72];
    assign G[15] = in1[71] & in2[71];
    assign P[15] = in1[71] ^ in2[71];
    assign G[16] = in1[70] & in2[70];
    assign P[16] = in1[70] ^ in2[70];
    assign G[17] = in1[69] & in2[69];
    assign P[17] = in1[69] ^ in2[69];
    assign G[18] = in1[68] & in2[68];
    assign P[18] = in1[68] ^ in2[68];
    assign G[19] = in1[67] & in2[67];
    assign P[19] = in1[67] ^ in2[67];
    assign G[20] = in1[66] & in2[66];
    assign P[20] = in1[66] ^ in2[66];
    assign G[21] = in1[65] & in2[65];
    assign P[21] = in1[65] ^ in2[65];
    assign G[22] = in1[64] & in2[64];
    assign P[22] = in1[64] ^ in2[64];
    assign G[23] = in1[63] & in2[63];
    assign P[23] = in1[63] ^ in2[63];
    assign G[24] = in1[62] & in2[62];
    assign P[24] = in1[62] ^ in2[62];
    assign G[25] = in1[61] & in2[61];
    assign P[25] = in1[61] ^ in2[61];
    assign G[26] = in1[60] & in2[60];
    assign P[26] = in1[60] ^ in2[60];
    assign G[27] = in1[59] & in2[59];
    assign P[27] = in1[59] ^ in2[59];
    assign G[28] = in1[58] & in2[58];
    assign P[28] = in1[58] ^ in2[58];
    assign G[29] = in1[57] & in2[57];
    assign P[29] = in1[57] ^ in2[57];
    assign G[30] = in1[56] & in2[56];
    assign P[30] = in1[56] ^ in2[56];
    assign G[31] = in1[55] & in2[55];
    assign P[31] = in1[55] ^ in2[55];
    assign G[32] = in1[54] & in2[54];
    assign P[32] = in1[54] ^ in2[54];
    assign G[33] = in1[53] & in2[53];
    assign P[33] = in1[53] ^ in2[53];
    assign G[34] = in1[52] & in2[52];
    assign P[34] = in1[52] ^ in2[52];
    assign G[35] = in1[51] & in2[51];
    assign P[35] = in1[51] ^ in2[51];
    assign G[36] = in1[50] & in2[50];
    assign P[36] = in1[50] ^ in2[50];
    assign G[37] = in1[49] & in2[49];
    assign P[37] = in1[49] ^ in2[49];
    assign G[38] = in1[48] & in2[48];
    assign P[38] = in1[48] ^ in2[48];
    assign G[39] = in1[47] & in2[47];
    assign P[39] = in1[47] ^ in2[47];
    assign G[40] = in1[46] & in2[46];
    assign P[40] = in1[46] ^ in2[46];
    assign G[41] = in1[45] & in2[45];
    assign P[41] = in1[45] ^ in2[45];
    assign G[42] = in1[44] & in2[44];
    assign P[42] = in1[44] ^ in2[44];
    assign G[43] = in1[43] & in2[43];
    assign P[43] = in1[43] ^ in2[43];
    assign G[44] = in1[42] & in2[42];
    assign P[44] = in1[42] ^ in2[42];
    assign G[45] = in1[41] & in2[41];
    assign P[45] = in1[41] ^ in2[41];
    assign G[46] = in1[40] & in2[40];
    assign P[46] = in1[40] ^ in2[40];
    assign G[47] = in1[39] & in2[39];
    assign P[47] = in1[39] ^ in2[39];
    assign G[48] = in1[38] & in2[38];
    assign P[48] = in1[38] ^ in2[38];
    assign G[49] = in1[37] & in2[37];
    assign P[49] = in1[37] ^ in2[37];
    assign G[50] = in1[36] & in2[36];
    assign P[50] = in1[36] ^ in2[36];
    assign G[51] = in1[35] & in2[35];
    assign P[51] = in1[35] ^ in2[35];
    assign G[52] = in1[34] & in2[34];
    assign P[52] = in1[34] ^ in2[34];
    assign G[53] = in1[33] & in2[33];
    assign P[53] = in1[33] ^ in2[33];
    assign G[54] = in1[32] & in2[32];
    assign P[54] = in1[32] ^ in2[32];
    assign G[55] = in1[31] & in2[31];
    assign P[55] = in1[31] ^ in2[31];
    assign G[56] = in1[30] & in2[30];
    assign P[56] = in1[30] ^ in2[30];
    assign G[57] = in1[29] & in2[29];
    assign P[57] = in1[29] ^ in2[29];
    assign G[58] = in1[28] & in2[28];
    assign P[58] = in1[28] ^ in2[28];
    assign G[59] = in1[27] & in2[27];
    assign P[59] = in1[27] ^ in2[27];
    assign G[60] = in1[26] & in2[26];
    assign P[60] = in1[26] ^ in2[26];
    assign G[61] = in1[25] & in2[25];
    assign P[61] = in1[25] ^ in2[25];
    assign G[62] = in1[24] & in2[24];
    assign P[62] = in1[24] ^ in2[24];
    assign G[63] = in1[23] & in2[23];
    assign P[63] = in1[23] ^ in2[23];
    assign G[64] = in1[22] & in2[22];
    assign P[64] = in1[22] ^ in2[22];
    assign G[65] = in1[21] & in2[21];
    assign P[65] = in1[21] ^ in2[21];
    assign G[66] = in1[20] & in2[20];
    assign P[66] = in1[20] ^ in2[20];
    assign G[67] = in1[19] & in2[19];
    assign P[67] = in1[19] ^ in2[19];
    assign G[68] = in1[18] & in2[18];
    assign P[68] = in1[18] ^ in2[18];
    assign G[69] = in1[17] & in2[17];
    assign P[69] = in1[17] ^ in2[17];
    assign G[70] = in1[16] & in2[16];
    assign P[70] = in1[16] ^ in2[16];
    assign G[71] = in1[15] & in2[15];
    assign P[71] = in1[15] ^ in2[15];
    assign G[72] = in1[14] & in2[14];
    assign P[72] = in1[14] ^ in2[14];
    assign G[73] = in1[13] & in2[13];
    assign P[73] = in1[13] ^ in2[13];
    assign G[74] = in1[12] & in2[12];
    assign P[74] = in1[12] ^ in2[12];
    assign G[75] = in1[11] & in2[11];
    assign P[75] = in1[11] ^ in2[11];
    assign G[76] = in1[10] & in2[10];
    assign P[76] = in1[10] ^ in2[10];
    assign G[77] = in1[9] & in2[9];
    assign P[77] = in1[9] ^ in2[9];
    assign G[78] = in1[8] & in2[8];
    assign P[78] = in1[8] ^ in2[8];
    assign G[79] = in1[7] & in2[7];
    assign P[79] = in1[7] ^ in2[7];
    assign G[80] = in1[6] & in2[6];
    assign P[80] = in1[6] ^ in2[6];
    assign G[81] = in1[5] & in2[5];
    assign P[81] = in1[5] ^ in2[5];
    assign G[82] = in1[4] & in2[4];
    assign P[82] = in1[4] ^ in2[4];
    assign G[83] = in1[3] & in2[3];
    assign P[83] = in1[3] ^ in2[3];
    assign G[84] = in1[2] & in2[2];
    assign P[84] = in1[2] ^ in2[2];
    assign G[85] = in1[1] & in2[1];
    assign P[85] = in1[1] ^ in2[1];
    assign G[86] = in1[0] & in2[0];
    assign P[86] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign cout = G[86] | (P[86] & C[86]);
    assign sum = P ^ C;
endmodule

module CLA_86(output [85:0] sum, output cout, input [85:0] in1, input [85:0] in2);

    wire[85:0] G;
    wire[85:0] C;
    wire[85:0] P;

    assign G[0] = in1[85] & in2[85];
    assign P[0] = in1[85] ^ in2[85];
    assign G[1] = in1[84] & in2[84];
    assign P[1] = in1[84] ^ in2[84];
    assign G[2] = in1[83] & in2[83];
    assign P[2] = in1[83] ^ in2[83];
    assign G[3] = in1[82] & in2[82];
    assign P[3] = in1[82] ^ in2[82];
    assign G[4] = in1[81] & in2[81];
    assign P[4] = in1[81] ^ in2[81];
    assign G[5] = in1[80] & in2[80];
    assign P[5] = in1[80] ^ in2[80];
    assign G[6] = in1[79] & in2[79];
    assign P[6] = in1[79] ^ in2[79];
    assign G[7] = in1[78] & in2[78];
    assign P[7] = in1[78] ^ in2[78];
    assign G[8] = in1[77] & in2[77];
    assign P[8] = in1[77] ^ in2[77];
    assign G[9] = in1[76] & in2[76];
    assign P[9] = in1[76] ^ in2[76];
    assign G[10] = in1[75] & in2[75];
    assign P[10] = in1[75] ^ in2[75];
    assign G[11] = in1[74] & in2[74];
    assign P[11] = in1[74] ^ in2[74];
    assign G[12] = in1[73] & in2[73];
    assign P[12] = in1[73] ^ in2[73];
    assign G[13] = in1[72] & in2[72];
    assign P[13] = in1[72] ^ in2[72];
    assign G[14] = in1[71] & in2[71];
    assign P[14] = in1[71] ^ in2[71];
    assign G[15] = in1[70] & in2[70];
    assign P[15] = in1[70] ^ in2[70];
    assign G[16] = in1[69] & in2[69];
    assign P[16] = in1[69] ^ in2[69];
    assign G[17] = in1[68] & in2[68];
    assign P[17] = in1[68] ^ in2[68];
    assign G[18] = in1[67] & in2[67];
    assign P[18] = in1[67] ^ in2[67];
    assign G[19] = in1[66] & in2[66];
    assign P[19] = in1[66] ^ in2[66];
    assign G[20] = in1[65] & in2[65];
    assign P[20] = in1[65] ^ in2[65];
    assign G[21] = in1[64] & in2[64];
    assign P[21] = in1[64] ^ in2[64];
    assign G[22] = in1[63] & in2[63];
    assign P[22] = in1[63] ^ in2[63];
    assign G[23] = in1[62] & in2[62];
    assign P[23] = in1[62] ^ in2[62];
    assign G[24] = in1[61] & in2[61];
    assign P[24] = in1[61] ^ in2[61];
    assign G[25] = in1[60] & in2[60];
    assign P[25] = in1[60] ^ in2[60];
    assign G[26] = in1[59] & in2[59];
    assign P[26] = in1[59] ^ in2[59];
    assign G[27] = in1[58] & in2[58];
    assign P[27] = in1[58] ^ in2[58];
    assign G[28] = in1[57] & in2[57];
    assign P[28] = in1[57] ^ in2[57];
    assign G[29] = in1[56] & in2[56];
    assign P[29] = in1[56] ^ in2[56];
    assign G[30] = in1[55] & in2[55];
    assign P[30] = in1[55] ^ in2[55];
    assign G[31] = in1[54] & in2[54];
    assign P[31] = in1[54] ^ in2[54];
    assign G[32] = in1[53] & in2[53];
    assign P[32] = in1[53] ^ in2[53];
    assign G[33] = in1[52] & in2[52];
    assign P[33] = in1[52] ^ in2[52];
    assign G[34] = in1[51] & in2[51];
    assign P[34] = in1[51] ^ in2[51];
    assign G[35] = in1[50] & in2[50];
    assign P[35] = in1[50] ^ in2[50];
    assign G[36] = in1[49] & in2[49];
    assign P[36] = in1[49] ^ in2[49];
    assign G[37] = in1[48] & in2[48];
    assign P[37] = in1[48] ^ in2[48];
    assign G[38] = in1[47] & in2[47];
    assign P[38] = in1[47] ^ in2[47];
    assign G[39] = in1[46] & in2[46];
    assign P[39] = in1[46] ^ in2[46];
    assign G[40] = in1[45] & in2[45];
    assign P[40] = in1[45] ^ in2[45];
    assign G[41] = in1[44] & in2[44];
    assign P[41] = in1[44] ^ in2[44];
    assign G[42] = in1[43] & in2[43];
    assign P[42] = in1[43] ^ in2[43];
    assign G[43] = in1[42] & in2[42];
    assign P[43] = in1[42] ^ in2[42];
    assign G[44] = in1[41] & in2[41];
    assign P[44] = in1[41] ^ in2[41];
    assign G[45] = in1[40] & in2[40];
    assign P[45] = in1[40] ^ in2[40];
    assign G[46] = in1[39] & in2[39];
    assign P[46] = in1[39] ^ in2[39];
    assign G[47] = in1[38] & in2[38];
    assign P[47] = in1[38] ^ in2[38];
    assign G[48] = in1[37] & in2[37];
    assign P[48] = in1[37] ^ in2[37];
    assign G[49] = in1[36] & in2[36];
    assign P[49] = in1[36] ^ in2[36];
    assign G[50] = in1[35] & in2[35];
    assign P[50] = in1[35] ^ in2[35];
    assign G[51] = in1[34] & in2[34];
    assign P[51] = in1[34] ^ in2[34];
    assign G[52] = in1[33] & in2[33];
    assign P[52] = in1[33] ^ in2[33];
    assign G[53] = in1[32] & in2[32];
    assign P[53] = in1[32] ^ in2[32];
    assign G[54] = in1[31] & in2[31];
    assign P[54] = in1[31] ^ in2[31];
    assign G[55] = in1[30] & in2[30];
    assign P[55] = in1[30] ^ in2[30];
    assign G[56] = in1[29] & in2[29];
    assign P[56] = in1[29] ^ in2[29];
    assign G[57] = in1[28] & in2[28];
    assign P[57] = in1[28] ^ in2[28];
    assign G[58] = in1[27] & in2[27];
    assign P[58] = in1[27] ^ in2[27];
    assign G[59] = in1[26] & in2[26];
    assign P[59] = in1[26] ^ in2[26];
    assign G[60] = in1[25] & in2[25];
    assign P[60] = in1[25] ^ in2[25];
    assign G[61] = in1[24] & in2[24];
    assign P[61] = in1[24] ^ in2[24];
    assign G[62] = in1[23] & in2[23];
    assign P[62] = in1[23] ^ in2[23];
    assign G[63] = in1[22] & in2[22];
    assign P[63] = in1[22] ^ in2[22];
    assign G[64] = in1[21] & in2[21];
    assign P[64] = in1[21] ^ in2[21];
    assign G[65] = in1[20] & in2[20];
    assign P[65] = in1[20] ^ in2[20];
    assign G[66] = in1[19] & in2[19];
    assign P[66] = in1[19] ^ in2[19];
    assign G[67] = in1[18] & in2[18];
    assign P[67] = in1[18] ^ in2[18];
    assign G[68] = in1[17] & in2[17];
    assign P[68] = in1[17] ^ in2[17];
    assign G[69] = in1[16] & in2[16];
    assign P[69] = in1[16] ^ in2[16];
    assign G[70] = in1[15] & in2[15];
    assign P[70] = in1[15] ^ in2[15];
    assign G[71] = in1[14] & in2[14];
    assign P[71] = in1[14] ^ in2[14];
    assign G[72] = in1[13] & in2[13];
    assign P[72] = in1[13] ^ in2[13];
    assign G[73] = in1[12] & in2[12];
    assign P[73] = in1[12] ^ in2[12];
    assign G[74] = in1[11] & in2[11];
    assign P[74] = in1[11] ^ in2[11];
    assign G[75] = in1[10] & in2[10];
    assign P[75] = in1[10] ^ in2[10];
    assign G[76] = in1[9] & in2[9];
    assign P[76] = in1[9] ^ in2[9];
    assign G[77] = in1[8] & in2[8];
    assign P[77] = in1[8] ^ in2[8];
    assign G[78] = in1[7] & in2[7];
    assign P[78] = in1[7] ^ in2[7];
    assign G[79] = in1[6] & in2[6];
    assign P[79] = in1[6] ^ in2[6];
    assign G[80] = in1[5] & in2[5];
    assign P[80] = in1[5] ^ in2[5];
    assign G[81] = in1[4] & in2[4];
    assign P[81] = in1[4] ^ in2[4];
    assign G[82] = in1[3] & in2[3];
    assign P[82] = in1[3] ^ in2[3];
    assign G[83] = in1[2] & in2[2];
    assign P[83] = in1[2] ^ in2[2];
    assign G[84] = in1[1] & in2[1];
    assign P[84] = in1[1] ^ in2[1];
    assign G[85] = in1[0] & in2[0];
    assign P[85] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign cout = G[85] | (P[85] & C[85]);
    assign sum = P ^ C;
endmodule

module CLA_85(output [84:0] sum, output cout, input [84:0] in1, input [84:0] in2);

    wire[84:0] G;
    wire[84:0] C;
    wire[84:0] P;

    assign G[0] = in1[84] & in2[84];
    assign P[0] = in1[84] ^ in2[84];
    assign G[1] = in1[83] & in2[83];
    assign P[1] = in1[83] ^ in2[83];
    assign G[2] = in1[82] & in2[82];
    assign P[2] = in1[82] ^ in2[82];
    assign G[3] = in1[81] & in2[81];
    assign P[3] = in1[81] ^ in2[81];
    assign G[4] = in1[80] & in2[80];
    assign P[4] = in1[80] ^ in2[80];
    assign G[5] = in1[79] & in2[79];
    assign P[5] = in1[79] ^ in2[79];
    assign G[6] = in1[78] & in2[78];
    assign P[6] = in1[78] ^ in2[78];
    assign G[7] = in1[77] & in2[77];
    assign P[7] = in1[77] ^ in2[77];
    assign G[8] = in1[76] & in2[76];
    assign P[8] = in1[76] ^ in2[76];
    assign G[9] = in1[75] & in2[75];
    assign P[9] = in1[75] ^ in2[75];
    assign G[10] = in1[74] & in2[74];
    assign P[10] = in1[74] ^ in2[74];
    assign G[11] = in1[73] & in2[73];
    assign P[11] = in1[73] ^ in2[73];
    assign G[12] = in1[72] & in2[72];
    assign P[12] = in1[72] ^ in2[72];
    assign G[13] = in1[71] & in2[71];
    assign P[13] = in1[71] ^ in2[71];
    assign G[14] = in1[70] & in2[70];
    assign P[14] = in1[70] ^ in2[70];
    assign G[15] = in1[69] & in2[69];
    assign P[15] = in1[69] ^ in2[69];
    assign G[16] = in1[68] & in2[68];
    assign P[16] = in1[68] ^ in2[68];
    assign G[17] = in1[67] & in2[67];
    assign P[17] = in1[67] ^ in2[67];
    assign G[18] = in1[66] & in2[66];
    assign P[18] = in1[66] ^ in2[66];
    assign G[19] = in1[65] & in2[65];
    assign P[19] = in1[65] ^ in2[65];
    assign G[20] = in1[64] & in2[64];
    assign P[20] = in1[64] ^ in2[64];
    assign G[21] = in1[63] & in2[63];
    assign P[21] = in1[63] ^ in2[63];
    assign G[22] = in1[62] & in2[62];
    assign P[22] = in1[62] ^ in2[62];
    assign G[23] = in1[61] & in2[61];
    assign P[23] = in1[61] ^ in2[61];
    assign G[24] = in1[60] & in2[60];
    assign P[24] = in1[60] ^ in2[60];
    assign G[25] = in1[59] & in2[59];
    assign P[25] = in1[59] ^ in2[59];
    assign G[26] = in1[58] & in2[58];
    assign P[26] = in1[58] ^ in2[58];
    assign G[27] = in1[57] & in2[57];
    assign P[27] = in1[57] ^ in2[57];
    assign G[28] = in1[56] & in2[56];
    assign P[28] = in1[56] ^ in2[56];
    assign G[29] = in1[55] & in2[55];
    assign P[29] = in1[55] ^ in2[55];
    assign G[30] = in1[54] & in2[54];
    assign P[30] = in1[54] ^ in2[54];
    assign G[31] = in1[53] & in2[53];
    assign P[31] = in1[53] ^ in2[53];
    assign G[32] = in1[52] & in2[52];
    assign P[32] = in1[52] ^ in2[52];
    assign G[33] = in1[51] & in2[51];
    assign P[33] = in1[51] ^ in2[51];
    assign G[34] = in1[50] & in2[50];
    assign P[34] = in1[50] ^ in2[50];
    assign G[35] = in1[49] & in2[49];
    assign P[35] = in1[49] ^ in2[49];
    assign G[36] = in1[48] & in2[48];
    assign P[36] = in1[48] ^ in2[48];
    assign G[37] = in1[47] & in2[47];
    assign P[37] = in1[47] ^ in2[47];
    assign G[38] = in1[46] & in2[46];
    assign P[38] = in1[46] ^ in2[46];
    assign G[39] = in1[45] & in2[45];
    assign P[39] = in1[45] ^ in2[45];
    assign G[40] = in1[44] & in2[44];
    assign P[40] = in1[44] ^ in2[44];
    assign G[41] = in1[43] & in2[43];
    assign P[41] = in1[43] ^ in2[43];
    assign G[42] = in1[42] & in2[42];
    assign P[42] = in1[42] ^ in2[42];
    assign G[43] = in1[41] & in2[41];
    assign P[43] = in1[41] ^ in2[41];
    assign G[44] = in1[40] & in2[40];
    assign P[44] = in1[40] ^ in2[40];
    assign G[45] = in1[39] & in2[39];
    assign P[45] = in1[39] ^ in2[39];
    assign G[46] = in1[38] & in2[38];
    assign P[46] = in1[38] ^ in2[38];
    assign G[47] = in1[37] & in2[37];
    assign P[47] = in1[37] ^ in2[37];
    assign G[48] = in1[36] & in2[36];
    assign P[48] = in1[36] ^ in2[36];
    assign G[49] = in1[35] & in2[35];
    assign P[49] = in1[35] ^ in2[35];
    assign G[50] = in1[34] & in2[34];
    assign P[50] = in1[34] ^ in2[34];
    assign G[51] = in1[33] & in2[33];
    assign P[51] = in1[33] ^ in2[33];
    assign G[52] = in1[32] & in2[32];
    assign P[52] = in1[32] ^ in2[32];
    assign G[53] = in1[31] & in2[31];
    assign P[53] = in1[31] ^ in2[31];
    assign G[54] = in1[30] & in2[30];
    assign P[54] = in1[30] ^ in2[30];
    assign G[55] = in1[29] & in2[29];
    assign P[55] = in1[29] ^ in2[29];
    assign G[56] = in1[28] & in2[28];
    assign P[56] = in1[28] ^ in2[28];
    assign G[57] = in1[27] & in2[27];
    assign P[57] = in1[27] ^ in2[27];
    assign G[58] = in1[26] & in2[26];
    assign P[58] = in1[26] ^ in2[26];
    assign G[59] = in1[25] & in2[25];
    assign P[59] = in1[25] ^ in2[25];
    assign G[60] = in1[24] & in2[24];
    assign P[60] = in1[24] ^ in2[24];
    assign G[61] = in1[23] & in2[23];
    assign P[61] = in1[23] ^ in2[23];
    assign G[62] = in1[22] & in2[22];
    assign P[62] = in1[22] ^ in2[22];
    assign G[63] = in1[21] & in2[21];
    assign P[63] = in1[21] ^ in2[21];
    assign G[64] = in1[20] & in2[20];
    assign P[64] = in1[20] ^ in2[20];
    assign G[65] = in1[19] & in2[19];
    assign P[65] = in1[19] ^ in2[19];
    assign G[66] = in1[18] & in2[18];
    assign P[66] = in1[18] ^ in2[18];
    assign G[67] = in1[17] & in2[17];
    assign P[67] = in1[17] ^ in2[17];
    assign G[68] = in1[16] & in2[16];
    assign P[68] = in1[16] ^ in2[16];
    assign G[69] = in1[15] & in2[15];
    assign P[69] = in1[15] ^ in2[15];
    assign G[70] = in1[14] & in2[14];
    assign P[70] = in1[14] ^ in2[14];
    assign G[71] = in1[13] & in2[13];
    assign P[71] = in1[13] ^ in2[13];
    assign G[72] = in1[12] & in2[12];
    assign P[72] = in1[12] ^ in2[12];
    assign G[73] = in1[11] & in2[11];
    assign P[73] = in1[11] ^ in2[11];
    assign G[74] = in1[10] & in2[10];
    assign P[74] = in1[10] ^ in2[10];
    assign G[75] = in1[9] & in2[9];
    assign P[75] = in1[9] ^ in2[9];
    assign G[76] = in1[8] & in2[8];
    assign P[76] = in1[8] ^ in2[8];
    assign G[77] = in1[7] & in2[7];
    assign P[77] = in1[7] ^ in2[7];
    assign G[78] = in1[6] & in2[6];
    assign P[78] = in1[6] ^ in2[6];
    assign G[79] = in1[5] & in2[5];
    assign P[79] = in1[5] ^ in2[5];
    assign G[80] = in1[4] & in2[4];
    assign P[80] = in1[4] ^ in2[4];
    assign G[81] = in1[3] & in2[3];
    assign P[81] = in1[3] ^ in2[3];
    assign G[82] = in1[2] & in2[2];
    assign P[82] = in1[2] ^ in2[2];
    assign G[83] = in1[1] & in2[1];
    assign P[83] = in1[1] ^ in2[1];
    assign G[84] = in1[0] & in2[0];
    assign P[84] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign cout = G[84] | (P[84] & C[84]);
    assign sum = P ^ C;
endmodule

module CLA_84(output [83:0] sum, output cout, input [83:0] in1, input [83:0] in2);

    wire[83:0] G;
    wire[83:0] C;
    wire[83:0] P;

    assign G[0] = in1[83] & in2[83];
    assign P[0] = in1[83] ^ in2[83];
    assign G[1] = in1[82] & in2[82];
    assign P[1] = in1[82] ^ in2[82];
    assign G[2] = in1[81] & in2[81];
    assign P[2] = in1[81] ^ in2[81];
    assign G[3] = in1[80] & in2[80];
    assign P[3] = in1[80] ^ in2[80];
    assign G[4] = in1[79] & in2[79];
    assign P[4] = in1[79] ^ in2[79];
    assign G[5] = in1[78] & in2[78];
    assign P[5] = in1[78] ^ in2[78];
    assign G[6] = in1[77] & in2[77];
    assign P[6] = in1[77] ^ in2[77];
    assign G[7] = in1[76] & in2[76];
    assign P[7] = in1[76] ^ in2[76];
    assign G[8] = in1[75] & in2[75];
    assign P[8] = in1[75] ^ in2[75];
    assign G[9] = in1[74] & in2[74];
    assign P[9] = in1[74] ^ in2[74];
    assign G[10] = in1[73] & in2[73];
    assign P[10] = in1[73] ^ in2[73];
    assign G[11] = in1[72] & in2[72];
    assign P[11] = in1[72] ^ in2[72];
    assign G[12] = in1[71] & in2[71];
    assign P[12] = in1[71] ^ in2[71];
    assign G[13] = in1[70] & in2[70];
    assign P[13] = in1[70] ^ in2[70];
    assign G[14] = in1[69] & in2[69];
    assign P[14] = in1[69] ^ in2[69];
    assign G[15] = in1[68] & in2[68];
    assign P[15] = in1[68] ^ in2[68];
    assign G[16] = in1[67] & in2[67];
    assign P[16] = in1[67] ^ in2[67];
    assign G[17] = in1[66] & in2[66];
    assign P[17] = in1[66] ^ in2[66];
    assign G[18] = in1[65] & in2[65];
    assign P[18] = in1[65] ^ in2[65];
    assign G[19] = in1[64] & in2[64];
    assign P[19] = in1[64] ^ in2[64];
    assign G[20] = in1[63] & in2[63];
    assign P[20] = in1[63] ^ in2[63];
    assign G[21] = in1[62] & in2[62];
    assign P[21] = in1[62] ^ in2[62];
    assign G[22] = in1[61] & in2[61];
    assign P[22] = in1[61] ^ in2[61];
    assign G[23] = in1[60] & in2[60];
    assign P[23] = in1[60] ^ in2[60];
    assign G[24] = in1[59] & in2[59];
    assign P[24] = in1[59] ^ in2[59];
    assign G[25] = in1[58] & in2[58];
    assign P[25] = in1[58] ^ in2[58];
    assign G[26] = in1[57] & in2[57];
    assign P[26] = in1[57] ^ in2[57];
    assign G[27] = in1[56] & in2[56];
    assign P[27] = in1[56] ^ in2[56];
    assign G[28] = in1[55] & in2[55];
    assign P[28] = in1[55] ^ in2[55];
    assign G[29] = in1[54] & in2[54];
    assign P[29] = in1[54] ^ in2[54];
    assign G[30] = in1[53] & in2[53];
    assign P[30] = in1[53] ^ in2[53];
    assign G[31] = in1[52] & in2[52];
    assign P[31] = in1[52] ^ in2[52];
    assign G[32] = in1[51] & in2[51];
    assign P[32] = in1[51] ^ in2[51];
    assign G[33] = in1[50] & in2[50];
    assign P[33] = in1[50] ^ in2[50];
    assign G[34] = in1[49] & in2[49];
    assign P[34] = in1[49] ^ in2[49];
    assign G[35] = in1[48] & in2[48];
    assign P[35] = in1[48] ^ in2[48];
    assign G[36] = in1[47] & in2[47];
    assign P[36] = in1[47] ^ in2[47];
    assign G[37] = in1[46] & in2[46];
    assign P[37] = in1[46] ^ in2[46];
    assign G[38] = in1[45] & in2[45];
    assign P[38] = in1[45] ^ in2[45];
    assign G[39] = in1[44] & in2[44];
    assign P[39] = in1[44] ^ in2[44];
    assign G[40] = in1[43] & in2[43];
    assign P[40] = in1[43] ^ in2[43];
    assign G[41] = in1[42] & in2[42];
    assign P[41] = in1[42] ^ in2[42];
    assign G[42] = in1[41] & in2[41];
    assign P[42] = in1[41] ^ in2[41];
    assign G[43] = in1[40] & in2[40];
    assign P[43] = in1[40] ^ in2[40];
    assign G[44] = in1[39] & in2[39];
    assign P[44] = in1[39] ^ in2[39];
    assign G[45] = in1[38] & in2[38];
    assign P[45] = in1[38] ^ in2[38];
    assign G[46] = in1[37] & in2[37];
    assign P[46] = in1[37] ^ in2[37];
    assign G[47] = in1[36] & in2[36];
    assign P[47] = in1[36] ^ in2[36];
    assign G[48] = in1[35] & in2[35];
    assign P[48] = in1[35] ^ in2[35];
    assign G[49] = in1[34] & in2[34];
    assign P[49] = in1[34] ^ in2[34];
    assign G[50] = in1[33] & in2[33];
    assign P[50] = in1[33] ^ in2[33];
    assign G[51] = in1[32] & in2[32];
    assign P[51] = in1[32] ^ in2[32];
    assign G[52] = in1[31] & in2[31];
    assign P[52] = in1[31] ^ in2[31];
    assign G[53] = in1[30] & in2[30];
    assign P[53] = in1[30] ^ in2[30];
    assign G[54] = in1[29] & in2[29];
    assign P[54] = in1[29] ^ in2[29];
    assign G[55] = in1[28] & in2[28];
    assign P[55] = in1[28] ^ in2[28];
    assign G[56] = in1[27] & in2[27];
    assign P[56] = in1[27] ^ in2[27];
    assign G[57] = in1[26] & in2[26];
    assign P[57] = in1[26] ^ in2[26];
    assign G[58] = in1[25] & in2[25];
    assign P[58] = in1[25] ^ in2[25];
    assign G[59] = in1[24] & in2[24];
    assign P[59] = in1[24] ^ in2[24];
    assign G[60] = in1[23] & in2[23];
    assign P[60] = in1[23] ^ in2[23];
    assign G[61] = in1[22] & in2[22];
    assign P[61] = in1[22] ^ in2[22];
    assign G[62] = in1[21] & in2[21];
    assign P[62] = in1[21] ^ in2[21];
    assign G[63] = in1[20] & in2[20];
    assign P[63] = in1[20] ^ in2[20];
    assign G[64] = in1[19] & in2[19];
    assign P[64] = in1[19] ^ in2[19];
    assign G[65] = in1[18] & in2[18];
    assign P[65] = in1[18] ^ in2[18];
    assign G[66] = in1[17] & in2[17];
    assign P[66] = in1[17] ^ in2[17];
    assign G[67] = in1[16] & in2[16];
    assign P[67] = in1[16] ^ in2[16];
    assign G[68] = in1[15] & in2[15];
    assign P[68] = in1[15] ^ in2[15];
    assign G[69] = in1[14] & in2[14];
    assign P[69] = in1[14] ^ in2[14];
    assign G[70] = in1[13] & in2[13];
    assign P[70] = in1[13] ^ in2[13];
    assign G[71] = in1[12] & in2[12];
    assign P[71] = in1[12] ^ in2[12];
    assign G[72] = in1[11] & in2[11];
    assign P[72] = in1[11] ^ in2[11];
    assign G[73] = in1[10] & in2[10];
    assign P[73] = in1[10] ^ in2[10];
    assign G[74] = in1[9] & in2[9];
    assign P[74] = in1[9] ^ in2[9];
    assign G[75] = in1[8] & in2[8];
    assign P[75] = in1[8] ^ in2[8];
    assign G[76] = in1[7] & in2[7];
    assign P[76] = in1[7] ^ in2[7];
    assign G[77] = in1[6] & in2[6];
    assign P[77] = in1[6] ^ in2[6];
    assign G[78] = in1[5] & in2[5];
    assign P[78] = in1[5] ^ in2[5];
    assign G[79] = in1[4] & in2[4];
    assign P[79] = in1[4] ^ in2[4];
    assign G[80] = in1[3] & in2[3];
    assign P[80] = in1[3] ^ in2[3];
    assign G[81] = in1[2] & in2[2];
    assign P[81] = in1[2] ^ in2[2];
    assign G[82] = in1[1] & in2[1];
    assign P[82] = in1[1] ^ in2[1];
    assign G[83] = in1[0] & in2[0];
    assign P[83] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign cout = G[83] | (P[83] & C[83]);
    assign sum = P ^ C;
endmodule

module CLA_83(output [82:0] sum, output cout, input [82:0] in1, input [82:0] in2);

    wire[82:0] G;
    wire[82:0] C;
    wire[82:0] P;

    assign G[0] = in1[82] & in2[82];
    assign P[0] = in1[82] ^ in2[82];
    assign G[1] = in1[81] & in2[81];
    assign P[1] = in1[81] ^ in2[81];
    assign G[2] = in1[80] & in2[80];
    assign P[2] = in1[80] ^ in2[80];
    assign G[3] = in1[79] & in2[79];
    assign P[3] = in1[79] ^ in2[79];
    assign G[4] = in1[78] & in2[78];
    assign P[4] = in1[78] ^ in2[78];
    assign G[5] = in1[77] & in2[77];
    assign P[5] = in1[77] ^ in2[77];
    assign G[6] = in1[76] & in2[76];
    assign P[6] = in1[76] ^ in2[76];
    assign G[7] = in1[75] & in2[75];
    assign P[7] = in1[75] ^ in2[75];
    assign G[8] = in1[74] & in2[74];
    assign P[8] = in1[74] ^ in2[74];
    assign G[9] = in1[73] & in2[73];
    assign P[9] = in1[73] ^ in2[73];
    assign G[10] = in1[72] & in2[72];
    assign P[10] = in1[72] ^ in2[72];
    assign G[11] = in1[71] & in2[71];
    assign P[11] = in1[71] ^ in2[71];
    assign G[12] = in1[70] & in2[70];
    assign P[12] = in1[70] ^ in2[70];
    assign G[13] = in1[69] & in2[69];
    assign P[13] = in1[69] ^ in2[69];
    assign G[14] = in1[68] & in2[68];
    assign P[14] = in1[68] ^ in2[68];
    assign G[15] = in1[67] & in2[67];
    assign P[15] = in1[67] ^ in2[67];
    assign G[16] = in1[66] & in2[66];
    assign P[16] = in1[66] ^ in2[66];
    assign G[17] = in1[65] & in2[65];
    assign P[17] = in1[65] ^ in2[65];
    assign G[18] = in1[64] & in2[64];
    assign P[18] = in1[64] ^ in2[64];
    assign G[19] = in1[63] & in2[63];
    assign P[19] = in1[63] ^ in2[63];
    assign G[20] = in1[62] & in2[62];
    assign P[20] = in1[62] ^ in2[62];
    assign G[21] = in1[61] & in2[61];
    assign P[21] = in1[61] ^ in2[61];
    assign G[22] = in1[60] & in2[60];
    assign P[22] = in1[60] ^ in2[60];
    assign G[23] = in1[59] & in2[59];
    assign P[23] = in1[59] ^ in2[59];
    assign G[24] = in1[58] & in2[58];
    assign P[24] = in1[58] ^ in2[58];
    assign G[25] = in1[57] & in2[57];
    assign P[25] = in1[57] ^ in2[57];
    assign G[26] = in1[56] & in2[56];
    assign P[26] = in1[56] ^ in2[56];
    assign G[27] = in1[55] & in2[55];
    assign P[27] = in1[55] ^ in2[55];
    assign G[28] = in1[54] & in2[54];
    assign P[28] = in1[54] ^ in2[54];
    assign G[29] = in1[53] & in2[53];
    assign P[29] = in1[53] ^ in2[53];
    assign G[30] = in1[52] & in2[52];
    assign P[30] = in1[52] ^ in2[52];
    assign G[31] = in1[51] & in2[51];
    assign P[31] = in1[51] ^ in2[51];
    assign G[32] = in1[50] & in2[50];
    assign P[32] = in1[50] ^ in2[50];
    assign G[33] = in1[49] & in2[49];
    assign P[33] = in1[49] ^ in2[49];
    assign G[34] = in1[48] & in2[48];
    assign P[34] = in1[48] ^ in2[48];
    assign G[35] = in1[47] & in2[47];
    assign P[35] = in1[47] ^ in2[47];
    assign G[36] = in1[46] & in2[46];
    assign P[36] = in1[46] ^ in2[46];
    assign G[37] = in1[45] & in2[45];
    assign P[37] = in1[45] ^ in2[45];
    assign G[38] = in1[44] & in2[44];
    assign P[38] = in1[44] ^ in2[44];
    assign G[39] = in1[43] & in2[43];
    assign P[39] = in1[43] ^ in2[43];
    assign G[40] = in1[42] & in2[42];
    assign P[40] = in1[42] ^ in2[42];
    assign G[41] = in1[41] & in2[41];
    assign P[41] = in1[41] ^ in2[41];
    assign G[42] = in1[40] & in2[40];
    assign P[42] = in1[40] ^ in2[40];
    assign G[43] = in1[39] & in2[39];
    assign P[43] = in1[39] ^ in2[39];
    assign G[44] = in1[38] & in2[38];
    assign P[44] = in1[38] ^ in2[38];
    assign G[45] = in1[37] & in2[37];
    assign P[45] = in1[37] ^ in2[37];
    assign G[46] = in1[36] & in2[36];
    assign P[46] = in1[36] ^ in2[36];
    assign G[47] = in1[35] & in2[35];
    assign P[47] = in1[35] ^ in2[35];
    assign G[48] = in1[34] & in2[34];
    assign P[48] = in1[34] ^ in2[34];
    assign G[49] = in1[33] & in2[33];
    assign P[49] = in1[33] ^ in2[33];
    assign G[50] = in1[32] & in2[32];
    assign P[50] = in1[32] ^ in2[32];
    assign G[51] = in1[31] & in2[31];
    assign P[51] = in1[31] ^ in2[31];
    assign G[52] = in1[30] & in2[30];
    assign P[52] = in1[30] ^ in2[30];
    assign G[53] = in1[29] & in2[29];
    assign P[53] = in1[29] ^ in2[29];
    assign G[54] = in1[28] & in2[28];
    assign P[54] = in1[28] ^ in2[28];
    assign G[55] = in1[27] & in2[27];
    assign P[55] = in1[27] ^ in2[27];
    assign G[56] = in1[26] & in2[26];
    assign P[56] = in1[26] ^ in2[26];
    assign G[57] = in1[25] & in2[25];
    assign P[57] = in1[25] ^ in2[25];
    assign G[58] = in1[24] & in2[24];
    assign P[58] = in1[24] ^ in2[24];
    assign G[59] = in1[23] & in2[23];
    assign P[59] = in1[23] ^ in2[23];
    assign G[60] = in1[22] & in2[22];
    assign P[60] = in1[22] ^ in2[22];
    assign G[61] = in1[21] & in2[21];
    assign P[61] = in1[21] ^ in2[21];
    assign G[62] = in1[20] & in2[20];
    assign P[62] = in1[20] ^ in2[20];
    assign G[63] = in1[19] & in2[19];
    assign P[63] = in1[19] ^ in2[19];
    assign G[64] = in1[18] & in2[18];
    assign P[64] = in1[18] ^ in2[18];
    assign G[65] = in1[17] & in2[17];
    assign P[65] = in1[17] ^ in2[17];
    assign G[66] = in1[16] & in2[16];
    assign P[66] = in1[16] ^ in2[16];
    assign G[67] = in1[15] & in2[15];
    assign P[67] = in1[15] ^ in2[15];
    assign G[68] = in1[14] & in2[14];
    assign P[68] = in1[14] ^ in2[14];
    assign G[69] = in1[13] & in2[13];
    assign P[69] = in1[13] ^ in2[13];
    assign G[70] = in1[12] & in2[12];
    assign P[70] = in1[12] ^ in2[12];
    assign G[71] = in1[11] & in2[11];
    assign P[71] = in1[11] ^ in2[11];
    assign G[72] = in1[10] & in2[10];
    assign P[72] = in1[10] ^ in2[10];
    assign G[73] = in1[9] & in2[9];
    assign P[73] = in1[9] ^ in2[9];
    assign G[74] = in1[8] & in2[8];
    assign P[74] = in1[8] ^ in2[8];
    assign G[75] = in1[7] & in2[7];
    assign P[75] = in1[7] ^ in2[7];
    assign G[76] = in1[6] & in2[6];
    assign P[76] = in1[6] ^ in2[6];
    assign G[77] = in1[5] & in2[5];
    assign P[77] = in1[5] ^ in2[5];
    assign G[78] = in1[4] & in2[4];
    assign P[78] = in1[4] ^ in2[4];
    assign G[79] = in1[3] & in2[3];
    assign P[79] = in1[3] ^ in2[3];
    assign G[80] = in1[2] & in2[2];
    assign P[80] = in1[2] ^ in2[2];
    assign G[81] = in1[1] & in2[1];
    assign P[81] = in1[1] ^ in2[1];
    assign G[82] = in1[0] & in2[0];
    assign P[82] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign cout = G[82] | (P[82] & C[82]);
    assign sum = P ^ C;
endmodule

module CLA_82(output [81:0] sum, output cout, input [81:0] in1, input [81:0] in2);

    wire[81:0] G;
    wire[81:0] C;
    wire[81:0] P;

    assign G[0] = in1[81] & in2[81];
    assign P[0] = in1[81] ^ in2[81];
    assign G[1] = in1[80] & in2[80];
    assign P[1] = in1[80] ^ in2[80];
    assign G[2] = in1[79] & in2[79];
    assign P[2] = in1[79] ^ in2[79];
    assign G[3] = in1[78] & in2[78];
    assign P[3] = in1[78] ^ in2[78];
    assign G[4] = in1[77] & in2[77];
    assign P[4] = in1[77] ^ in2[77];
    assign G[5] = in1[76] & in2[76];
    assign P[5] = in1[76] ^ in2[76];
    assign G[6] = in1[75] & in2[75];
    assign P[6] = in1[75] ^ in2[75];
    assign G[7] = in1[74] & in2[74];
    assign P[7] = in1[74] ^ in2[74];
    assign G[8] = in1[73] & in2[73];
    assign P[8] = in1[73] ^ in2[73];
    assign G[9] = in1[72] & in2[72];
    assign P[9] = in1[72] ^ in2[72];
    assign G[10] = in1[71] & in2[71];
    assign P[10] = in1[71] ^ in2[71];
    assign G[11] = in1[70] & in2[70];
    assign P[11] = in1[70] ^ in2[70];
    assign G[12] = in1[69] & in2[69];
    assign P[12] = in1[69] ^ in2[69];
    assign G[13] = in1[68] & in2[68];
    assign P[13] = in1[68] ^ in2[68];
    assign G[14] = in1[67] & in2[67];
    assign P[14] = in1[67] ^ in2[67];
    assign G[15] = in1[66] & in2[66];
    assign P[15] = in1[66] ^ in2[66];
    assign G[16] = in1[65] & in2[65];
    assign P[16] = in1[65] ^ in2[65];
    assign G[17] = in1[64] & in2[64];
    assign P[17] = in1[64] ^ in2[64];
    assign G[18] = in1[63] & in2[63];
    assign P[18] = in1[63] ^ in2[63];
    assign G[19] = in1[62] & in2[62];
    assign P[19] = in1[62] ^ in2[62];
    assign G[20] = in1[61] & in2[61];
    assign P[20] = in1[61] ^ in2[61];
    assign G[21] = in1[60] & in2[60];
    assign P[21] = in1[60] ^ in2[60];
    assign G[22] = in1[59] & in2[59];
    assign P[22] = in1[59] ^ in2[59];
    assign G[23] = in1[58] & in2[58];
    assign P[23] = in1[58] ^ in2[58];
    assign G[24] = in1[57] & in2[57];
    assign P[24] = in1[57] ^ in2[57];
    assign G[25] = in1[56] & in2[56];
    assign P[25] = in1[56] ^ in2[56];
    assign G[26] = in1[55] & in2[55];
    assign P[26] = in1[55] ^ in2[55];
    assign G[27] = in1[54] & in2[54];
    assign P[27] = in1[54] ^ in2[54];
    assign G[28] = in1[53] & in2[53];
    assign P[28] = in1[53] ^ in2[53];
    assign G[29] = in1[52] & in2[52];
    assign P[29] = in1[52] ^ in2[52];
    assign G[30] = in1[51] & in2[51];
    assign P[30] = in1[51] ^ in2[51];
    assign G[31] = in1[50] & in2[50];
    assign P[31] = in1[50] ^ in2[50];
    assign G[32] = in1[49] & in2[49];
    assign P[32] = in1[49] ^ in2[49];
    assign G[33] = in1[48] & in2[48];
    assign P[33] = in1[48] ^ in2[48];
    assign G[34] = in1[47] & in2[47];
    assign P[34] = in1[47] ^ in2[47];
    assign G[35] = in1[46] & in2[46];
    assign P[35] = in1[46] ^ in2[46];
    assign G[36] = in1[45] & in2[45];
    assign P[36] = in1[45] ^ in2[45];
    assign G[37] = in1[44] & in2[44];
    assign P[37] = in1[44] ^ in2[44];
    assign G[38] = in1[43] & in2[43];
    assign P[38] = in1[43] ^ in2[43];
    assign G[39] = in1[42] & in2[42];
    assign P[39] = in1[42] ^ in2[42];
    assign G[40] = in1[41] & in2[41];
    assign P[40] = in1[41] ^ in2[41];
    assign G[41] = in1[40] & in2[40];
    assign P[41] = in1[40] ^ in2[40];
    assign G[42] = in1[39] & in2[39];
    assign P[42] = in1[39] ^ in2[39];
    assign G[43] = in1[38] & in2[38];
    assign P[43] = in1[38] ^ in2[38];
    assign G[44] = in1[37] & in2[37];
    assign P[44] = in1[37] ^ in2[37];
    assign G[45] = in1[36] & in2[36];
    assign P[45] = in1[36] ^ in2[36];
    assign G[46] = in1[35] & in2[35];
    assign P[46] = in1[35] ^ in2[35];
    assign G[47] = in1[34] & in2[34];
    assign P[47] = in1[34] ^ in2[34];
    assign G[48] = in1[33] & in2[33];
    assign P[48] = in1[33] ^ in2[33];
    assign G[49] = in1[32] & in2[32];
    assign P[49] = in1[32] ^ in2[32];
    assign G[50] = in1[31] & in2[31];
    assign P[50] = in1[31] ^ in2[31];
    assign G[51] = in1[30] & in2[30];
    assign P[51] = in1[30] ^ in2[30];
    assign G[52] = in1[29] & in2[29];
    assign P[52] = in1[29] ^ in2[29];
    assign G[53] = in1[28] & in2[28];
    assign P[53] = in1[28] ^ in2[28];
    assign G[54] = in1[27] & in2[27];
    assign P[54] = in1[27] ^ in2[27];
    assign G[55] = in1[26] & in2[26];
    assign P[55] = in1[26] ^ in2[26];
    assign G[56] = in1[25] & in2[25];
    assign P[56] = in1[25] ^ in2[25];
    assign G[57] = in1[24] & in2[24];
    assign P[57] = in1[24] ^ in2[24];
    assign G[58] = in1[23] & in2[23];
    assign P[58] = in1[23] ^ in2[23];
    assign G[59] = in1[22] & in2[22];
    assign P[59] = in1[22] ^ in2[22];
    assign G[60] = in1[21] & in2[21];
    assign P[60] = in1[21] ^ in2[21];
    assign G[61] = in1[20] & in2[20];
    assign P[61] = in1[20] ^ in2[20];
    assign G[62] = in1[19] & in2[19];
    assign P[62] = in1[19] ^ in2[19];
    assign G[63] = in1[18] & in2[18];
    assign P[63] = in1[18] ^ in2[18];
    assign G[64] = in1[17] & in2[17];
    assign P[64] = in1[17] ^ in2[17];
    assign G[65] = in1[16] & in2[16];
    assign P[65] = in1[16] ^ in2[16];
    assign G[66] = in1[15] & in2[15];
    assign P[66] = in1[15] ^ in2[15];
    assign G[67] = in1[14] & in2[14];
    assign P[67] = in1[14] ^ in2[14];
    assign G[68] = in1[13] & in2[13];
    assign P[68] = in1[13] ^ in2[13];
    assign G[69] = in1[12] & in2[12];
    assign P[69] = in1[12] ^ in2[12];
    assign G[70] = in1[11] & in2[11];
    assign P[70] = in1[11] ^ in2[11];
    assign G[71] = in1[10] & in2[10];
    assign P[71] = in1[10] ^ in2[10];
    assign G[72] = in1[9] & in2[9];
    assign P[72] = in1[9] ^ in2[9];
    assign G[73] = in1[8] & in2[8];
    assign P[73] = in1[8] ^ in2[8];
    assign G[74] = in1[7] & in2[7];
    assign P[74] = in1[7] ^ in2[7];
    assign G[75] = in1[6] & in2[6];
    assign P[75] = in1[6] ^ in2[6];
    assign G[76] = in1[5] & in2[5];
    assign P[76] = in1[5] ^ in2[5];
    assign G[77] = in1[4] & in2[4];
    assign P[77] = in1[4] ^ in2[4];
    assign G[78] = in1[3] & in2[3];
    assign P[78] = in1[3] ^ in2[3];
    assign G[79] = in1[2] & in2[2];
    assign P[79] = in1[2] ^ in2[2];
    assign G[80] = in1[1] & in2[1];
    assign P[80] = in1[1] ^ in2[1];
    assign G[81] = in1[0] & in2[0];
    assign P[81] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign cout = G[81] | (P[81] & C[81]);
    assign sum = P ^ C;
endmodule

module CLA_81(output [80:0] sum, output cout, input [80:0] in1, input [80:0] in2);

    wire[80:0] G;
    wire[80:0] C;
    wire[80:0] P;

    assign G[0] = in1[80] & in2[80];
    assign P[0] = in1[80] ^ in2[80];
    assign G[1] = in1[79] & in2[79];
    assign P[1] = in1[79] ^ in2[79];
    assign G[2] = in1[78] & in2[78];
    assign P[2] = in1[78] ^ in2[78];
    assign G[3] = in1[77] & in2[77];
    assign P[3] = in1[77] ^ in2[77];
    assign G[4] = in1[76] & in2[76];
    assign P[4] = in1[76] ^ in2[76];
    assign G[5] = in1[75] & in2[75];
    assign P[5] = in1[75] ^ in2[75];
    assign G[6] = in1[74] & in2[74];
    assign P[6] = in1[74] ^ in2[74];
    assign G[7] = in1[73] & in2[73];
    assign P[7] = in1[73] ^ in2[73];
    assign G[8] = in1[72] & in2[72];
    assign P[8] = in1[72] ^ in2[72];
    assign G[9] = in1[71] & in2[71];
    assign P[9] = in1[71] ^ in2[71];
    assign G[10] = in1[70] & in2[70];
    assign P[10] = in1[70] ^ in2[70];
    assign G[11] = in1[69] & in2[69];
    assign P[11] = in1[69] ^ in2[69];
    assign G[12] = in1[68] & in2[68];
    assign P[12] = in1[68] ^ in2[68];
    assign G[13] = in1[67] & in2[67];
    assign P[13] = in1[67] ^ in2[67];
    assign G[14] = in1[66] & in2[66];
    assign P[14] = in1[66] ^ in2[66];
    assign G[15] = in1[65] & in2[65];
    assign P[15] = in1[65] ^ in2[65];
    assign G[16] = in1[64] & in2[64];
    assign P[16] = in1[64] ^ in2[64];
    assign G[17] = in1[63] & in2[63];
    assign P[17] = in1[63] ^ in2[63];
    assign G[18] = in1[62] & in2[62];
    assign P[18] = in1[62] ^ in2[62];
    assign G[19] = in1[61] & in2[61];
    assign P[19] = in1[61] ^ in2[61];
    assign G[20] = in1[60] & in2[60];
    assign P[20] = in1[60] ^ in2[60];
    assign G[21] = in1[59] & in2[59];
    assign P[21] = in1[59] ^ in2[59];
    assign G[22] = in1[58] & in2[58];
    assign P[22] = in1[58] ^ in2[58];
    assign G[23] = in1[57] & in2[57];
    assign P[23] = in1[57] ^ in2[57];
    assign G[24] = in1[56] & in2[56];
    assign P[24] = in1[56] ^ in2[56];
    assign G[25] = in1[55] & in2[55];
    assign P[25] = in1[55] ^ in2[55];
    assign G[26] = in1[54] & in2[54];
    assign P[26] = in1[54] ^ in2[54];
    assign G[27] = in1[53] & in2[53];
    assign P[27] = in1[53] ^ in2[53];
    assign G[28] = in1[52] & in2[52];
    assign P[28] = in1[52] ^ in2[52];
    assign G[29] = in1[51] & in2[51];
    assign P[29] = in1[51] ^ in2[51];
    assign G[30] = in1[50] & in2[50];
    assign P[30] = in1[50] ^ in2[50];
    assign G[31] = in1[49] & in2[49];
    assign P[31] = in1[49] ^ in2[49];
    assign G[32] = in1[48] & in2[48];
    assign P[32] = in1[48] ^ in2[48];
    assign G[33] = in1[47] & in2[47];
    assign P[33] = in1[47] ^ in2[47];
    assign G[34] = in1[46] & in2[46];
    assign P[34] = in1[46] ^ in2[46];
    assign G[35] = in1[45] & in2[45];
    assign P[35] = in1[45] ^ in2[45];
    assign G[36] = in1[44] & in2[44];
    assign P[36] = in1[44] ^ in2[44];
    assign G[37] = in1[43] & in2[43];
    assign P[37] = in1[43] ^ in2[43];
    assign G[38] = in1[42] & in2[42];
    assign P[38] = in1[42] ^ in2[42];
    assign G[39] = in1[41] & in2[41];
    assign P[39] = in1[41] ^ in2[41];
    assign G[40] = in1[40] & in2[40];
    assign P[40] = in1[40] ^ in2[40];
    assign G[41] = in1[39] & in2[39];
    assign P[41] = in1[39] ^ in2[39];
    assign G[42] = in1[38] & in2[38];
    assign P[42] = in1[38] ^ in2[38];
    assign G[43] = in1[37] & in2[37];
    assign P[43] = in1[37] ^ in2[37];
    assign G[44] = in1[36] & in2[36];
    assign P[44] = in1[36] ^ in2[36];
    assign G[45] = in1[35] & in2[35];
    assign P[45] = in1[35] ^ in2[35];
    assign G[46] = in1[34] & in2[34];
    assign P[46] = in1[34] ^ in2[34];
    assign G[47] = in1[33] & in2[33];
    assign P[47] = in1[33] ^ in2[33];
    assign G[48] = in1[32] & in2[32];
    assign P[48] = in1[32] ^ in2[32];
    assign G[49] = in1[31] & in2[31];
    assign P[49] = in1[31] ^ in2[31];
    assign G[50] = in1[30] & in2[30];
    assign P[50] = in1[30] ^ in2[30];
    assign G[51] = in1[29] & in2[29];
    assign P[51] = in1[29] ^ in2[29];
    assign G[52] = in1[28] & in2[28];
    assign P[52] = in1[28] ^ in2[28];
    assign G[53] = in1[27] & in2[27];
    assign P[53] = in1[27] ^ in2[27];
    assign G[54] = in1[26] & in2[26];
    assign P[54] = in1[26] ^ in2[26];
    assign G[55] = in1[25] & in2[25];
    assign P[55] = in1[25] ^ in2[25];
    assign G[56] = in1[24] & in2[24];
    assign P[56] = in1[24] ^ in2[24];
    assign G[57] = in1[23] & in2[23];
    assign P[57] = in1[23] ^ in2[23];
    assign G[58] = in1[22] & in2[22];
    assign P[58] = in1[22] ^ in2[22];
    assign G[59] = in1[21] & in2[21];
    assign P[59] = in1[21] ^ in2[21];
    assign G[60] = in1[20] & in2[20];
    assign P[60] = in1[20] ^ in2[20];
    assign G[61] = in1[19] & in2[19];
    assign P[61] = in1[19] ^ in2[19];
    assign G[62] = in1[18] & in2[18];
    assign P[62] = in1[18] ^ in2[18];
    assign G[63] = in1[17] & in2[17];
    assign P[63] = in1[17] ^ in2[17];
    assign G[64] = in1[16] & in2[16];
    assign P[64] = in1[16] ^ in2[16];
    assign G[65] = in1[15] & in2[15];
    assign P[65] = in1[15] ^ in2[15];
    assign G[66] = in1[14] & in2[14];
    assign P[66] = in1[14] ^ in2[14];
    assign G[67] = in1[13] & in2[13];
    assign P[67] = in1[13] ^ in2[13];
    assign G[68] = in1[12] & in2[12];
    assign P[68] = in1[12] ^ in2[12];
    assign G[69] = in1[11] & in2[11];
    assign P[69] = in1[11] ^ in2[11];
    assign G[70] = in1[10] & in2[10];
    assign P[70] = in1[10] ^ in2[10];
    assign G[71] = in1[9] & in2[9];
    assign P[71] = in1[9] ^ in2[9];
    assign G[72] = in1[8] & in2[8];
    assign P[72] = in1[8] ^ in2[8];
    assign G[73] = in1[7] & in2[7];
    assign P[73] = in1[7] ^ in2[7];
    assign G[74] = in1[6] & in2[6];
    assign P[74] = in1[6] ^ in2[6];
    assign G[75] = in1[5] & in2[5];
    assign P[75] = in1[5] ^ in2[5];
    assign G[76] = in1[4] & in2[4];
    assign P[76] = in1[4] ^ in2[4];
    assign G[77] = in1[3] & in2[3];
    assign P[77] = in1[3] ^ in2[3];
    assign G[78] = in1[2] & in2[2];
    assign P[78] = in1[2] ^ in2[2];
    assign G[79] = in1[1] & in2[1];
    assign P[79] = in1[1] ^ in2[1];
    assign G[80] = in1[0] & in2[0];
    assign P[80] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign cout = G[80] | (P[80] & C[80]);
    assign sum = P ^ C;
endmodule

module CLA_80(output [79:0] sum, output cout, input [79:0] in1, input [79:0] in2);

    wire[79:0] G;
    wire[79:0] C;
    wire[79:0] P;

    assign G[0] = in1[79] & in2[79];
    assign P[0] = in1[79] ^ in2[79];
    assign G[1] = in1[78] & in2[78];
    assign P[1] = in1[78] ^ in2[78];
    assign G[2] = in1[77] & in2[77];
    assign P[2] = in1[77] ^ in2[77];
    assign G[3] = in1[76] & in2[76];
    assign P[3] = in1[76] ^ in2[76];
    assign G[4] = in1[75] & in2[75];
    assign P[4] = in1[75] ^ in2[75];
    assign G[5] = in1[74] & in2[74];
    assign P[5] = in1[74] ^ in2[74];
    assign G[6] = in1[73] & in2[73];
    assign P[6] = in1[73] ^ in2[73];
    assign G[7] = in1[72] & in2[72];
    assign P[7] = in1[72] ^ in2[72];
    assign G[8] = in1[71] & in2[71];
    assign P[8] = in1[71] ^ in2[71];
    assign G[9] = in1[70] & in2[70];
    assign P[9] = in1[70] ^ in2[70];
    assign G[10] = in1[69] & in2[69];
    assign P[10] = in1[69] ^ in2[69];
    assign G[11] = in1[68] & in2[68];
    assign P[11] = in1[68] ^ in2[68];
    assign G[12] = in1[67] & in2[67];
    assign P[12] = in1[67] ^ in2[67];
    assign G[13] = in1[66] & in2[66];
    assign P[13] = in1[66] ^ in2[66];
    assign G[14] = in1[65] & in2[65];
    assign P[14] = in1[65] ^ in2[65];
    assign G[15] = in1[64] & in2[64];
    assign P[15] = in1[64] ^ in2[64];
    assign G[16] = in1[63] & in2[63];
    assign P[16] = in1[63] ^ in2[63];
    assign G[17] = in1[62] & in2[62];
    assign P[17] = in1[62] ^ in2[62];
    assign G[18] = in1[61] & in2[61];
    assign P[18] = in1[61] ^ in2[61];
    assign G[19] = in1[60] & in2[60];
    assign P[19] = in1[60] ^ in2[60];
    assign G[20] = in1[59] & in2[59];
    assign P[20] = in1[59] ^ in2[59];
    assign G[21] = in1[58] & in2[58];
    assign P[21] = in1[58] ^ in2[58];
    assign G[22] = in1[57] & in2[57];
    assign P[22] = in1[57] ^ in2[57];
    assign G[23] = in1[56] & in2[56];
    assign P[23] = in1[56] ^ in2[56];
    assign G[24] = in1[55] & in2[55];
    assign P[24] = in1[55] ^ in2[55];
    assign G[25] = in1[54] & in2[54];
    assign P[25] = in1[54] ^ in2[54];
    assign G[26] = in1[53] & in2[53];
    assign P[26] = in1[53] ^ in2[53];
    assign G[27] = in1[52] & in2[52];
    assign P[27] = in1[52] ^ in2[52];
    assign G[28] = in1[51] & in2[51];
    assign P[28] = in1[51] ^ in2[51];
    assign G[29] = in1[50] & in2[50];
    assign P[29] = in1[50] ^ in2[50];
    assign G[30] = in1[49] & in2[49];
    assign P[30] = in1[49] ^ in2[49];
    assign G[31] = in1[48] & in2[48];
    assign P[31] = in1[48] ^ in2[48];
    assign G[32] = in1[47] & in2[47];
    assign P[32] = in1[47] ^ in2[47];
    assign G[33] = in1[46] & in2[46];
    assign P[33] = in1[46] ^ in2[46];
    assign G[34] = in1[45] & in2[45];
    assign P[34] = in1[45] ^ in2[45];
    assign G[35] = in1[44] & in2[44];
    assign P[35] = in1[44] ^ in2[44];
    assign G[36] = in1[43] & in2[43];
    assign P[36] = in1[43] ^ in2[43];
    assign G[37] = in1[42] & in2[42];
    assign P[37] = in1[42] ^ in2[42];
    assign G[38] = in1[41] & in2[41];
    assign P[38] = in1[41] ^ in2[41];
    assign G[39] = in1[40] & in2[40];
    assign P[39] = in1[40] ^ in2[40];
    assign G[40] = in1[39] & in2[39];
    assign P[40] = in1[39] ^ in2[39];
    assign G[41] = in1[38] & in2[38];
    assign P[41] = in1[38] ^ in2[38];
    assign G[42] = in1[37] & in2[37];
    assign P[42] = in1[37] ^ in2[37];
    assign G[43] = in1[36] & in2[36];
    assign P[43] = in1[36] ^ in2[36];
    assign G[44] = in1[35] & in2[35];
    assign P[44] = in1[35] ^ in2[35];
    assign G[45] = in1[34] & in2[34];
    assign P[45] = in1[34] ^ in2[34];
    assign G[46] = in1[33] & in2[33];
    assign P[46] = in1[33] ^ in2[33];
    assign G[47] = in1[32] & in2[32];
    assign P[47] = in1[32] ^ in2[32];
    assign G[48] = in1[31] & in2[31];
    assign P[48] = in1[31] ^ in2[31];
    assign G[49] = in1[30] & in2[30];
    assign P[49] = in1[30] ^ in2[30];
    assign G[50] = in1[29] & in2[29];
    assign P[50] = in1[29] ^ in2[29];
    assign G[51] = in1[28] & in2[28];
    assign P[51] = in1[28] ^ in2[28];
    assign G[52] = in1[27] & in2[27];
    assign P[52] = in1[27] ^ in2[27];
    assign G[53] = in1[26] & in2[26];
    assign P[53] = in1[26] ^ in2[26];
    assign G[54] = in1[25] & in2[25];
    assign P[54] = in1[25] ^ in2[25];
    assign G[55] = in1[24] & in2[24];
    assign P[55] = in1[24] ^ in2[24];
    assign G[56] = in1[23] & in2[23];
    assign P[56] = in1[23] ^ in2[23];
    assign G[57] = in1[22] & in2[22];
    assign P[57] = in1[22] ^ in2[22];
    assign G[58] = in1[21] & in2[21];
    assign P[58] = in1[21] ^ in2[21];
    assign G[59] = in1[20] & in2[20];
    assign P[59] = in1[20] ^ in2[20];
    assign G[60] = in1[19] & in2[19];
    assign P[60] = in1[19] ^ in2[19];
    assign G[61] = in1[18] & in2[18];
    assign P[61] = in1[18] ^ in2[18];
    assign G[62] = in1[17] & in2[17];
    assign P[62] = in1[17] ^ in2[17];
    assign G[63] = in1[16] & in2[16];
    assign P[63] = in1[16] ^ in2[16];
    assign G[64] = in1[15] & in2[15];
    assign P[64] = in1[15] ^ in2[15];
    assign G[65] = in1[14] & in2[14];
    assign P[65] = in1[14] ^ in2[14];
    assign G[66] = in1[13] & in2[13];
    assign P[66] = in1[13] ^ in2[13];
    assign G[67] = in1[12] & in2[12];
    assign P[67] = in1[12] ^ in2[12];
    assign G[68] = in1[11] & in2[11];
    assign P[68] = in1[11] ^ in2[11];
    assign G[69] = in1[10] & in2[10];
    assign P[69] = in1[10] ^ in2[10];
    assign G[70] = in1[9] & in2[9];
    assign P[70] = in1[9] ^ in2[9];
    assign G[71] = in1[8] & in2[8];
    assign P[71] = in1[8] ^ in2[8];
    assign G[72] = in1[7] & in2[7];
    assign P[72] = in1[7] ^ in2[7];
    assign G[73] = in1[6] & in2[6];
    assign P[73] = in1[6] ^ in2[6];
    assign G[74] = in1[5] & in2[5];
    assign P[74] = in1[5] ^ in2[5];
    assign G[75] = in1[4] & in2[4];
    assign P[75] = in1[4] ^ in2[4];
    assign G[76] = in1[3] & in2[3];
    assign P[76] = in1[3] ^ in2[3];
    assign G[77] = in1[2] & in2[2];
    assign P[77] = in1[2] ^ in2[2];
    assign G[78] = in1[1] & in2[1];
    assign P[78] = in1[1] ^ in2[1];
    assign G[79] = in1[0] & in2[0];
    assign P[79] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign cout = G[79] | (P[79] & C[79]);
    assign sum = P ^ C;
endmodule

module CLA_79(output [78:0] sum, output cout, input [78:0] in1, input [78:0] in2);

    wire[78:0] G;
    wire[78:0] C;
    wire[78:0] P;

    assign G[0] = in1[78] & in2[78];
    assign P[0] = in1[78] ^ in2[78];
    assign G[1] = in1[77] & in2[77];
    assign P[1] = in1[77] ^ in2[77];
    assign G[2] = in1[76] & in2[76];
    assign P[2] = in1[76] ^ in2[76];
    assign G[3] = in1[75] & in2[75];
    assign P[3] = in1[75] ^ in2[75];
    assign G[4] = in1[74] & in2[74];
    assign P[4] = in1[74] ^ in2[74];
    assign G[5] = in1[73] & in2[73];
    assign P[5] = in1[73] ^ in2[73];
    assign G[6] = in1[72] & in2[72];
    assign P[6] = in1[72] ^ in2[72];
    assign G[7] = in1[71] & in2[71];
    assign P[7] = in1[71] ^ in2[71];
    assign G[8] = in1[70] & in2[70];
    assign P[8] = in1[70] ^ in2[70];
    assign G[9] = in1[69] & in2[69];
    assign P[9] = in1[69] ^ in2[69];
    assign G[10] = in1[68] & in2[68];
    assign P[10] = in1[68] ^ in2[68];
    assign G[11] = in1[67] & in2[67];
    assign P[11] = in1[67] ^ in2[67];
    assign G[12] = in1[66] & in2[66];
    assign P[12] = in1[66] ^ in2[66];
    assign G[13] = in1[65] & in2[65];
    assign P[13] = in1[65] ^ in2[65];
    assign G[14] = in1[64] & in2[64];
    assign P[14] = in1[64] ^ in2[64];
    assign G[15] = in1[63] & in2[63];
    assign P[15] = in1[63] ^ in2[63];
    assign G[16] = in1[62] & in2[62];
    assign P[16] = in1[62] ^ in2[62];
    assign G[17] = in1[61] & in2[61];
    assign P[17] = in1[61] ^ in2[61];
    assign G[18] = in1[60] & in2[60];
    assign P[18] = in1[60] ^ in2[60];
    assign G[19] = in1[59] & in2[59];
    assign P[19] = in1[59] ^ in2[59];
    assign G[20] = in1[58] & in2[58];
    assign P[20] = in1[58] ^ in2[58];
    assign G[21] = in1[57] & in2[57];
    assign P[21] = in1[57] ^ in2[57];
    assign G[22] = in1[56] & in2[56];
    assign P[22] = in1[56] ^ in2[56];
    assign G[23] = in1[55] & in2[55];
    assign P[23] = in1[55] ^ in2[55];
    assign G[24] = in1[54] & in2[54];
    assign P[24] = in1[54] ^ in2[54];
    assign G[25] = in1[53] & in2[53];
    assign P[25] = in1[53] ^ in2[53];
    assign G[26] = in1[52] & in2[52];
    assign P[26] = in1[52] ^ in2[52];
    assign G[27] = in1[51] & in2[51];
    assign P[27] = in1[51] ^ in2[51];
    assign G[28] = in1[50] & in2[50];
    assign P[28] = in1[50] ^ in2[50];
    assign G[29] = in1[49] & in2[49];
    assign P[29] = in1[49] ^ in2[49];
    assign G[30] = in1[48] & in2[48];
    assign P[30] = in1[48] ^ in2[48];
    assign G[31] = in1[47] & in2[47];
    assign P[31] = in1[47] ^ in2[47];
    assign G[32] = in1[46] & in2[46];
    assign P[32] = in1[46] ^ in2[46];
    assign G[33] = in1[45] & in2[45];
    assign P[33] = in1[45] ^ in2[45];
    assign G[34] = in1[44] & in2[44];
    assign P[34] = in1[44] ^ in2[44];
    assign G[35] = in1[43] & in2[43];
    assign P[35] = in1[43] ^ in2[43];
    assign G[36] = in1[42] & in2[42];
    assign P[36] = in1[42] ^ in2[42];
    assign G[37] = in1[41] & in2[41];
    assign P[37] = in1[41] ^ in2[41];
    assign G[38] = in1[40] & in2[40];
    assign P[38] = in1[40] ^ in2[40];
    assign G[39] = in1[39] & in2[39];
    assign P[39] = in1[39] ^ in2[39];
    assign G[40] = in1[38] & in2[38];
    assign P[40] = in1[38] ^ in2[38];
    assign G[41] = in1[37] & in2[37];
    assign P[41] = in1[37] ^ in2[37];
    assign G[42] = in1[36] & in2[36];
    assign P[42] = in1[36] ^ in2[36];
    assign G[43] = in1[35] & in2[35];
    assign P[43] = in1[35] ^ in2[35];
    assign G[44] = in1[34] & in2[34];
    assign P[44] = in1[34] ^ in2[34];
    assign G[45] = in1[33] & in2[33];
    assign P[45] = in1[33] ^ in2[33];
    assign G[46] = in1[32] & in2[32];
    assign P[46] = in1[32] ^ in2[32];
    assign G[47] = in1[31] & in2[31];
    assign P[47] = in1[31] ^ in2[31];
    assign G[48] = in1[30] & in2[30];
    assign P[48] = in1[30] ^ in2[30];
    assign G[49] = in1[29] & in2[29];
    assign P[49] = in1[29] ^ in2[29];
    assign G[50] = in1[28] & in2[28];
    assign P[50] = in1[28] ^ in2[28];
    assign G[51] = in1[27] & in2[27];
    assign P[51] = in1[27] ^ in2[27];
    assign G[52] = in1[26] & in2[26];
    assign P[52] = in1[26] ^ in2[26];
    assign G[53] = in1[25] & in2[25];
    assign P[53] = in1[25] ^ in2[25];
    assign G[54] = in1[24] & in2[24];
    assign P[54] = in1[24] ^ in2[24];
    assign G[55] = in1[23] & in2[23];
    assign P[55] = in1[23] ^ in2[23];
    assign G[56] = in1[22] & in2[22];
    assign P[56] = in1[22] ^ in2[22];
    assign G[57] = in1[21] & in2[21];
    assign P[57] = in1[21] ^ in2[21];
    assign G[58] = in1[20] & in2[20];
    assign P[58] = in1[20] ^ in2[20];
    assign G[59] = in1[19] & in2[19];
    assign P[59] = in1[19] ^ in2[19];
    assign G[60] = in1[18] & in2[18];
    assign P[60] = in1[18] ^ in2[18];
    assign G[61] = in1[17] & in2[17];
    assign P[61] = in1[17] ^ in2[17];
    assign G[62] = in1[16] & in2[16];
    assign P[62] = in1[16] ^ in2[16];
    assign G[63] = in1[15] & in2[15];
    assign P[63] = in1[15] ^ in2[15];
    assign G[64] = in1[14] & in2[14];
    assign P[64] = in1[14] ^ in2[14];
    assign G[65] = in1[13] & in2[13];
    assign P[65] = in1[13] ^ in2[13];
    assign G[66] = in1[12] & in2[12];
    assign P[66] = in1[12] ^ in2[12];
    assign G[67] = in1[11] & in2[11];
    assign P[67] = in1[11] ^ in2[11];
    assign G[68] = in1[10] & in2[10];
    assign P[68] = in1[10] ^ in2[10];
    assign G[69] = in1[9] & in2[9];
    assign P[69] = in1[9] ^ in2[9];
    assign G[70] = in1[8] & in2[8];
    assign P[70] = in1[8] ^ in2[8];
    assign G[71] = in1[7] & in2[7];
    assign P[71] = in1[7] ^ in2[7];
    assign G[72] = in1[6] & in2[6];
    assign P[72] = in1[6] ^ in2[6];
    assign G[73] = in1[5] & in2[5];
    assign P[73] = in1[5] ^ in2[5];
    assign G[74] = in1[4] & in2[4];
    assign P[74] = in1[4] ^ in2[4];
    assign G[75] = in1[3] & in2[3];
    assign P[75] = in1[3] ^ in2[3];
    assign G[76] = in1[2] & in2[2];
    assign P[76] = in1[2] ^ in2[2];
    assign G[77] = in1[1] & in2[1];
    assign P[77] = in1[1] ^ in2[1];
    assign G[78] = in1[0] & in2[0];
    assign P[78] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign cout = G[78] | (P[78] & C[78]);
    assign sum = P ^ C;
endmodule

module CLA_78(output [77:0] sum, output cout, input [77:0] in1, input [77:0] in2);

    wire[77:0] G;
    wire[77:0] C;
    wire[77:0] P;

    assign G[0] = in1[77] & in2[77];
    assign P[0] = in1[77] ^ in2[77];
    assign G[1] = in1[76] & in2[76];
    assign P[1] = in1[76] ^ in2[76];
    assign G[2] = in1[75] & in2[75];
    assign P[2] = in1[75] ^ in2[75];
    assign G[3] = in1[74] & in2[74];
    assign P[3] = in1[74] ^ in2[74];
    assign G[4] = in1[73] & in2[73];
    assign P[4] = in1[73] ^ in2[73];
    assign G[5] = in1[72] & in2[72];
    assign P[5] = in1[72] ^ in2[72];
    assign G[6] = in1[71] & in2[71];
    assign P[6] = in1[71] ^ in2[71];
    assign G[7] = in1[70] & in2[70];
    assign P[7] = in1[70] ^ in2[70];
    assign G[8] = in1[69] & in2[69];
    assign P[8] = in1[69] ^ in2[69];
    assign G[9] = in1[68] & in2[68];
    assign P[9] = in1[68] ^ in2[68];
    assign G[10] = in1[67] & in2[67];
    assign P[10] = in1[67] ^ in2[67];
    assign G[11] = in1[66] & in2[66];
    assign P[11] = in1[66] ^ in2[66];
    assign G[12] = in1[65] & in2[65];
    assign P[12] = in1[65] ^ in2[65];
    assign G[13] = in1[64] & in2[64];
    assign P[13] = in1[64] ^ in2[64];
    assign G[14] = in1[63] & in2[63];
    assign P[14] = in1[63] ^ in2[63];
    assign G[15] = in1[62] & in2[62];
    assign P[15] = in1[62] ^ in2[62];
    assign G[16] = in1[61] & in2[61];
    assign P[16] = in1[61] ^ in2[61];
    assign G[17] = in1[60] & in2[60];
    assign P[17] = in1[60] ^ in2[60];
    assign G[18] = in1[59] & in2[59];
    assign P[18] = in1[59] ^ in2[59];
    assign G[19] = in1[58] & in2[58];
    assign P[19] = in1[58] ^ in2[58];
    assign G[20] = in1[57] & in2[57];
    assign P[20] = in1[57] ^ in2[57];
    assign G[21] = in1[56] & in2[56];
    assign P[21] = in1[56] ^ in2[56];
    assign G[22] = in1[55] & in2[55];
    assign P[22] = in1[55] ^ in2[55];
    assign G[23] = in1[54] & in2[54];
    assign P[23] = in1[54] ^ in2[54];
    assign G[24] = in1[53] & in2[53];
    assign P[24] = in1[53] ^ in2[53];
    assign G[25] = in1[52] & in2[52];
    assign P[25] = in1[52] ^ in2[52];
    assign G[26] = in1[51] & in2[51];
    assign P[26] = in1[51] ^ in2[51];
    assign G[27] = in1[50] & in2[50];
    assign P[27] = in1[50] ^ in2[50];
    assign G[28] = in1[49] & in2[49];
    assign P[28] = in1[49] ^ in2[49];
    assign G[29] = in1[48] & in2[48];
    assign P[29] = in1[48] ^ in2[48];
    assign G[30] = in1[47] & in2[47];
    assign P[30] = in1[47] ^ in2[47];
    assign G[31] = in1[46] & in2[46];
    assign P[31] = in1[46] ^ in2[46];
    assign G[32] = in1[45] & in2[45];
    assign P[32] = in1[45] ^ in2[45];
    assign G[33] = in1[44] & in2[44];
    assign P[33] = in1[44] ^ in2[44];
    assign G[34] = in1[43] & in2[43];
    assign P[34] = in1[43] ^ in2[43];
    assign G[35] = in1[42] & in2[42];
    assign P[35] = in1[42] ^ in2[42];
    assign G[36] = in1[41] & in2[41];
    assign P[36] = in1[41] ^ in2[41];
    assign G[37] = in1[40] & in2[40];
    assign P[37] = in1[40] ^ in2[40];
    assign G[38] = in1[39] & in2[39];
    assign P[38] = in1[39] ^ in2[39];
    assign G[39] = in1[38] & in2[38];
    assign P[39] = in1[38] ^ in2[38];
    assign G[40] = in1[37] & in2[37];
    assign P[40] = in1[37] ^ in2[37];
    assign G[41] = in1[36] & in2[36];
    assign P[41] = in1[36] ^ in2[36];
    assign G[42] = in1[35] & in2[35];
    assign P[42] = in1[35] ^ in2[35];
    assign G[43] = in1[34] & in2[34];
    assign P[43] = in1[34] ^ in2[34];
    assign G[44] = in1[33] & in2[33];
    assign P[44] = in1[33] ^ in2[33];
    assign G[45] = in1[32] & in2[32];
    assign P[45] = in1[32] ^ in2[32];
    assign G[46] = in1[31] & in2[31];
    assign P[46] = in1[31] ^ in2[31];
    assign G[47] = in1[30] & in2[30];
    assign P[47] = in1[30] ^ in2[30];
    assign G[48] = in1[29] & in2[29];
    assign P[48] = in1[29] ^ in2[29];
    assign G[49] = in1[28] & in2[28];
    assign P[49] = in1[28] ^ in2[28];
    assign G[50] = in1[27] & in2[27];
    assign P[50] = in1[27] ^ in2[27];
    assign G[51] = in1[26] & in2[26];
    assign P[51] = in1[26] ^ in2[26];
    assign G[52] = in1[25] & in2[25];
    assign P[52] = in1[25] ^ in2[25];
    assign G[53] = in1[24] & in2[24];
    assign P[53] = in1[24] ^ in2[24];
    assign G[54] = in1[23] & in2[23];
    assign P[54] = in1[23] ^ in2[23];
    assign G[55] = in1[22] & in2[22];
    assign P[55] = in1[22] ^ in2[22];
    assign G[56] = in1[21] & in2[21];
    assign P[56] = in1[21] ^ in2[21];
    assign G[57] = in1[20] & in2[20];
    assign P[57] = in1[20] ^ in2[20];
    assign G[58] = in1[19] & in2[19];
    assign P[58] = in1[19] ^ in2[19];
    assign G[59] = in1[18] & in2[18];
    assign P[59] = in1[18] ^ in2[18];
    assign G[60] = in1[17] & in2[17];
    assign P[60] = in1[17] ^ in2[17];
    assign G[61] = in1[16] & in2[16];
    assign P[61] = in1[16] ^ in2[16];
    assign G[62] = in1[15] & in2[15];
    assign P[62] = in1[15] ^ in2[15];
    assign G[63] = in1[14] & in2[14];
    assign P[63] = in1[14] ^ in2[14];
    assign G[64] = in1[13] & in2[13];
    assign P[64] = in1[13] ^ in2[13];
    assign G[65] = in1[12] & in2[12];
    assign P[65] = in1[12] ^ in2[12];
    assign G[66] = in1[11] & in2[11];
    assign P[66] = in1[11] ^ in2[11];
    assign G[67] = in1[10] & in2[10];
    assign P[67] = in1[10] ^ in2[10];
    assign G[68] = in1[9] & in2[9];
    assign P[68] = in1[9] ^ in2[9];
    assign G[69] = in1[8] & in2[8];
    assign P[69] = in1[8] ^ in2[8];
    assign G[70] = in1[7] & in2[7];
    assign P[70] = in1[7] ^ in2[7];
    assign G[71] = in1[6] & in2[6];
    assign P[71] = in1[6] ^ in2[6];
    assign G[72] = in1[5] & in2[5];
    assign P[72] = in1[5] ^ in2[5];
    assign G[73] = in1[4] & in2[4];
    assign P[73] = in1[4] ^ in2[4];
    assign G[74] = in1[3] & in2[3];
    assign P[74] = in1[3] ^ in2[3];
    assign G[75] = in1[2] & in2[2];
    assign P[75] = in1[2] ^ in2[2];
    assign G[76] = in1[1] & in2[1];
    assign P[76] = in1[1] ^ in2[1];
    assign G[77] = in1[0] & in2[0];
    assign P[77] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign cout = G[77] | (P[77] & C[77]);
    assign sum = P ^ C;
endmodule

module CLA_77(output [76:0] sum, output cout, input [76:0] in1, input [76:0] in2);

    wire[76:0] G;
    wire[76:0] C;
    wire[76:0] P;

    assign G[0] = in1[76] & in2[76];
    assign P[0] = in1[76] ^ in2[76];
    assign G[1] = in1[75] & in2[75];
    assign P[1] = in1[75] ^ in2[75];
    assign G[2] = in1[74] & in2[74];
    assign P[2] = in1[74] ^ in2[74];
    assign G[3] = in1[73] & in2[73];
    assign P[3] = in1[73] ^ in2[73];
    assign G[4] = in1[72] & in2[72];
    assign P[4] = in1[72] ^ in2[72];
    assign G[5] = in1[71] & in2[71];
    assign P[5] = in1[71] ^ in2[71];
    assign G[6] = in1[70] & in2[70];
    assign P[6] = in1[70] ^ in2[70];
    assign G[7] = in1[69] & in2[69];
    assign P[7] = in1[69] ^ in2[69];
    assign G[8] = in1[68] & in2[68];
    assign P[8] = in1[68] ^ in2[68];
    assign G[9] = in1[67] & in2[67];
    assign P[9] = in1[67] ^ in2[67];
    assign G[10] = in1[66] & in2[66];
    assign P[10] = in1[66] ^ in2[66];
    assign G[11] = in1[65] & in2[65];
    assign P[11] = in1[65] ^ in2[65];
    assign G[12] = in1[64] & in2[64];
    assign P[12] = in1[64] ^ in2[64];
    assign G[13] = in1[63] & in2[63];
    assign P[13] = in1[63] ^ in2[63];
    assign G[14] = in1[62] & in2[62];
    assign P[14] = in1[62] ^ in2[62];
    assign G[15] = in1[61] & in2[61];
    assign P[15] = in1[61] ^ in2[61];
    assign G[16] = in1[60] & in2[60];
    assign P[16] = in1[60] ^ in2[60];
    assign G[17] = in1[59] & in2[59];
    assign P[17] = in1[59] ^ in2[59];
    assign G[18] = in1[58] & in2[58];
    assign P[18] = in1[58] ^ in2[58];
    assign G[19] = in1[57] & in2[57];
    assign P[19] = in1[57] ^ in2[57];
    assign G[20] = in1[56] & in2[56];
    assign P[20] = in1[56] ^ in2[56];
    assign G[21] = in1[55] & in2[55];
    assign P[21] = in1[55] ^ in2[55];
    assign G[22] = in1[54] & in2[54];
    assign P[22] = in1[54] ^ in2[54];
    assign G[23] = in1[53] & in2[53];
    assign P[23] = in1[53] ^ in2[53];
    assign G[24] = in1[52] & in2[52];
    assign P[24] = in1[52] ^ in2[52];
    assign G[25] = in1[51] & in2[51];
    assign P[25] = in1[51] ^ in2[51];
    assign G[26] = in1[50] & in2[50];
    assign P[26] = in1[50] ^ in2[50];
    assign G[27] = in1[49] & in2[49];
    assign P[27] = in1[49] ^ in2[49];
    assign G[28] = in1[48] & in2[48];
    assign P[28] = in1[48] ^ in2[48];
    assign G[29] = in1[47] & in2[47];
    assign P[29] = in1[47] ^ in2[47];
    assign G[30] = in1[46] & in2[46];
    assign P[30] = in1[46] ^ in2[46];
    assign G[31] = in1[45] & in2[45];
    assign P[31] = in1[45] ^ in2[45];
    assign G[32] = in1[44] & in2[44];
    assign P[32] = in1[44] ^ in2[44];
    assign G[33] = in1[43] & in2[43];
    assign P[33] = in1[43] ^ in2[43];
    assign G[34] = in1[42] & in2[42];
    assign P[34] = in1[42] ^ in2[42];
    assign G[35] = in1[41] & in2[41];
    assign P[35] = in1[41] ^ in2[41];
    assign G[36] = in1[40] & in2[40];
    assign P[36] = in1[40] ^ in2[40];
    assign G[37] = in1[39] & in2[39];
    assign P[37] = in1[39] ^ in2[39];
    assign G[38] = in1[38] & in2[38];
    assign P[38] = in1[38] ^ in2[38];
    assign G[39] = in1[37] & in2[37];
    assign P[39] = in1[37] ^ in2[37];
    assign G[40] = in1[36] & in2[36];
    assign P[40] = in1[36] ^ in2[36];
    assign G[41] = in1[35] & in2[35];
    assign P[41] = in1[35] ^ in2[35];
    assign G[42] = in1[34] & in2[34];
    assign P[42] = in1[34] ^ in2[34];
    assign G[43] = in1[33] & in2[33];
    assign P[43] = in1[33] ^ in2[33];
    assign G[44] = in1[32] & in2[32];
    assign P[44] = in1[32] ^ in2[32];
    assign G[45] = in1[31] & in2[31];
    assign P[45] = in1[31] ^ in2[31];
    assign G[46] = in1[30] & in2[30];
    assign P[46] = in1[30] ^ in2[30];
    assign G[47] = in1[29] & in2[29];
    assign P[47] = in1[29] ^ in2[29];
    assign G[48] = in1[28] & in2[28];
    assign P[48] = in1[28] ^ in2[28];
    assign G[49] = in1[27] & in2[27];
    assign P[49] = in1[27] ^ in2[27];
    assign G[50] = in1[26] & in2[26];
    assign P[50] = in1[26] ^ in2[26];
    assign G[51] = in1[25] & in2[25];
    assign P[51] = in1[25] ^ in2[25];
    assign G[52] = in1[24] & in2[24];
    assign P[52] = in1[24] ^ in2[24];
    assign G[53] = in1[23] & in2[23];
    assign P[53] = in1[23] ^ in2[23];
    assign G[54] = in1[22] & in2[22];
    assign P[54] = in1[22] ^ in2[22];
    assign G[55] = in1[21] & in2[21];
    assign P[55] = in1[21] ^ in2[21];
    assign G[56] = in1[20] & in2[20];
    assign P[56] = in1[20] ^ in2[20];
    assign G[57] = in1[19] & in2[19];
    assign P[57] = in1[19] ^ in2[19];
    assign G[58] = in1[18] & in2[18];
    assign P[58] = in1[18] ^ in2[18];
    assign G[59] = in1[17] & in2[17];
    assign P[59] = in1[17] ^ in2[17];
    assign G[60] = in1[16] & in2[16];
    assign P[60] = in1[16] ^ in2[16];
    assign G[61] = in1[15] & in2[15];
    assign P[61] = in1[15] ^ in2[15];
    assign G[62] = in1[14] & in2[14];
    assign P[62] = in1[14] ^ in2[14];
    assign G[63] = in1[13] & in2[13];
    assign P[63] = in1[13] ^ in2[13];
    assign G[64] = in1[12] & in2[12];
    assign P[64] = in1[12] ^ in2[12];
    assign G[65] = in1[11] & in2[11];
    assign P[65] = in1[11] ^ in2[11];
    assign G[66] = in1[10] & in2[10];
    assign P[66] = in1[10] ^ in2[10];
    assign G[67] = in1[9] & in2[9];
    assign P[67] = in1[9] ^ in2[9];
    assign G[68] = in1[8] & in2[8];
    assign P[68] = in1[8] ^ in2[8];
    assign G[69] = in1[7] & in2[7];
    assign P[69] = in1[7] ^ in2[7];
    assign G[70] = in1[6] & in2[6];
    assign P[70] = in1[6] ^ in2[6];
    assign G[71] = in1[5] & in2[5];
    assign P[71] = in1[5] ^ in2[5];
    assign G[72] = in1[4] & in2[4];
    assign P[72] = in1[4] ^ in2[4];
    assign G[73] = in1[3] & in2[3];
    assign P[73] = in1[3] ^ in2[3];
    assign G[74] = in1[2] & in2[2];
    assign P[74] = in1[2] ^ in2[2];
    assign G[75] = in1[1] & in2[1];
    assign P[75] = in1[1] ^ in2[1];
    assign G[76] = in1[0] & in2[0];
    assign P[76] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign cout = G[76] | (P[76] & C[76]);
    assign sum = P ^ C;
endmodule

module CLA_76(output [75:0] sum, output cout, input [75:0] in1, input [75:0] in2);

    wire[75:0] G;
    wire[75:0] C;
    wire[75:0] P;

    assign G[0] = in1[75] & in2[75];
    assign P[0] = in1[75] ^ in2[75];
    assign G[1] = in1[74] & in2[74];
    assign P[1] = in1[74] ^ in2[74];
    assign G[2] = in1[73] & in2[73];
    assign P[2] = in1[73] ^ in2[73];
    assign G[3] = in1[72] & in2[72];
    assign P[3] = in1[72] ^ in2[72];
    assign G[4] = in1[71] & in2[71];
    assign P[4] = in1[71] ^ in2[71];
    assign G[5] = in1[70] & in2[70];
    assign P[5] = in1[70] ^ in2[70];
    assign G[6] = in1[69] & in2[69];
    assign P[6] = in1[69] ^ in2[69];
    assign G[7] = in1[68] & in2[68];
    assign P[7] = in1[68] ^ in2[68];
    assign G[8] = in1[67] & in2[67];
    assign P[8] = in1[67] ^ in2[67];
    assign G[9] = in1[66] & in2[66];
    assign P[9] = in1[66] ^ in2[66];
    assign G[10] = in1[65] & in2[65];
    assign P[10] = in1[65] ^ in2[65];
    assign G[11] = in1[64] & in2[64];
    assign P[11] = in1[64] ^ in2[64];
    assign G[12] = in1[63] & in2[63];
    assign P[12] = in1[63] ^ in2[63];
    assign G[13] = in1[62] & in2[62];
    assign P[13] = in1[62] ^ in2[62];
    assign G[14] = in1[61] & in2[61];
    assign P[14] = in1[61] ^ in2[61];
    assign G[15] = in1[60] & in2[60];
    assign P[15] = in1[60] ^ in2[60];
    assign G[16] = in1[59] & in2[59];
    assign P[16] = in1[59] ^ in2[59];
    assign G[17] = in1[58] & in2[58];
    assign P[17] = in1[58] ^ in2[58];
    assign G[18] = in1[57] & in2[57];
    assign P[18] = in1[57] ^ in2[57];
    assign G[19] = in1[56] & in2[56];
    assign P[19] = in1[56] ^ in2[56];
    assign G[20] = in1[55] & in2[55];
    assign P[20] = in1[55] ^ in2[55];
    assign G[21] = in1[54] & in2[54];
    assign P[21] = in1[54] ^ in2[54];
    assign G[22] = in1[53] & in2[53];
    assign P[22] = in1[53] ^ in2[53];
    assign G[23] = in1[52] & in2[52];
    assign P[23] = in1[52] ^ in2[52];
    assign G[24] = in1[51] & in2[51];
    assign P[24] = in1[51] ^ in2[51];
    assign G[25] = in1[50] & in2[50];
    assign P[25] = in1[50] ^ in2[50];
    assign G[26] = in1[49] & in2[49];
    assign P[26] = in1[49] ^ in2[49];
    assign G[27] = in1[48] & in2[48];
    assign P[27] = in1[48] ^ in2[48];
    assign G[28] = in1[47] & in2[47];
    assign P[28] = in1[47] ^ in2[47];
    assign G[29] = in1[46] & in2[46];
    assign P[29] = in1[46] ^ in2[46];
    assign G[30] = in1[45] & in2[45];
    assign P[30] = in1[45] ^ in2[45];
    assign G[31] = in1[44] & in2[44];
    assign P[31] = in1[44] ^ in2[44];
    assign G[32] = in1[43] & in2[43];
    assign P[32] = in1[43] ^ in2[43];
    assign G[33] = in1[42] & in2[42];
    assign P[33] = in1[42] ^ in2[42];
    assign G[34] = in1[41] & in2[41];
    assign P[34] = in1[41] ^ in2[41];
    assign G[35] = in1[40] & in2[40];
    assign P[35] = in1[40] ^ in2[40];
    assign G[36] = in1[39] & in2[39];
    assign P[36] = in1[39] ^ in2[39];
    assign G[37] = in1[38] & in2[38];
    assign P[37] = in1[38] ^ in2[38];
    assign G[38] = in1[37] & in2[37];
    assign P[38] = in1[37] ^ in2[37];
    assign G[39] = in1[36] & in2[36];
    assign P[39] = in1[36] ^ in2[36];
    assign G[40] = in1[35] & in2[35];
    assign P[40] = in1[35] ^ in2[35];
    assign G[41] = in1[34] & in2[34];
    assign P[41] = in1[34] ^ in2[34];
    assign G[42] = in1[33] & in2[33];
    assign P[42] = in1[33] ^ in2[33];
    assign G[43] = in1[32] & in2[32];
    assign P[43] = in1[32] ^ in2[32];
    assign G[44] = in1[31] & in2[31];
    assign P[44] = in1[31] ^ in2[31];
    assign G[45] = in1[30] & in2[30];
    assign P[45] = in1[30] ^ in2[30];
    assign G[46] = in1[29] & in2[29];
    assign P[46] = in1[29] ^ in2[29];
    assign G[47] = in1[28] & in2[28];
    assign P[47] = in1[28] ^ in2[28];
    assign G[48] = in1[27] & in2[27];
    assign P[48] = in1[27] ^ in2[27];
    assign G[49] = in1[26] & in2[26];
    assign P[49] = in1[26] ^ in2[26];
    assign G[50] = in1[25] & in2[25];
    assign P[50] = in1[25] ^ in2[25];
    assign G[51] = in1[24] & in2[24];
    assign P[51] = in1[24] ^ in2[24];
    assign G[52] = in1[23] & in2[23];
    assign P[52] = in1[23] ^ in2[23];
    assign G[53] = in1[22] & in2[22];
    assign P[53] = in1[22] ^ in2[22];
    assign G[54] = in1[21] & in2[21];
    assign P[54] = in1[21] ^ in2[21];
    assign G[55] = in1[20] & in2[20];
    assign P[55] = in1[20] ^ in2[20];
    assign G[56] = in1[19] & in2[19];
    assign P[56] = in1[19] ^ in2[19];
    assign G[57] = in1[18] & in2[18];
    assign P[57] = in1[18] ^ in2[18];
    assign G[58] = in1[17] & in2[17];
    assign P[58] = in1[17] ^ in2[17];
    assign G[59] = in1[16] & in2[16];
    assign P[59] = in1[16] ^ in2[16];
    assign G[60] = in1[15] & in2[15];
    assign P[60] = in1[15] ^ in2[15];
    assign G[61] = in1[14] & in2[14];
    assign P[61] = in1[14] ^ in2[14];
    assign G[62] = in1[13] & in2[13];
    assign P[62] = in1[13] ^ in2[13];
    assign G[63] = in1[12] & in2[12];
    assign P[63] = in1[12] ^ in2[12];
    assign G[64] = in1[11] & in2[11];
    assign P[64] = in1[11] ^ in2[11];
    assign G[65] = in1[10] & in2[10];
    assign P[65] = in1[10] ^ in2[10];
    assign G[66] = in1[9] & in2[9];
    assign P[66] = in1[9] ^ in2[9];
    assign G[67] = in1[8] & in2[8];
    assign P[67] = in1[8] ^ in2[8];
    assign G[68] = in1[7] & in2[7];
    assign P[68] = in1[7] ^ in2[7];
    assign G[69] = in1[6] & in2[6];
    assign P[69] = in1[6] ^ in2[6];
    assign G[70] = in1[5] & in2[5];
    assign P[70] = in1[5] ^ in2[5];
    assign G[71] = in1[4] & in2[4];
    assign P[71] = in1[4] ^ in2[4];
    assign G[72] = in1[3] & in2[3];
    assign P[72] = in1[3] ^ in2[3];
    assign G[73] = in1[2] & in2[2];
    assign P[73] = in1[2] ^ in2[2];
    assign G[74] = in1[1] & in2[1];
    assign P[74] = in1[1] ^ in2[1];
    assign G[75] = in1[0] & in2[0];
    assign P[75] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign cout = G[75] | (P[75] & C[75]);
    assign sum = P ^ C;
endmodule

module CLA_75(output [74:0] sum, output cout, input [74:0] in1, input [74:0] in2);

    wire[74:0] G;
    wire[74:0] C;
    wire[74:0] P;

    assign G[0] = in1[74] & in2[74];
    assign P[0] = in1[74] ^ in2[74];
    assign G[1] = in1[73] & in2[73];
    assign P[1] = in1[73] ^ in2[73];
    assign G[2] = in1[72] & in2[72];
    assign P[2] = in1[72] ^ in2[72];
    assign G[3] = in1[71] & in2[71];
    assign P[3] = in1[71] ^ in2[71];
    assign G[4] = in1[70] & in2[70];
    assign P[4] = in1[70] ^ in2[70];
    assign G[5] = in1[69] & in2[69];
    assign P[5] = in1[69] ^ in2[69];
    assign G[6] = in1[68] & in2[68];
    assign P[6] = in1[68] ^ in2[68];
    assign G[7] = in1[67] & in2[67];
    assign P[7] = in1[67] ^ in2[67];
    assign G[8] = in1[66] & in2[66];
    assign P[8] = in1[66] ^ in2[66];
    assign G[9] = in1[65] & in2[65];
    assign P[9] = in1[65] ^ in2[65];
    assign G[10] = in1[64] & in2[64];
    assign P[10] = in1[64] ^ in2[64];
    assign G[11] = in1[63] & in2[63];
    assign P[11] = in1[63] ^ in2[63];
    assign G[12] = in1[62] & in2[62];
    assign P[12] = in1[62] ^ in2[62];
    assign G[13] = in1[61] & in2[61];
    assign P[13] = in1[61] ^ in2[61];
    assign G[14] = in1[60] & in2[60];
    assign P[14] = in1[60] ^ in2[60];
    assign G[15] = in1[59] & in2[59];
    assign P[15] = in1[59] ^ in2[59];
    assign G[16] = in1[58] & in2[58];
    assign P[16] = in1[58] ^ in2[58];
    assign G[17] = in1[57] & in2[57];
    assign P[17] = in1[57] ^ in2[57];
    assign G[18] = in1[56] & in2[56];
    assign P[18] = in1[56] ^ in2[56];
    assign G[19] = in1[55] & in2[55];
    assign P[19] = in1[55] ^ in2[55];
    assign G[20] = in1[54] & in2[54];
    assign P[20] = in1[54] ^ in2[54];
    assign G[21] = in1[53] & in2[53];
    assign P[21] = in1[53] ^ in2[53];
    assign G[22] = in1[52] & in2[52];
    assign P[22] = in1[52] ^ in2[52];
    assign G[23] = in1[51] & in2[51];
    assign P[23] = in1[51] ^ in2[51];
    assign G[24] = in1[50] & in2[50];
    assign P[24] = in1[50] ^ in2[50];
    assign G[25] = in1[49] & in2[49];
    assign P[25] = in1[49] ^ in2[49];
    assign G[26] = in1[48] & in2[48];
    assign P[26] = in1[48] ^ in2[48];
    assign G[27] = in1[47] & in2[47];
    assign P[27] = in1[47] ^ in2[47];
    assign G[28] = in1[46] & in2[46];
    assign P[28] = in1[46] ^ in2[46];
    assign G[29] = in1[45] & in2[45];
    assign P[29] = in1[45] ^ in2[45];
    assign G[30] = in1[44] & in2[44];
    assign P[30] = in1[44] ^ in2[44];
    assign G[31] = in1[43] & in2[43];
    assign P[31] = in1[43] ^ in2[43];
    assign G[32] = in1[42] & in2[42];
    assign P[32] = in1[42] ^ in2[42];
    assign G[33] = in1[41] & in2[41];
    assign P[33] = in1[41] ^ in2[41];
    assign G[34] = in1[40] & in2[40];
    assign P[34] = in1[40] ^ in2[40];
    assign G[35] = in1[39] & in2[39];
    assign P[35] = in1[39] ^ in2[39];
    assign G[36] = in1[38] & in2[38];
    assign P[36] = in1[38] ^ in2[38];
    assign G[37] = in1[37] & in2[37];
    assign P[37] = in1[37] ^ in2[37];
    assign G[38] = in1[36] & in2[36];
    assign P[38] = in1[36] ^ in2[36];
    assign G[39] = in1[35] & in2[35];
    assign P[39] = in1[35] ^ in2[35];
    assign G[40] = in1[34] & in2[34];
    assign P[40] = in1[34] ^ in2[34];
    assign G[41] = in1[33] & in2[33];
    assign P[41] = in1[33] ^ in2[33];
    assign G[42] = in1[32] & in2[32];
    assign P[42] = in1[32] ^ in2[32];
    assign G[43] = in1[31] & in2[31];
    assign P[43] = in1[31] ^ in2[31];
    assign G[44] = in1[30] & in2[30];
    assign P[44] = in1[30] ^ in2[30];
    assign G[45] = in1[29] & in2[29];
    assign P[45] = in1[29] ^ in2[29];
    assign G[46] = in1[28] & in2[28];
    assign P[46] = in1[28] ^ in2[28];
    assign G[47] = in1[27] & in2[27];
    assign P[47] = in1[27] ^ in2[27];
    assign G[48] = in1[26] & in2[26];
    assign P[48] = in1[26] ^ in2[26];
    assign G[49] = in1[25] & in2[25];
    assign P[49] = in1[25] ^ in2[25];
    assign G[50] = in1[24] & in2[24];
    assign P[50] = in1[24] ^ in2[24];
    assign G[51] = in1[23] & in2[23];
    assign P[51] = in1[23] ^ in2[23];
    assign G[52] = in1[22] & in2[22];
    assign P[52] = in1[22] ^ in2[22];
    assign G[53] = in1[21] & in2[21];
    assign P[53] = in1[21] ^ in2[21];
    assign G[54] = in1[20] & in2[20];
    assign P[54] = in1[20] ^ in2[20];
    assign G[55] = in1[19] & in2[19];
    assign P[55] = in1[19] ^ in2[19];
    assign G[56] = in1[18] & in2[18];
    assign P[56] = in1[18] ^ in2[18];
    assign G[57] = in1[17] & in2[17];
    assign P[57] = in1[17] ^ in2[17];
    assign G[58] = in1[16] & in2[16];
    assign P[58] = in1[16] ^ in2[16];
    assign G[59] = in1[15] & in2[15];
    assign P[59] = in1[15] ^ in2[15];
    assign G[60] = in1[14] & in2[14];
    assign P[60] = in1[14] ^ in2[14];
    assign G[61] = in1[13] & in2[13];
    assign P[61] = in1[13] ^ in2[13];
    assign G[62] = in1[12] & in2[12];
    assign P[62] = in1[12] ^ in2[12];
    assign G[63] = in1[11] & in2[11];
    assign P[63] = in1[11] ^ in2[11];
    assign G[64] = in1[10] & in2[10];
    assign P[64] = in1[10] ^ in2[10];
    assign G[65] = in1[9] & in2[9];
    assign P[65] = in1[9] ^ in2[9];
    assign G[66] = in1[8] & in2[8];
    assign P[66] = in1[8] ^ in2[8];
    assign G[67] = in1[7] & in2[7];
    assign P[67] = in1[7] ^ in2[7];
    assign G[68] = in1[6] & in2[6];
    assign P[68] = in1[6] ^ in2[6];
    assign G[69] = in1[5] & in2[5];
    assign P[69] = in1[5] ^ in2[5];
    assign G[70] = in1[4] & in2[4];
    assign P[70] = in1[4] ^ in2[4];
    assign G[71] = in1[3] & in2[3];
    assign P[71] = in1[3] ^ in2[3];
    assign G[72] = in1[2] & in2[2];
    assign P[72] = in1[2] ^ in2[2];
    assign G[73] = in1[1] & in2[1];
    assign P[73] = in1[1] ^ in2[1];
    assign G[74] = in1[0] & in2[0];
    assign P[74] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign cout = G[74] | (P[74] & C[74]);
    assign sum = P ^ C;
endmodule

module CLA_74(output [73:0] sum, output cout, input [73:0] in1, input [73:0] in2);

    wire[73:0] G;
    wire[73:0] C;
    wire[73:0] P;

    assign G[0] = in1[73] & in2[73];
    assign P[0] = in1[73] ^ in2[73];
    assign G[1] = in1[72] & in2[72];
    assign P[1] = in1[72] ^ in2[72];
    assign G[2] = in1[71] & in2[71];
    assign P[2] = in1[71] ^ in2[71];
    assign G[3] = in1[70] & in2[70];
    assign P[3] = in1[70] ^ in2[70];
    assign G[4] = in1[69] & in2[69];
    assign P[4] = in1[69] ^ in2[69];
    assign G[5] = in1[68] & in2[68];
    assign P[5] = in1[68] ^ in2[68];
    assign G[6] = in1[67] & in2[67];
    assign P[6] = in1[67] ^ in2[67];
    assign G[7] = in1[66] & in2[66];
    assign P[7] = in1[66] ^ in2[66];
    assign G[8] = in1[65] & in2[65];
    assign P[8] = in1[65] ^ in2[65];
    assign G[9] = in1[64] & in2[64];
    assign P[9] = in1[64] ^ in2[64];
    assign G[10] = in1[63] & in2[63];
    assign P[10] = in1[63] ^ in2[63];
    assign G[11] = in1[62] & in2[62];
    assign P[11] = in1[62] ^ in2[62];
    assign G[12] = in1[61] & in2[61];
    assign P[12] = in1[61] ^ in2[61];
    assign G[13] = in1[60] & in2[60];
    assign P[13] = in1[60] ^ in2[60];
    assign G[14] = in1[59] & in2[59];
    assign P[14] = in1[59] ^ in2[59];
    assign G[15] = in1[58] & in2[58];
    assign P[15] = in1[58] ^ in2[58];
    assign G[16] = in1[57] & in2[57];
    assign P[16] = in1[57] ^ in2[57];
    assign G[17] = in1[56] & in2[56];
    assign P[17] = in1[56] ^ in2[56];
    assign G[18] = in1[55] & in2[55];
    assign P[18] = in1[55] ^ in2[55];
    assign G[19] = in1[54] & in2[54];
    assign P[19] = in1[54] ^ in2[54];
    assign G[20] = in1[53] & in2[53];
    assign P[20] = in1[53] ^ in2[53];
    assign G[21] = in1[52] & in2[52];
    assign P[21] = in1[52] ^ in2[52];
    assign G[22] = in1[51] & in2[51];
    assign P[22] = in1[51] ^ in2[51];
    assign G[23] = in1[50] & in2[50];
    assign P[23] = in1[50] ^ in2[50];
    assign G[24] = in1[49] & in2[49];
    assign P[24] = in1[49] ^ in2[49];
    assign G[25] = in1[48] & in2[48];
    assign P[25] = in1[48] ^ in2[48];
    assign G[26] = in1[47] & in2[47];
    assign P[26] = in1[47] ^ in2[47];
    assign G[27] = in1[46] & in2[46];
    assign P[27] = in1[46] ^ in2[46];
    assign G[28] = in1[45] & in2[45];
    assign P[28] = in1[45] ^ in2[45];
    assign G[29] = in1[44] & in2[44];
    assign P[29] = in1[44] ^ in2[44];
    assign G[30] = in1[43] & in2[43];
    assign P[30] = in1[43] ^ in2[43];
    assign G[31] = in1[42] & in2[42];
    assign P[31] = in1[42] ^ in2[42];
    assign G[32] = in1[41] & in2[41];
    assign P[32] = in1[41] ^ in2[41];
    assign G[33] = in1[40] & in2[40];
    assign P[33] = in1[40] ^ in2[40];
    assign G[34] = in1[39] & in2[39];
    assign P[34] = in1[39] ^ in2[39];
    assign G[35] = in1[38] & in2[38];
    assign P[35] = in1[38] ^ in2[38];
    assign G[36] = in1[37] & in2[37];
    assign P[36] = in1[37] ^ in2[37];
    assign G[37] = in1[36] & in2[36];
    assign P[37] = in1[36] ^ in2[36];
    assign G[38] = in1[35] & in2[35];
    assign P[38] = in1[35] ^ in2[35];
    assign G[39] = in1[34] & in2[34];
    assign P[39] = in1[34] ^ in2[34];
    assign G[40] = in1[33] & in2[33];
    assign P[40] = in1[33] ^ in2[33];
    assign G[41] = in1[32] & in2[32];
    assign P[41] = in1[32] ^ in2[32];
    assign G[42] = in1[31] & in2[31];
    assign P[42] = in1[31] ^ in2[31];
    assign G[43] = in1[30] & in2[30];
    assign P[43] = in1[30] ^ in2[30];
    assign G[44] = in1[29] & in2[29];
    assign P[44] = in1[29] ^ in2[29];
    assign G[45] = in1[28] & in2[28];
    assign P[45] = in1[28] ^ in2[28];
    assign G[46] = in1[27] & in2[27];
    assign P[46] = in1[27] ^ in2[27];
    assign G[47] = in1[26] & in2[26];
    assign P[47] = in1[26] ^ in2[26];
    assign G[48] = in1[25] & in2[25];
    assign P[48] = in1[25] ^ in2[25];
    assign G[49] = in1[24] & in2[24];
    assign P[49] = in1[24] ^ in2[24];
    assign G[50] = in1[23] & in2[23];
    assign P[50] = in1[23] ^ in2[23];
    assign G[51] = in1[22] & in2[22];
    assign P[51] = in1[22] ^ in2[22];
    assign G[52] = in1[21] & in2[21];
    assign P[52] = in1[21] ^ in2[21];
    assign G[53] = in1[20] & in2[20];
    assign P[53] = in1[20] ^ in2[20];
    assign G[54] = in1[19] & in2[19];
    assign P[54] = in1[19] ^ in2[19];
    assign G[55] = in1[18] & in2[18];
    assign P[55] = in1[18] ^ in2[18];
    assign G[56] = in1[17] & in2[17];
    assign P[56] = in1[17] ^ in2[17];
    assign G[57] = in1[16] & in2[16];
    assign P[57] = in1[16] ^ in2[16];
    assign G[58] = in1[15] & in2[15];
    assign P[58] = in1[15] ^ in2[15];
    assign G[59] = in1[14] & in2[14];
    assign P[59] = in1[14] ^ in2[14];
    assign G[60] = in1[13] & in2[13];
    assign P[60] = in1[13] ^ in2[13];
    assign G[61] = in1[12] & in2[12];
    assign P[61] = in1[12] ^ in2[12];
    assign G[62] = in1[11] & in2[11];
    assign P[62] = in1[11] ^ in2[11];
    assign G[63] = in1[10] & in2[10];
    assign P[63] = in1[10] ^ in2[10];
    assign G[64] = in1[9] & in2[9];
    assign P[64] = in1[9] ^ in2[9];
    assign G[65] = in1[8] & in2[8];
    assign P[65] = in1[8] ^ in2[8];
    assign G[66] = in1[7] & in2[7];
    assign P[66] = in1[7] ^ in2[7];
    assign G[67] = in1[6] & in2[6];
    assign P[67] = in1[6] ^ in2[6];
    assign G[68] = in1[5] & in2[5];
    assign P[68] = in1[5] ^ in2[5];
    assign G[69] = in1[4] & in2[4];
    assign P[69] = in1[4] ^ in2[4];
    assign G[70] = in1[3] & in2[3];
    assign P[70] = in1[3] ^ in2[3];
    assign G[71] = in1[2] & in2[2];
    assign P[71] = in1[2] ^ in2[2];
    assign G[72] = in1[1] & in2[1];
    assign P[72] = in1[1] ^ in2[1];
    assign G[73] = in1[0] & in2[0];
    assign P[73] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign cout = G[73] | (P[73] & C[73]);
    assign sum = P ^ C;
endmodule

module CLA_73(output [72:0] sum, output cout, input [72:0] in1, input [72:0] in2);

    wire[72:0] G;
    wire[72:0] C;
    wire[72:0] P;

    assign G[0] = in1[72] & in2[72];
    assign P[0] = in1[72] ^ in2[72];
    assign G[1] = in1[71] & in2[71];
    assign P[1] = in1[71] ^ in2[71];
    assign G[2] = in1[70] & in2[70];
    assign P[2] = in1[70] ^ in2[70];
    assign G[3] = in1[69] & in2[69];
    assign P[3] = in1[69] ^ in2[69];
    assign G[4] = in1[68] & in2[68];
    assign P[4] = in1[68] ^ in2[68];
    assign G[5] = in1[67] & in2[67];
    assign P[5] = in1[67] ^ in2[67];
    assign G[6] = in1[66] & in2[66];
    assign P[6] = in1[66] ^ in2[66];
    assign G[7] = in1[65] & in2[65];
    assign P[7] = in1[65] ^ in2[65];
    assign G[8] = in1[64] & in2[64];
    assign P[8] = in1[64] ^ in2[64];
    assign G[9] = in1[63] & in2[63];
    assign P[9] = in1[63] ^ in2[63];
    assign G[10] = in1[62] & in2[62];
    assign P[10] = in1[62] ^ in2[62];
    assign G[11] = in1[61] & in2[61];
    assign P[11] = in1[61] ^ in2[61];
    assign G[12] = in1[60] & in2[60];
    assign P[12] = in1[60] ^ in2[60];
    assign G[13] = in1[59] & in2[59];
    assign P[13] = in1[59] ^ in2[59];
    assign G[14] = in1[58] & in2[58];
    assign P[14] = in1[58] ^ in2[58];
    assign G[15] = in1[57] & in2[57];
    assign P[15] = in1[57] ^ in2[57];
    assign G[16] = in1[56] & in2[56];
    assign P[16] = in1[56] ^ in2[56];
    assign G[17] = in1[55] & in2[55];
    assign P[17] = in1[55] ^ in2[55];
    assign G[18] = in1[54] & in2[54];
    assign P[18] = in1[54] ^ in2[54];
    assign G[19] = in1[53] & in2[53];
    assign P[19] = in1[53] ^ in2[53];
    assign G[20] = in1[52] & in2[52];
    assign P[20] = in1[52] ^ in2[52];
    assign G[21] = in1[51] & in2[51];
    assign P[21] = in1[51] ^ in2[51];
    assign G[22] = in1[50] & in2[50];
    assign P[22] = in1[50] ^ in2[50];
    assign G[23] = in1[49] & in2[49];
    assign P[23] = in1[49] ^ in2[49];
    assign G[24] = in1[48] & in2[48];
    assign P[24] = in1[48] ^ in2[48];
    assign G[25] = in1[47] & in2[47];
    assign P[25] = in1[47] ^ in2[47];
    assign G[26] = in1[46] & in2[46];
    assign P[26] = in1[46] ^ in2[46];
    assign G[27] = in1[45] & in2[45];
    assign P[27] = in1[45] ^ in2[45];
    assign G[28] = in1[44] & in2[44];
    assign P[28] = in1[44] ^ in2[44];
    assign G[29] = in1[43] & in2[43];
    assign P[29] = in1[43] ^ in2[43];
    assign G[30] = in1[42] & in2[42];
    assign P[30] = in1[42] ^ in2[42];
    assign G[31] = in1[41] & in2[41];
    assign P[31] = in1[41] ^ in2[41];
    assign G[32] = in1[40] & in2[40];
    assign P[32] = in1[40] ^ in2[40];
    assign G[33] = in1[39] & in2[39];
    assign P[33] = in1[39] ^ in2[39];
    assign G[34] = in1[38] & in2[38];
    assign P[34] = in1[38] ^ in2[38];
    assign G[35] = in1[37] & in2[37];
    assign P[35] = in1[37] ^ in2[37];
    assign G[36] = in1[36] & in2[36];
    assign P[36] = in1[36] ^ in2[36];
    assign G[37] = in1[35] & in2[35];
    assign P[37] = in1[35] ^ in2[35];
    assign G[38] = in1[34] & in2[34];
    assign P[38] = in1[34] ^ in2[34];
    assign G[39] = in1[33] & in2[33];
    assign P[39] = in1[33] ^ in2[33];
    assign G[40] = in1[32] & in2[32];
    assign P[40] = in1[32] ^ in2[32];
    assign G[41] = in1[31] & in2[31];
    assign P[41] = in1[31] ^ in2[31];
    assign G[42] = in1[30] & in2[30];
    assign P[42] = in1[30] ^ in2[30];
    assign G[43] = in1[29] & in2[29];
    assign P[43] = in1[29] ^ in2[29];
    assign G[44] = in1[28] & in2[28];
    assign P[44] = in1[28] ^ in2[28];
    assign G[45] = in1[27] & in2[27];
    assign P[45] = in1[27] ^ in2[27];
    assign G[46] = in1[26] & in2[26];
    assign P[46] = in1[26] ^ in2[26];
    assign G[47] = in1[25] & in2[25];
    assign P[47] = in1[25] ^ in2[25];
    assign G[48] = in1[24] & in2[24];
    assign P[48] = in1[24] ^ in2[24];
    assign G[49] = in1[23] & in2[23];
    assign P[49] = in1[23] ^ in2[23];
    assign G[50] = in1[22] & in2[22];
    assign P[50] = in1[22] ^ in2[22];
    assign G[51] = in1[21] & in2[21];
    assign P[51] = in1[21] ^ in2[21];
    assign G[52] = in1[20] & in2[20];
    assign P[52] = in1[20] ^ in2[20];
    assign G[53] = in1[19] & in2[19];
    assign P[53] = in1[19] ^ in2[19];
    assign G[54] = in1[18] & in2[18];
    assign P[54] = in1[18] ^ in2[18];
    assign G[55] = in1[17] & in2[17];
    assign P[55] = in1[17] ^ in2[17];
    assign G[56] = in1[16] & in2[16];
    assign P[56] = in1[16] ^ in2[16];
    assign G[57] = in1[15] & in2[15];
    assign P[57] = in1[15] ^ in2[15];
    assign G[58] = in1[14] & in2[14];
    assign P[58] = in1[14] ^ in2[14];
    assign G[59] = in1[13] & in2[13];
    assign P[59] = in1[13] ^ in2[13];
    assign G[60] = in1[12] & in2[12];
    assign P[60] = in1[12] ^ in2[12];
    assign G[61] = in1[11] & in2[11];
    assign P[61] = in1[11] ^ in2[11];
    assign G[62] = in1[10] & in2[10];
    assign P[62] = in1[10] ^ in2[10];
    assign G[63] = in1[9] & in2[9];
    assign P[63] = in1[9] ^ in2[9];
    assign G[64] = in1[8] & in2[8];
    assign P[64] = in1[8] ^ in2[8];
    assign G[65] = in1[7] & in2[7];
    assign P[65] = in1[7] ^ in2[7];
    assign G[66] = in1[6] & in2[6];
    assign P[66] = in1[6] ^ in2[6];
    assign G[67] = in1[5] & in2[5];
    assign P[67] = in1[5] ^ in2[5];
    assign G[68] = in1[4] & in2[4];
    assign P[68] = in1[4] ^ in2[4];
    assign G[69] = in1[3] & in2[3];
    assign P[69] = in1[3] ^ in2[3];
    assign G[70] = in1[2] & in2[2];
    assign P[70] = in1[2] ^ in2[2];
    assign G[71] = in1[1] & in2[1];
    assign P[71] = in1[1] ^ in2[1];
    assign G[72] = in1[0] & in2[0];
    assign P[72] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign cout = G[72] | (P[72] & C[72]);
    assign sum = P ^ C;
endmodule

module CLA_72(output [71:0] sum, output cout, input [71:0] in1, input [71:0] in2);

    wire[71:0] G;
    wire[71:0] C;
    wire[71:0] P;

    assign G[0] = in1[71] & in2[71];
    assign P[0] = in1[71] ^ in2[71];
    assign G[1] = in1[70] & in2[70];
    assign P[1] = in1[70] ^ in2[70];
    assign G[2] = in1[69] & in2[69];
    assign P[2] = in1[69] ^ in2[69];
    assign G[3] = in1[68] & in2[68];
    assign P[3] = in1[68] ^ in2[68];
    assign G[4] = in1[67] & in2[67];
    assign P[4] = in1[67] ^ in2[67];
    assign G[5] = in1[66] & in2[66];
    assign P[5] = in1[66] ^ in2[66];
    assign G[6] = in1[65] & in2[65];
    assign P[6] = in1[65] ^ in2[65];
    assign G[7] = in1[64] & in2[64];
    assign P[7] = in1[64] ^ in2[64];
    assign G[8] = in1[63] & in2[63];
    assign P[8] = in1[63] ^ in2[63];
    assign G[9] = in1[62] & in2[62];
    assign P[9] = in1[62] ^ in2[62];
    assign G[10] = in1[61] & in2[61];
    assign P[10] = in1[61] ^ in2[61];
    assign G[11] = in1[60] & in2[60];
    assign P[11] = in1[60] ^ in2[60];
    assign G[12] = in1[59] & in2[59];
    assign P[12] = in1[59] ^ in2[59];
    assign G[13] = in1[58] & in2[58];
    assign P[13] = in1[58] ^ in2[58];
    assign G[14] = in1[57] & in2[57];
    assign P[14] = in1[57] ^ in2[57];
    assign G[15] = in1[56] & in2[56];
    assign P[15] = in1[56] ^ in2[56];
    assign G[16] = in1[55] & in2[55];
    assign P[16] = in1[55] ^ in2[55];
    assign G[17] = in1[54] & in2[54];
    assign P[17] = in1[54] ^ in2[54];
    assign G[18] = in1[53] & in2[53];
    assign P[18] = in1[53] ^ in2[53];
    assign G[19] = in1[52] & in2[52];
    assign P[19] = in1[52] ^ in2[52];
    assign G[20] = in1[51] & in2[51];
    assign P[20] = in1[51] ^ in2[51];
    assign G[21] = in1[50] & in2[50];
    assign P[21] = in1[50] ^ in2[50];
    assign G[22] = in1[49] & in2[49];
    assign P[22] = in1[49] ^ in2[49];
    assign G[23] = in1[48] & in2[48];
    assign P[23] = in1[48] ^ in2[48];
    assign G[24] = in1[47] & in2[47];
    assign P[24] = in1[47] ^ in2[47];
    assign G[25] = in1[46] & in2[46];
    assign P[25] = in1[46] ^ in2[46];
    assign G[26] = in1[45] & in2[45];
    assign P[26] = in1[45] ^ in2[45];
    assign G[27] = in1[44] & in2[44];
    assign P[27] = in1[44] ^ in2[44];
    assign G[28] = in1[43] & in2[43];
    assign P[28] = in1[43] ^ in2[43];
    assign G[29] = in1[42] & in2[42];
    assign P[29] = in1[42] ^ in2[42];
    assign G[30] = in1[41] & in2[41];
    assign P[30] = in1[41] ^ in2[41];
    assign G[31] = in1[40] & in2[40];
    assign P[31] = in1[40] ^ in2[40];
    assign G[32] = in1[39] & in2[39];
    assign P[32] = in1[39] ^ in2[39];
    assign G[33] = in1[38] & in2[38];
    assign P[33] = in1[38] ^ in2[38];
    assign G[34] = in1[37] & in2[37];
    assign P[34] = in1[37] ^ in2[37];
    assign G[35] = in1[36] & in2[36];
    assign P[35] = in1[36] ^ in2[36];
    assign G[36] = in1[35] & in2[35];
    assign P[36] = in1[35] ^ in2[35];
    assign G[37] = in1[34] & in2[34];
    assign P[37] = in1[34] ^ in2[34];
    assign G[38] = in1[33] & in2[33];
    assign P[38] = in1[33] ^ in2[33];
    assign G[39] = in1[32] & in2[32];
    assign P[39] = in1[32] ^ in2[32];
    assign G[40] = in1[31] & in2[31];
    assign P[40] = in1[31] ^ in2[31];
    assign G[41] = in1[30] & in2[30];
    assign P[41] = in1[30] ^ in2[30];
    assign G[42] = in1[29] & in2[29];
    assign P[42] = in1[29] ^ in2[29];
    assign G[43] = in1[28] & in2[28];
    assign P[43] = in1[28] ^ in2[28];
    assign G[44] = in1[27] & in2[27];
    assign P[44] = in1[27] ^ in2[27];
    assign G[45] = in1[26] & in2[26];
    assign P[45] = in1[26] ^ in2[26];
    assign G[46] = in1[25] & in2[25];
    assign P[46] = in1[25] ^ in2[25];
    assign G[47] = in1[24] & in2[24];
    assign P[47] = in1[24] ^ in2[24];
    assign G[48] = in1[23] & in2[23];
    assign P[48] = in1[23] ^ in2[23];
    assign G[49] = in1[22] & in2[22];
    assign P[49] = in1[22] ^ in2[22];
    assign G[50] = in1[21] & in2[21];
    assign P[50] = in1[21] ^ in2[21];
    assign G[51] = in1[20] & in2[20];
    assign P[51] = in1[20] ^ in2[20];
    assign G[52] = in1[19] & in2[19];
    assign P[52] = in1[19] ^ in2[19];
    assign G[53] = in1[18] & in2[18];
    assign P[53] = in1[18] ^ in2[18];
    assign G[54] = in1[17] & in2[17];
    assign P[54] = in1[17] ^ in2[17];
    assign G[55] = in1[16] & in2[16];
    assign P[55] = in1[16] ^ in2[16];
    assign G[56] = in1[15] & in2[15];
    assign P[56] = in1[15] ^ in2[15];
    assign G[57] = in1[14] & in2[14];
    assign P[57] = in1[14] ^ in2[14];
    assign G[58] = in1[13] & in2[13];
    assign P[58] = in1[13] ^ in2[13];
    assign G[59] = in1[12] & in2[12];
    assign P[59] = in1[12] ^ in2[12];
    assign G[60] = in1[11] & in2[11];
    assign P[60] = in1[11] ^ in2[11];
    assign G[61] = in1[10] & in2[10];
    assign P[61] = in1[10] ^ in2[10];
    assign G[62] = in1[9] & in2[9];
    assign P[62] = in1[9] ^ in2[9];
    assign G[63] = in1[8] & in2[8];
    assign P[63] = in1[8] ^ in2[8];
    assign G[64] = in1[7] & in2[7];
    assign P[64] = in1[7] ^ in2[7];
    assign G[65] = in1[6] & in2[6];
    assign P[65] = in1[6] ^ in2[6];
    assign G[66] = in1[5] & in2[5];
    assign P[66] = in1[5] ^ in2[5];
    assign G[67] = in1[4] & in2[4];
    assign P[67] = in1[4] ^ in2[4];
    assign G[68] = in1[3] & in2[3];
    assign P[68] = in1[3] ^ in2[3];
    assign G[69] = in1[2] & in2[2];
    assign P[69] = in1[2] ^ in2[2];
    assign G[70] = in1[1] & in2[1];
    assign P[70] = in1[1] ^ in2[1];
    assign G[71] = in1[0] & in2[0];
    assign P[71] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign cout = G[71] | (P[71] & C[71]);
    assign sum = P ^ C;
endmodule

module CLA_71(output [70:0] sum, output cout, input [70:0] in1, input [70:0] in2);

    wire[70:0] G;
    wire[70:0] C;
    wire[70:0] P;

    assign G[0] = in1[70] & in2[70];
    assign P[0] = in1[70] ^ in2[70];
    assign G[1] = in1[69] & in2[69];
    assign P[1] = in1[69] ^ in2[69];
    assign G[2] = in1[68] & in2[68];
    assign P[2] = in1[68] ^ in2[68];
    assign G[3] = in1[67] & in2[67];
    assign P[3] = in1[67] ^ in2[67];
    assign G[4] = in1[66] & in2[66];
    assign P[4] = in1[66] ^ in2[66];
    assign G[5] = in1[65] & in2[65];
    assign P[5] = in1[65] ^ in2[65];
    assign G[6] = in1[64] & in2[64];
    assign P[6] = in1[64] ^ in2[64];
    assign G[7] = in1[63] & in2[63];
    assign P[7] = in1[63] ^ in2[63];
    assign G[8] = in1[62] & in2[62];
    assign P[8] = in1[62] ^ in2[62];
    assign G[9] = in1[61] & in2[61];
    assign P[9] = in1[61] ^ in2[61];
    assign G[10] = in1[60] & in2[60];
    assign P[10] = in1[60] ^ in2[60];
    assign G[11] = in1[59] & in2[59];
    assign P[11] = in1[59] ^ in2[59];
    assign G[12] = in1[58] & in2[58];
    assign P[12] = in1[58] ^ in2[58];
    assign G[13] = in1[57] & in2[57];
    assign P[13] = in1[57] ^ in2[57];
    assign G[14] = in1[56] & in2[56];
    assign P[14] = in1[56] ^ in2[56];
    assign G[15] = in1[55] & in2[55];
    assign P[15] = in1[55] ^ in2[55];
    assign G[16] = in1[54] & in2[54];
    assign P[16] = in1[54] ^ in2[54];
    assign G[17] = in1[53] & in2[53];
    assign P[17] = in1[53] ^ in2[53];
    assign G[18] = in1[52] & in2[52];
    assign P[18] = in1[52] ^ in2[52];
    assign G[19] = in1[51] & in2[51];
    assign P[19] = in1[51] ^ in2[51];
    assign G[20] = in1[50] & in2[50];
    assign P[20] = in1[50] ^ in2[50];
    assign G[21] = in1[49] & in2[49];
    assign P[21] = in1[49] ^ in2[49];
    assign G[22] = in1[48] & in2[48];
    assign P[22] = in1[48] ^ in2[48];
    assign G[23] = in1[47] & in2[47];
    assign P[23] = in1[47] ^ in2[47];
    assign G[24] = in1[46] & in2[46];
    assign P[24] = in1[46] ^ in2[46];
    assign G[25] = in1[45] & in2[45];
    assign P[25] = in1[45] ^ in2[45];
    assign G[26] = in1[44] & in2[44];
    assign P[26] = in1[44] ^ in2[44];
    assign G[27] = in1[43] & in2[43];
    assign P[27] = in1[43] ^ in2[43];
    assign G[28] = in1[42] & in2[42];
    assign P[28] = in1[42] ^ in2[42];
    assign G[29] = in1[41] & in2[41];
    assign P[29] = in1[41] ^ in2[41];
    assign G[30] = in1[40] & in2[40];
    assign P[30] = in1[40] ^ in2[40];
    assign G[31] = in1[39] & in2[39];
    assign P[31] = in1[39] ^ in2[39];
    assign G[32] = in1[38] & in2[38];
    assign P[32] = in1[38] ^ in2[38];
    assign G[33] = in1[37] & in2[37];
    assign P[33] = in1[37] ^ in2[37];
    assign G[34] = in1[36] & in2[36];
    assign P[34] = in1[36] ^ in2[36];
    assign G[35] = in1[35] & in2[35];
    assign P[35] = in1[35] ^ in2[35];
    assign G[36] = in1[34] & in2[34];
    assign P[36] = in1[34] ^ in2[34];
    assign G[37] = in1[33] & in2[33];
    assign P[37] = in1[33] ^ in2[33];
    assign G[38] = in1[32] & in2[32];
    assign P[38] = in1[32] ^ in2[32];
    assign G[39] = in1[31] & in2[31];
    assign P[39] = in1[31] ^ in2[31];
    assign G[40] = in1[30] & in2[30];
    assign P[40] = in1[30] ^ in2[30];
    assign G[41] = in1[29] & in2[29];
    assign P[41] = in1[29] ^ in2[29];
    assign G[42] = in1[28] & in2[28];
    assign P[42] = in1[28] ^ in2[28];
    assign G[43] = in1[27] & in2[27];
    assign P[43] = in1[27] ^ in2[27];
    assign G[44] = in1[26] & in2[26];
    assign P[44] = in1[26] ^ in2[26];
    assign G[45] = in1[25] & in2[25];
    assign P[45] = in1[25] ^ in2[25];
    assign G[46] = in1[24] & in2[24];
    assign P[46] = in1[24] ^ in2[24];
    assign G[47] = in1[23] & in2[23];
    assign P[47] = in1[23] ^ in2[23];
    assign G[48] = in1[22] & in2[22];
    assign P[48] = in1[22] ^ in2[22];
    assign G[49] = in1[21] & in2[21];
    assign P[49] = in1[21] ^ in2[21];
    assign G[50] = in1[20] & in2[20];
    assign P[50] = in1[20] ^ in2[20];
    assign G[51] = in1[19] & in2[19];
    assign P[51] = in1[19] ^ in2[19];
    assign G[52] = in1[18] & in2[18];
    assign P[52] = in1[18] ^ in2[18];
    assign G[53] = in1[17] & in2[17];
    assign P[53] = in1[17] ^ in2[17];
    assign G[54] = in1[16] & in2[16];
    assign P[54] = in1[16] ^ in2[16];
    assign G[55] = in1[15] & in2[15];
    assign P[55] = in1[15] ^ in2[15];
    assign G[56] = in1[14] & in2[14];
    assign P[56] = in1[14] ^ in2[14];
    assign G[57] = in1[13] & in2[13];
    assign P[57] = in1[13] ^ in2[13];
    assign G[58] = in1[12] & in2[12];
    assign P[58] = in1[12] ^ in2[12];
    assign G[59] = in1[11] & in2[11];
    assign P[59] = in1[11] ^ in2[11];
    assign G[60] = in1[10] & in2[10];
    assign P[60] = in1[10] ^ in2[10];
    assign G[61] = in1[9] & in2[9];
    assign P[61] = in1[9] ^ in2[9];
    assign G[62] = in1[8] & in2[8];
    assign P[62] = in1[8] ^ in2[8];
    assign G[63] = in1[7] & in2[7];
    assign P[63] = in1[7] ^ in2[7];
    assign G[64] = in1[6] & in2[6];
    assign P[64] = in1[6] ^ in2[6];
    assign G[65] = in1[5] & in2[5];
    assign P[65] = in1[5] ^ in2[5];
    assign G[66] = in1[4] & in2[4];
    assign P[66] = in1[4] ^ in2[4];
    assign G[67] = in1[3] & in2[3];
    assign P[67] = in1[3] ^ in2[3];
    assign G[68] = in1[2] & in2[2];
    assign P[68] = in1[2] ^ in2[2];
    assign G[69] = in1[1] & in2[1];
    assign P[69] = in1[1] ^ in2[1];
    assign G[70] = in1[0] & in2[0];
    assign P[70] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign cout = G[70] | (P[70] & C[70]);
    assign sum = P ^ C;
endmodule

module CLA_70(output [69:0] sum, output cout, input [69:0] in1, input [69:0] in2);

    wire[69:0] G;
    wire[69:0] C;
    wire[69:0] P;

    assign G[0] = in1[69] & in2[69];
    assign P[0] = in1[69] ^ in2[69];
    assign G[1] = in1[68] & in2[68];
    assign P[1] = in1[68] ^ in2[68];
    assign G[2] = in1[67] & in2[67];
    assign P[2] = in1[67] ^ in2[67];
    assign G[3] = in1[66] & in2[66];
    assign P[3] = in1[66] ^ in2[66];
    assign G[4] = in1[65] & in2[65];
    assign P[4] = in1[65] ^ in2[65];
    assign G[5] = in1[64] & in2[64];
    assign P[5] = in1[64] ^ in2[64];
    assign G[6] = in1[63] & in2[63];
    assign P[6] = in1[63] ^ in2[63];
    assign G[7] = in1[62] & in2[62];
    assign P[7] = in1[62] ^ in2[62];
    assign G[8] = in1[61] & in2[61];
    assign P[8] = in1[61] ^ in2[61];
    assign G[9] = in1[60] & in2[60];
    assign P[9] = in1[60] ^ in2[60];
    assign G[10] = in1[59] & in2[59];
    assign P[10] = in1[59] ^ in2[59];
    assign G[11] = in1[58] & in2[58];
    assign P[11] = in1[58] ^ in2[58];
    assign G[12] = in1[57] & in2[57];
    assign P[12] = in1[57] ^ in2[57];
    assign G[13] = in1[56] & in2[56];
    assign P[13] = in1[56] ^ in2[56];
    assign G[14] = in1[55] & in2[55];
    assign P[14] = in1[55] ^ in2[55];
    assign G[15] = in1[54] & in2[54];
    assign P[15] = in1[54] ^ in2[54];
    assign G[16] = in1[53] & in2[53];
    assign P[16] = in1[53] ^ in2[53];
    assign G[17] = in1[52] & in2[52];
    assign P[17] = in1[52] ^ in2[52];
    assign G[18] = in1[51] & in2[51];
    assign P[18] = in1[51] ^ in2[51];
    assign G[19] = in1[50] & in2[50];
    assign P[19] = in1[50] ^ in2[50];
    assign G[20] = in1[49] & in2[49];
    assign P[20] = in1[49] ^ in2[49];
    assign G[21] = in1[48] & in2[48];
    assign P[21] = in1[48] ^ in2[48];
    assign G[22] = in1[47] & in2[47];
    assign P[22] = in1[47] ^ in2[47];
    assign G[23] = in1[46] & in2[46];
    assign P[23] = in1[46] ^ in2[46];
    assign G[24] = in1[45] & in2[45];
    assign P[24] = in1[45] ^ in2[45];
    assign G[25] = in1[44] & in2[44];
    assign P[25] = in1[44] ^ in2[44];
    assign G[26] = in1[43] & in2[43];
    assign P[26] = in1[43] ^ in2[43];
    assign G[27] = in1[42] & in2[42];
    assign P[27] = in1[42] ^ in2[42];
    assign G[28] = in1[41] & in2[41];
    assign P[28] = in1[41] ^ in2[41];
    assign G[29] = in1[40] & in2[40];
    assign P[29] = in1[40] ^ in2[40];
    assign G[30] = in1[39] & in2[39];
    assign P[30] = in1[39] ^ in2[39];
    assign G[31] = in1[38] & in2[38];
    assign P[31] = in1[38] ^ in2[38];
    assign G[32] = in1[37] & in2[37];
    assign P[32] = in1[37] ^ in2[37];
    assign G[33] = in1[36] & in2[36];
    assign P[33] = in1[36] ^ in2[36];
    assign G[34] = in1[35] & in2[35];
    assign P[34] = in1[35] ^ in2[35];
    assign G[35] = in1[34] & in2[34];
    assign P[35] = in1[34] ^ in2[34];
    assign G[36] = in1[33] & in2[33];
    assign P[36] = in1[33] ^ in2[33];
    assign G[37] = in1[32] & in2[32];
    assign P[37] = in1[32] ^ in2[32];
    assign G[38] = in1[31] & in2[31];
    assign P[38] = in1[31] ^ in2[31];
    assign G[39] = in1[30] & in2[30];
    assign P[39] = in1[30] ^ in2[30];
    assign G[40] = in1[29] & in2[29];
    assign P[40] = in1[29] ^ in2[29];
    assign G[41] = in1[28] & in2[28];
    assign P[41] = in1[28] ^ in2[28];
    assign G[42] = in1[27] & in2[27];
    assign P[42] = in1[27] ^ in2[27];
    assign G[43] = in1[26] & in2[26];
    assign P[43] = in1[26] ^ in2[26];
    assign G[44] = in1[25] & in2[25];
    assign P[44] = in1[25] ^ in2[25];
    assign G[45] = in1[24] & in2[24];
    assign P[45] = in1[24] ^ in2[24];
    assign G[46] = in1[23] & in2[23];
    assign P[46] = in1[23] ^ in2[23];
    assign G[47] = in1[22] & in2[22];
    assign P[47] = in1[22] ^ in2[22];
    assign G[48] = in1[21] & in2[21];
    assign P[48] = in1[21] ^ in2[21];
    assign G[49] = in1[20] & in2[20];
    assign P[49] = in1[20] ^ in2[20];
    assign G[50] = in1[19] & in2[19];
    assign P[50] = in1[19] ^ in2[19];
    assign G[51] = in1[18] & in2[18];
    assign P[51] = in1[18] ^ in2[18];
    assign G[52] = in1[17] & in2[17];
    assign P[52] = in1[17] ^ in2[17];
    assign G[53] = in1[16] & in2[16];
    assign P[53] = in1[16] ^ in2[16];
    assign G[54] = in1[15] & in2[15];
    assign P[54] = in1[15] ^ in2[15];
    assign G[55] = in1[14] & in2[14];
    assign P[55] = in1[14] ^ in2[14];
    assign G[56] = in1[13] & in2[13];
    assign P[56] = in1[13] ^ in2[13];
    assign G[57] = in1[12] & in2[12];
    assign P[57] = in1[12] ^ in2[12];
    assign G[58] = in1[11] & in2[11];
    assign P[58] = in1[11] ^ in2[11];
    assign G[59] = in1[10] & in2[10];
    assign P[59] = in1[10] ^ in2[10];
    assign G[60] = in1[9] & in2[9];
    assign P[60] = in1[9] ^ in2[9];
    assign G[61] = in1[8] & in2[8];
    assign P[61] = in1[8] ^ in2[8];
    assign G[62] = in1[7] & in2[7];
    assign P[62] = in1[7] ^ in2[7];
    assign G[63] = in1[6] & in2[6];
    assign P[63] = in1[6] ^ in2[6];
    assign G[64] = in1[5] & in2[5];
    assign P[64] = in1[5] ^ in2[5];
    assign G[65] = in1[4] & in2[4];
    assign P[65] = in1[4] ^ in2[4];
    assign G[66] = in1[3] & in2[3];
    assign P[66] = in1[3] ^ in2[3];
    assign G[67] = in1[2] & in2[2];
    assign P[67] = in1[2] ^ in2[2];
    assign G[68] = in1[1] & in2[1];
    assign P[68] = in1[1] ^ in2[1];
    assign G[69] = in1[0] & in2[0];
    assign P[69] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign cout = G[69] | (P[69] & C[69]);
    assign sum = P ^ C;
endmodule

module CLA_69(output [68:0] sum, output cout, input [68:0] in1, input [68:0] in2);

    wire[68:0] G;
    wire[68:0] C;
    wire[68:0] P;

    assign G[0] = in1[68] & in2[68];
    assign P[0] = in1[68] ^ in2[68];
    assign G[1] = in1[67] & in2[67];
    assign P[1] = in1[67] ^ in2[67];
    assign G[2] = in1[66] & in2[66];
    assign P[2] = in1[66] ^ in2[66];
    assign G[3] = in1[65] & in2[65];
    assign P[3] = in1[65] ^ in2[65];
    assign G[4] = in1[64] & in2[64];
    assign P[4] = in1[64] ^ in2[64];
    assign G[5] = in1[63] & in2[63];
    assign P[5] = in1[63] ^ in2[63];
    assign G[6] = in1[62] & in2[62];
    assign P[6] = in1[62] ^ in2[62];
    assign G[7] = in1[61] & in2[61];
    assign P[7] = in1[61] ^ in2[61];
    assign G[8] = in1[60] & in2[60];
    assign P[8] = in1[60] ^ in2[60];
    assign G[9] = in1[59] & in2[59];
    assign P[9] = in1[59] ^ in2[59];
    assign G[10] = in1[58] & in2[58];
    assign P[10] = in1[58] ^ in2[58];
    assign G[11] = in1[57] & in2[57];
    assign P[11] = in1[57] ^ in2[57];
    assign G[12] = in1[56] & in2[56];
    assign P[12] = in1[56] ^ in2[56];
    assign G[13] = in1[55] & in2[55];
    assign P[13] = in1[55] ^ in2[55];
    assign G[14] = in1[54] & in2[54];
    assign P[14] = in1[54] ^ in2[54];
    assign G[15] = in1[53] & in2[53];
    assign P[15] = in1[53] ^ in2[53];
    assign G[16] = in1[52] & in2[52];
    assign P[16] = in1[52] ^ in2[52];
    assign G[17] = in1[51] & in2[51];
    assign P[17] = in1[51] ^ in2[51];
    assign G[18] = in1[50] & in2[50];
    assign P[18] = in1[50] ^ in2[50];
    assign G[19] = in1[49] & in2[49];
    assign P[19] = in1[49] ^ in2[49];
    assign G[20] = in1[48] & in2[48];
    assign P[20] = in1[48] ^ in2[48];
    assign G[21] = in1[47] & in2[47];
    assign P[21] = in1[47] ^ in2[47];
    assign G[22] = in1[46] & in2[46];
    assign P[22] = in1[46] ^ in2[46];
    assign G[23] = in1[45] & in2[45];
    assign P[23] = in1[45] ^ in2[45];
    assign G[24] = in1[44] & in2[44];
    assign P[24] = in1[44] ^ in2[44];
    assign G[25] = in1[43] & in2[43];
    assign P[25] = in1[43] ^ in2[43];
    assign G[26] = in1[42] & in2[42];
    assign P[26] = in1[42] ^ in2[42];
    assign G[27] = in1[41] & in2[41];
    assign P[27] = in1[41] ^ in2[41];
    assign G[28] = in1[40] & in2[40];
    assign P[28] = in1[40] ^ in2[40];
    assign G[29] = in1[39] & in2[39];
    assign P[29] = in1[39] ^ in2[39];
    assign G[30] = in1[38] & in2[38];
    assign P[30] = in1[38] ^ in2[38];
    assign G[31] = in1[37] & in2[37];
    assign P[31] = in1[37] ^ in2[37];
    assign G[32] = in1[36] & in2[36];
    assign P[32] = in1[36] ^ in2[36];
    assign G[33] = in1[35] & in2[35];
    assign P[33] = in1[35] ^ in2[35];
    assign G[34] = in1[34] & in2[34];
    assign P[34] = in1[34] ^ in2[34];
    assign G[35] = in1[33] & in2[33];
    assign P[35] = in1[33] ^ in2[33];
    assign G[36] = in1[32] & in2[32];
    assign P[36] = in1[32] ^ in2[32];
    assign G[37] = in1[31] & in2[31];
    assign P[37] = in1[31] ^ in2[31];
    assign G[38] = in1[30] & in2[30];
    assign P[38] = in1[30] ^ in2[30];
    assign G[39] = in1[29] & in2[29];
    assign P[39] = in1[29] ^ in2[29];
    assign G[40] = in1[28] & in2[28];
    assign P[40] = in1[28] ^ in2[28];
    assign G[41] = in1[27] & in2[27];
    assign P[41] = in1[27] ^ in2[27];
    assign G[42] = in1[26] & in2[26];
    assign P[42] = in1[26] ^ in2[26];
    assign G[43] = in1[25] & in2[25];
    assign P[43] = in1[25] ^ in2[25];
    assign G[44] = in1[24] & in2[24];
    assign P[44] = in1[24] ^ in2[24];
    assign G[45] = in1[23] & in2[23];
    assign P[45] = in1[23] ^ in2[23];
    assign G[46] = in1[22] & in2[22];
    assign P[46] = in1[22] ^ in2[22];
    assign G[47] = in1[21] & in2[21];
    assign P[47] = in1[21] ^ in2[21];
    assign G[48] = in1[20] & in2[20];
    assign P[48] = in1[20] ^ in2[20];
    assign G[49] = in1[19] & in2[19];
    assign P[49] = in1[19] ^ in2[19];
    assign G[50] = in1[18] & in2[18];
    assign P[50] = in1[18] ^ in2[18];
    assign G[51] = in1[17] & in2[17];
    assign P[51] = in1[17] ^ in2[17];
    assign G[52] = in1[16] & in2[16];
    assign P[52] = in1[16] ^ in2[16];
    assign G[53] = in1[15] & in2[15];
    assign P[53] = in1[15] ^ in2[15];
    assign G[54] = in1[14] & in2[14];
    assign P[54] = in1[14] ^ in2[14];
    assign G[55] = in1[13] & in2[13];
    assign P[55] = in1[13] ^ in2[13];
    assign G[56] = in1[12] & in2[12];
    assign P[56] = in1[12] ^ in2[12];
    assign G[57] = in1[11] & in2[11];
    assign P[57] = in1[11] ^ in2[11];
    assign G[58] = in1[10] & in2[10];
    assign P[58] = in1[10] ^ in2[10];
    assign G[59] = in1[9] & in2[9];
    assign P[59] = in1[9] ^ in2[9];
    assign G[60] = in1[8] & in2[8];
    assign P[60] = in1[8] ^ in2[8];
    assign G[61] = in1[7] & in2[7];
    assign P[61] = in1[7] ^ in2[7];
    assign G[62] = in1[6] & in2[6];
    assign P[62] = in1[6] ^ in2[6];
    assign G[63] = in1[5] & in2[5];
    assign P[63] = in1[5] ^ in2[5];
    assign G[64] = in1[4] & in2[4];
    assign P[64] = in1[4] ^ in2[4];
    assign G[65] = in1[3] & in2[3];
    assign P[65] = in1[3] ^ in2[3];
    assign G[66] = in1[2] & in2[2];
    assign P[66] = in1[2] ^ in2[2];
    assign G[67] = in1[1] & in2[1];
    assign P[67] = in1[1] ^ in2[1];
    assign G[68] = in1[0] & in2[0];
    assign P[68] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign cout = G[68] | (P[68] & C[68]);
    assign sum = P ^ C;
endmodule

module CLA_68(output [67:0] sum, output cout, input [67:0] in1, input [67:0] in2);

    wire[67:0] G;
    wire[67:0] C;
    wire[67:0] P;

    assign G[0] = in1[67] & in2[67];
    assign P[0] = in1[67] ^ in2[67];
    assign G[1] = in1[66] & in2[66];
    assign P[1] = in1[66] ^ in2[66];
    assign G[2] = in1[65] & in2[65];
    assign P[2] = in1[65] ^ in2[65];
    assign G[3] = in1[64] & in2[64];
    assign P[3] = in1[64] ^ in2[64];
    assign G[4] = in1[63] & in2[63];
    assign P[4] = in1[63] ^ in2[63];
    assign G[5] = in1[62] & in2[62];
    assign P[5] = in1[62] ^ in2[62];
    assign G[6] = in1[61] & in2[61];
    assign P[6] = in1[61] ^ in2[61];
    assign G[7] = in1[60] & in2[60];
    assign P[7] = in1[60] ^ in2[60];
    assign G[8] = in1[59] & in2[59];
    assign P[8] = in1[59] ^ in2[59];
    assign G[9] = in1[58] & in2[58];
    assign P[9] = in1[58] ^ in2[58];
    assign G[10] = in1[57] & in2[57];
    assign P[10] = in1[57] ^ in2[57];
    assign G[11] = in1[56] & in2[56];
    assign P[11] = in1[56] ^ in2[56];
    assign G[12] = in1[55] & in2[55];
    assign P[12] = in1[55] ^ in2[55];
    assign G[13] = in1[54] & in2[54];
    assign P[13] = in1[54] ^ in2[54];
    assign G[14] = in1[53] & in2[53];
    assign P[14] = in1[53] ^ in2[53];
    assign G[15] = in1[52] & in2[52];
    assign P[15] = in1[52] ^ in2[52];
    assign G[16] = in1[51] & in2[51];
    assign P[16] = in1[51] ^ in2[51];
    assign G[17] = in1[50] & in2[50];
    assign P[17] = in1[50] ^ in2[50];
    assign G[18] = in1[49] & in2[49];
    assign P[18] = in1[49] ^ in2[49];
    assign G[19] = in1[48] & in2[48];
    assign P[19] = in1[48] ^ in2[48];
    assign G[20] = in1[47] & in2[47];
    assign P[20] = in1[47] ^ in2[47];
    assign G[21] = in1[46] & in2[46];
    assign P[21] = in1[46] ^ in2[46];
    assign G[22] = in1[45] & in2[45];
    assign P[22] = in1[45] ^ in2[45];
    assign G[23] = in1[44] & in2[44];
    assign P[23] = in1[44] ^ in2[44];
    assign G[24] = in1[43] & in2[43];
    assign P[24] = in1[43] ^ in2[43];
    assign G[25] = in1[42] & in2[42];
    assign P[25] = in1[42] ^ in2[42];
    assign G[26] = in1[41] & in2[41];
    assign P[26] = in1[41] ^ in2[41];
    assign G[27] = in1[40] & in2[40];
    assign P[27] = in1[40] ^ in2[40];
    assign G[28] = in1[39] & in2[39];
    assign P[28] = in1[39] ^ in2[39];
    assign G[29] = in1[38] & in2[38];
    assign P[29] = in1[38] ^ in2[38];
    assign G[30] = in1[37] & in2[37];
    assign P[30] = in1[37] ^ in2[37];
    assign G[31] = in1[36] & in2[36];
    assign P[31] = in1[36] ^ in2[36];
    assign G[32] = in1[35] & in2[35];
    assign P[32] = in1[35] ^ in2[35];
    assign G[33] = in1[34] & in2[34];
    assign P[33] = in1[34] ^ in2[34];
    assign G[34] = in1[33] & in2[33];
    assign P[34] = in1[33] ^ in2[33];
    assign G[35] = in1[32] & in2[32];
    assign P[35] = in1[32] ^ in2[32];
    assign G[36] = in1[31] & in2[31];
    assign P[36] = in1[31] ^ in2[31];
    assign G[37] = in1[30] & in2[30];
    assign P[37] = in1[30] ^ in2[30];
    assign G[38] = in1[29] & in2[29];
    assign P[38] = in1[29] ^ in2[29];
    assign G[39] = in1[28] & in2[28];
    assign P[39] = in1[28] ^ in2[28];
    assign G[40] = in1[27] & in2[27];
    assign P[40] = in1[27] ^ in2[27];
    assign G[41] = in1[26] & in2[26];
    assign P[41] = in1[26] ^ in2[26];
    assign G[42] = in1[25] & in2[25];
    assign P[42] = in1[25] ^ in2[25];
    assign G[43] = in1[24] & in2[24];
    assign P[43] = in1[24] ^ in2[24];
    assign G[44] = in1[23] & in2[23];
    assign P[44] = in1[23] ^ in2[23];
    assign G[45] = in1[22] & in2[22];
    assign P[45] = in1[22] ^ in2[22];
    assign G[46] = in1[21] & in2[21];
    assign P[46] = in1[21] ^ in2[21];
    assign G[47] = in1[20] & in2[20];
    assign P[47] = in1[20] ^ in2[20];
    assign G[48] = in1[19] & in2[19];
    assign P[48] = in1[19] ^ in2[19];
    assign G[49] = in1[18] & in2[18];
    assign P[49] = in1[18] ^ in2[18];
    assign G[50] = in1[17] & in2[17];
    assign P[50] = in1[17] ^ in2[17];
    assign G[51] = in1[16] & in2[16];
    assign P[51] = in1[16] ^ in2[16];
    assign G[52] = in1[15] & in2[15];
    assign P[52] = in1[15] ^ in2[15];
    assign G[53] = in1[14] & in2[14];
    assign P[53] = in1[14] ^ in2[14];
    assign G[54] = in1[13] & in2[13];
    assign P[54] = in1[13] ^ in2[13];
    assign G[55] = in1[12] & in2[12];
    assign P[55] = in1[12] ^ in2[12];
    assign G[56] = in1[11] & in2[11];
    assign P[56] = in1[11] ^ in2[11];
    assign G[57] = in1[10] & in2[10];
    assign P[57] = in1[10] ^ in2[10];
    assign G[58] = in1[9] & in2[9];
    assign P[58] = in1[9] ^ in2[9];
    assign G[59] = in1[8] & in2[8];
    assign P[59] = in1[8] ^ in2[8];
    assign G[60] = in1[7] & in2[7];
    assign P[60] = in1[7] ^ in2[7];
    assign G[61] = in1[6] & in2[6];
    assign P[61] = in1[6] ^ in2[6];
    assign G[62] = in1[5] & in2[5];
    assign P[62] = in1[5] ^ in2[5];
    assign G[63] = in1[4] & in2[4];
    assign P[63] = in1[4] ^ in2[4];
    assign G[64] = in1[3] & in2[3];
    assign P[64] = in1[3] ^ in2[3];
    assign G[65] = in1[2] & in2[2];
    assign P[65] = in1[2] ^ in2[2];
    assign G[66] = in1[1] & in2[1];
    assign P[66] = in1[1] ^ in2[1];
    assign G[67] = in1[0] & in2[0];
    assign P[67] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign cout = G[67] | (P[67] & C[67]);
    assign sum = P ^ C;
endmodule

module CLA_67(output [66:0] sum, output cout, input [66:0] in1, input [66:0] in2);

    wire[66:0] G;
    wire[66:0] C;
    wire[66:0] P;

    assign G[0] = in1[66] & in2[66];
    assign P[0] = in1[66] ^ in2[66];
    assign G[1] = in1[65] & in2[65];
    assign P[1] = in1[65] ^ in2[65];
    assign G[2] = in1[64] & in2[64];
    assign P[2] = in1[64] ^ in2[64];
    assign G[3] = in1[63] & in2[63];
    assign P[3] = in1[63] ^ in2[63];
    assign G[4] = in1[62] & in2[62];
    assign P[4] = in1[62] ^ in2[62];
    assign G[5] = in1[61] & in2[61];
    assign P[5] = in1[61] ^ in2[61];
    assign G[6] = in1[60] & in2[60];
    assign P[6] = in1[60] ^ in2[60];
    assign G[7] = in1[59] & in2[59];
    assign P[7] = in1[59] ^ in2[59];
    assign G[8] = in1[58] & in2[58];
    assign P[8] = in1[58] ^ in2[58];
    assign G[9] = in1[57] & in2[57];
    assign P[9] = in1[57] ^ in2[57];
    assign G[10] = in1[56] & in2[56];
    assign P[10] = in1[56] ^ in2[56];
    assign G[11] = in1[55] & in2[55];
    assign P[11] = in1[55] ^ in2[55];
    assign G[12] = in1[54] & in2[54];
    assign P[12] = in1[54] ^ in2[54];
    assign G[13] = in1[53] & in2[53];
    assign P[13] = in1[53] ^ in2[53];
    assign G[14] = in1[52] & in2[52];
    assign P[14] = in1[52] ^ in2[52];
    assign G[15] = in1[51] & in2[51];
    assign P[15] = in1[51] ^ in2[51];
    assign G[16] = in1[50] & in2[50];
    assign P[16] = in1[50] ^ in2[50];
    assign G[17] = in1[49] & in2[49];
    assign P[17] = in1[49] ^ in2[49];
    assign G[18] = in1[48] & in2[48];
    assign P[18] = in1[48] ^ in2[48];
    assign G[19] = in1[47] & in2[47];
    assign P[19] = in1[47] ^ in2[47];
    assign G[20] = in1[46] & in2[46];
    assign P[20] = in1[46] ^ in2[46];
    assign G[21] = in1[45] & in2[45];
    assign P[21] = in1[45] ^ in2[45];
    assign G[22] = in1[44] & in2[44];
    assign P[22] = in1[44] ^ in2[44];
    assign G[23] = in1[43] & in2[43];
    assign P[23] = in1[43] ^ in2[43];
    assign G[24] = in1[42] & in2[42];
    assign P[24] = in1[42] ^ in2[42];
    assign G[25] = in1[41] & in2[41];
    assign P[25] = in1[41] ^ in2[41];
    assign G[26] = in1[40] & in2[40];
    assign P[26] = in1[40] ^ in2[40];
    assign G[27] = in1[39] & in2[39];
    assign P[27] = in1[39] ^ in2[39];
    assign G[28] = in1[38] & in2[38];
    assign P[28] = in1[38] ^ in2[38];
    assign G[29] = in1[37] & in2[37];
    assign P[29] = in1[37] ^ in2[37];
    assign G[30] = in1[36] & in2[36];
    assign P[30] = in1[36] ^ in2[36];
    assign G[31] = in1[35] & in2[35];
    assign P[31] = in1[35] ^ in2[35];
    assign G[32] = in1[34] & in2[34];
    assign P[32] = in1[34] ^ in2[34];
    assign G[33] = in1[33] & in2[33];
    assign P[33] = in1[33] ^ in2[33];
    assign G[34] = in1[32] & in2[32];
    assign P[34] = in1[32] ^ in2[32];
    assign G[35] = in1[31] & in2[31];
    assign P[35] = in1[31] ^ in2[31];
    assign G[36] = in1[30] & in2[30];
    assign P[36] = in1[30] ^ in2[30];
    assign G[37] = in1[29] & in2[29];
    assign P[37] = in1[29] ^ in2[29];
    assign G[38] = in1[28] & in2[28];
    assign P[38] = in1[28] ^ in2[28];
    assign G[39] = in1[27] & in2[27];
    assign P[39] = in1[27] ^ in2[27];
    assign G[40] = in1[26] & in2[26];
    assign P[40] = in1[26] ^ in2[26];
    assign G[41] = in1[25] & in2[25];
    assign P[41] = in1[25] ^ in2[25];
    assign G[42] = in1[24] & in2[24];
    assign P[42] = in1[24] ^ in2[24];
    assign G[43] = in1[23] & in2[23];
    assign P[43] = in1[23] ^ in2[23];
    assign G[44] = in1[22] & in2[22];
    assign P[44] = in1[22] ^ in2[22];
    assign G[45] = in1[21] & in2[21];
    assign P[45] = in1[21] ^ in2[21];
    assign G[46] = in1[20] & in2[20];
    assign P[46] = in1[20] ^ in2[20];
    assign G[47] = in1[19] & in2[19];
    assign P[47] = in1[19] ^ in2[19];
    assign G[48] = in1[18] & in2[18];
    assign P[48] = in1[18] ^ in2[18];
    assign G[49] = in1[17] & in2[17];
    assign P[49] = in1[17] ^ in2[17];
    assign G[50] = in1[16] & in2[16];
    assign P[50] = in1[16] ^ in2[16];
    assign G[51] = in1[15] & in2[15];
    assign P[51] = in1[15] ^ in2[15];
    assign G[52] = in1[14] & in2[14];
    assign P[52] = in1[14] ^ in2[14];
    assign G[53] = in1[13] & in2[13];
    assign P[53] = in1[13] ^ in2[13];
    assign G[54] = in1[12] & in2[12];
    assign P[54] = in1[12] ^ in2[12];
    assign G[55] = in1[11] & in2[11];
    assign P[55] = in1[11] ^ in2[11];
    assign G[56] = in1[10] & in2[10];
    assign P[56] = in1[10] ^ in2[10];
    assign G[57] = in1[9] & in2[9];
    assign P[57] = in1[9] ^ in2[9];
    assign G[58] = in1[8] & in2[8];
    assign P[58] = in1[8] ^ in2[8];
    assign G[59] = in1[7] & in2[7];
    assign P[59] = in1[7] ^ in2[7];
    assign G[60] = in1[6] & in2[6];
    assign P[60] = in1[6] ^ in2[6];
    assign G[61] = in1[5] & in2[5];
    assign P[61] = in1[5] ^ in2[5];
    assign G[62] = in1[4] & in2[4];
    assign P[62] = in1[4] ^ in2[4];
    assign G[63] = in1[3] & in2[3];
    assign P[63] = in1[3] ^ in2[3];
    assign G[64] = in1[2] & in2[2];
    assign P[64] = in1[2] ^ in2[2];
    assign G[65] = in1[1] & in2[1];
    assign P[65] = in1[1] ^ in2[1];
    assign G[66] = in1[0] & in2[0];
    assign P[66] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign cout = G[66] | (P[66] & C[66]);
    assign sum = P ^ C;
endmodule

module CLA_66(output [65:0] sum, output cout, input [65:0] in1, input [65:0] in2);

    wire[65:0] G;
    wire[65:0] C;
    wire[65:0] P;

    assign G[0] = in1[65] & in2[65];
    assign P[0] = in1[65] ^ in2[65];
    assign G[1] = in1[64] & in2[64];
    assign P[1] = in1[64] ^ in2[64];
    assign G[2] = in1[63] & in2[63];
    assign P[2] = in1[63] ^ in2[63];
    assign G[3] = in1[62] & in2[62];
    assign P[3] = in1[62] ^ in2[62];
    assign G[4] = in1[61] & in2[61];
    assign P[4] = in1[61] ^ in2[61];
    assign G[5] = in1[60] & in2[60];
    assign P[5] = in1[60] ^ in2[60];
    assign G[6] = in1[59] & in2[59];
    assign P[6] = in1[59] ^ in2[59];
    assign G[7] = in1[58] & in2[58];
    assign P[7] = in1[58] ^ in2[58];
    assign G[8] = in1[57] & in2[57];
    assign P[8] = in1[57] ^ in2[57];
    assign G[9] = in1[56] & in2[56];
    assign P[9] = in1[56] ^ in2[56];
    assign G[10] = in1[55] & in2[55];
    assign P[10] = in1[55] ^ in2[55];
    assign G[11] = in1[54] & in2[54];
    assign P[11] = in1[54] ^ in2[54];
    assign G[12] = in1[53] & in2[53];
    assign P[12] = in1[53] ^ in2[53];
    assign G[13] = in1[52] & in2[52];
    assign P[13] = in1[52] ^ in2[52];
    assign G[14] = in1[51] & in2[51];
    assign P[14] = in1[51] ^ in2[51];
    assign G[15] = in1[50] & in2[50];
    assign P[15] = in1[50] ^ in2[50];
    assign G[16] = in1[49] & in2[49];
    assign P[16] = in1[49] ^ in2[49];
    assign G[17] = in1[48] & in2[48];
    assign P[17] = in1[48] ^ in2[48];
    assign G[18] = in1[47] & in2[47];
    assign P[18] = in1[47] ^ in2[47];
    assign G[19] = in1[46] & in2[46];
    assign P[19] = in1[46] ^ in2[46];
    assign G[20] = in1[45] & in2[45];
    assign P[20] = in1[45] ^ in2[45];
    assign G[21] = in1[44] & in2[44];
    assign P[21] = in1[44] ^ in2[44];
    assign G[22] = in1[43] & in2[43];
    assign P[22] = in1[43] ^ in2[43];
    assign G[23] = in1[42] & in2[42];
    assign P[23] = in1[42] ^ in2[42];
    assign G[24] = in1[41] & in2[41];
    assign P[24] = in1[41] ^ in2[41];
    assign G[25] = in1[40] & in2[40];
    assign P[25] = in1[40] ^ in2[40];
    assign G[26] = in1[39] & in2[39];
    assign P[26] = in1[39] ^ in2[39];
    assign G[27] = in1[38] & in2[38];
    assign P[27] = in1[38] ^ in2[38];
    assign G[28] = in1[37] & in2[37];
    assign P[28] = in1[37] ^ in2[37];
    assign G[29] = in1[36] & in2[36];
    assign P[29] = in1[36] ^ in2[36];
    assign G[30] = in1[35] & in2[35];
    assign P[30] = in1[35] ^ in2[35];
    assign G[31] = in1[34] & in2[34];
    assign P[31] = in1[34] ^ in2[34];
    assign G[32] = in1[33] & in2[33];
    assign P[32] = in1[33] ^ in2[33];
    assign G[33] = in1[32] & in2[32];
    assign P[33] = in1[32] ^ in2[32];
    assign G[34] = in1[31] & in2[31];
    assign P[34] = in1[31] ^ in2[31];
    assign G[35] = in1[30] & in2[30];
    assign P[35] = in1[30] ^ in2[30];
    assign G[36] = in1[29] & in2[29];
    assign P[36] = in1[29] ^ in2[29];
    assign G[37] = in1[28] & in2[28];
    assign P[37] = in1[28] ^ in2[28];
    assign G[38] = in1[27] & in2[27];
    assign P[38] = in1[27] ^ in2[27];
    assign G[39] = in1[26] & in2[26];
    assign P[39] = in1[26] ^ in2[26];
    assign G[40] = in1[25] & in2[25];
    assign P[40] = in1[25] ^ in2[25];
    assign G[41] = in1[24] & in2[24];
    assign P[41] = in1[24] ^ in2[24];
    assign G[42] = in1[23] & in2[23];
    assign P[42] = in1[23] ^ in2[23];
    assign G[43] = in1[22] & in2[22];
    assign P[43] = in1[22] ^ in2[22];
    assign G[44] = in1[21] & in2[21];
    assign P[44] = in1[21] ^ in2[21];
    assign G[45] = in1[20] & in2[20];
    assign P[45] = in1[20] ^ in2[20];
    assign G[46] = in1[19] & in2[19];
    assign P[46] = in1[19] ^ in2[19];
    assign G[47] = in1[18] & in2[18];
    assign P[47] = in1[18] ^ in2[18];
    assign G[48] = in1[17] & in2[17];
    assign P[48] = in1[17] ^ in2[17];
    assign G[49] = in1[16] & in2[16];
    assign P[49] = in1[16] ^ in2[16];
    assign G[50] = in1[15] & in2[15];
    assign P[50] = in1[15] ^ in2[15];
    assign G[51] = in1[14] & in2[14];
    assign P[51] = in1[14] ^ in2[14];
    assign G[52] = in1[13] & in2[13];
    assign P[52] = in1[13] ^ in2[13];
    assign G[53] = in1[12] & in2[12];
    assign P[53] = in1[12] ^ in2[12];
    assign G[54] = in1[11] & in2[11];
    assign P[54] = in1[11] ^ in2[11];
    assign G[55] = in1[10] & in2[10];
    assign P[55] = in1[10] ^ in2[10];
    assign G[56] = in1[9] & in2[9];
    assign P[56] = in1[9] ^ in2[9];
    assign G[57] = in1[8] & in2[8];
    assign P[57] = in1[8] ^ in2[8];
    assign G[58] = in1[7] & in2[7];
    assign P[58] = in1[7] ^ in2[7];
    assign G[59] = in1[6] & in2[6];
    assign P[59] = in1[6] ^ in2[6];
    assign G[60] = in1[5] & in2[5];
    assign P[60] = in1[5] ^ in2[5];
    assign G[61] = in1[4] & in2[4];
    assign P[61] = in1[4] ^ in2[4];
    assign G[62] = in1[3] & in2[3];
    assign P[62] = in1[3] ^ in2[3];
    assign G[63] = in1[2] & in2[2];
    assign P[63] = in1[2] ^ in2[2];
    assign G[64] = in1[1] & in2[1];
    assign P[64] = in1[1] ^ in2[1];
    assign G[65] = in1[0] & in2[0];
    assign P[65] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign cout = G[65] | (P[65] & C[65]);
    assign sum = P ^ C;
endmodule

module CLA_65(output [64:0] sum, output cout, input [64:0] in1, input [64:0] in2);

    wire[64:0] G;
    wire[64:0] C;
    wire[64:0] P;

    assign G[0] = in1[64] & in2[64];
    assign P[0] = in1[64] ^ in2[64];
    assign G[1] = in1[63] & in2[63];
    assign P[1] = in1[63] ^ in2[63];
    assign G[2] = in1[62] & in2[62];
    assign P[2] = in1[62] ^ in2[62];
    assign G[3] = in1[61] & in2[61];
    assign P[3] = in1[61] ^ in2[61];
    assign G[4] = in1[60] & in2[60];
    assign P[4] = in1[60] ^ in2[60];
    assign G[5] = in1[59] & in2[59];
    assign P[5] = in1[59] ^ in2[59];
    assign G[6] = in1[58] & in2[58];
    assign P[6] = in1[58] ^ in2[58];
    assign G[7] = in1[57] & in2[57];
    assign P[7] = in1[57] ^ in2[57];
    assign G[8] = in1[56] & in2[56];
    assign P[8] = in1[56] ^ in2[56];
    assign G[9] = in1[55] & in2[55];
    assign P[9] = in1[55] ^ in2[55];
    assign G[10] = in1[54] & in2[54];
    assign P[10] = in1[54] ^ in2[54];
    assign G[11] = in1[53] & in2[53];
    assign P[11] = in1[53] ^ in2[53];
    assign G[12] = in1[52] & in2[52];
    assign P[12] = in1[52] ^ in2[52];
    assign G[13] = in1[51] & in2[51];
    assign P[13] = in1[51] ^ in2[51];
    assign G[14] = in1[50] & in2[50];
    assign P[14] = in1[50] ^ in2[50];
    assign G[15] = in1[49] & in2[49];
    assign P[15] = in1[49] ^ in2[49];
    assign G[16] = in1[48] & in2[48];
    assign P[16] = in1[48] ^ in2[48];
    assign G[17] = in1[47] & in2[47];
    assign P[17] = in1[47] ^ in2[47];
    assign G[18] = in1[46] & in2[46];
    assign P[18] = in1[46] ^ in2[46];
    assign G[19] = in1[45] & in2[45];
    assign P[19] = in1[45] ^ in2[45];
    assign G[20] = in1[44] & in2[44];
    assign P[20] = in1[44] ^ in2[44];
    assign G[21] = in1[43] & in2[43];
    assign P[21] = in1[43] ^ in2[43];
    assign G[22] = in1[42] & in2[42];
    assign P[22] = in1[42] ^ in2[42];
    assign G[23] = in1[41] & in2[41];
    assign P[23] = in1[41] ^ in2[41];
    assign G[24] = in1[40] & in2[40];
    assign P[24] = in1[40] ^ in2[40];
    assign G[25] = in1[39] & in2[39];
    assign P[25] = in1[39] ^ in2[39];
    assign G[26] = in1[38] & in2[38];
    assign P[26] = in1[38] ^ in2[38];
    assign G[27] = in1[37] & in2[37];
    assign P[27] = in1[37] ^ in2[37];
    assign G[28] = in1[36] & in2[36];
    assign P[28] = in1[36] ^ in2[36];
    assign G[29] = in1[35] & in2[35];
    assign P[29] = in1[35] ^ in2[35];
    assign G[30] = in1[34] & in2[34];
    assign P[30] = in1[34] ^ in2[34];
    assign G[31] = in1[33] & in2[33];
    assign P[31] = in1[33] ^ in2[33];
    assign G[32] = in1[32] & in2[32];
    assign P[32] = in1[32] ^ in2[32];
    assign G[33] = in1[31] & in2[31];
    assign P[33] = in1[31] ^ in2[31];
    assign G[34] = in1[30] & in2[30];
    assign P[34] = in1[30] ^ in2[30];
    assign G[35] = in1[29] & in2[29];
    assign P[35] = in1[29] ^ in2[29];
    assign G[36] = in1[28] & in2[28];
    assign P[36] = in1[28] ^ in2[28];
    assign G[37] = in1[27] & in2[27];
    assign P[37] = in1[27] ^ in2[27];
    assign G[38] = in1[26] & in2[26];
    assign P[38] = in1[26] ^ in2[26];
    assign G[39] = in1[25] & in2[25];
    assign P[39] = in1[25] ^ in2[25];
    assign G[40] = in1[24] & in2[24];
    assign P[40] = in1[24] ^ in2[24];
    assign G[41] = in1[23] & in2[23];
    assign P[41] = in1[23] ^ in2[23];
    assign G[42] = in1[22] & in2[22];
    assign P[42] = in1[22] ^ in2[22];
    assign G[43] = in1[21] & in2[21];
    assign P[43] = in1[21] ^ in2[21];
    assign G[44] = in1[20] & in2[20];
    assign P[44] = in1[20] ^ in2[20];
    assign G[45] = in1[19] & in2[19];
    assign P[45] = in1[19] ^ in2[19];
    assign G[46] = in1[18] & in2[18];
    assign P[46] = in1[18] ^ in2[18];
    assign G[47] = in1[17] & in2[17];
    assign P[47] = in1[17] ^ in2[17];
    assign G[48] = in1[16] & in2[16];
    assign P[48] = in1[16] ^ in2[16];
    assign G[49] = in1[15] & in2[15];
    assign P[49] = in1[15] ^ in2[15];
    assign G[50] = in1[14] & in2[14];
    assign P[50] = in1[14] ^ in2[14];
    assign G[51] = in1[13] & in2[13];
    assign P[51] = in1[13] ^ in2[13];
    assign G[52] = in1[12] & in2[12];
    assign P[52] = in1[12] ^ in2[12];
    assign G[53] = in1[11] & in2[11];
    assign P[53] = in1[11] ^ in2[11];
    assign G[54] = in1[10] & in2[10];
    assign P[54] = in1[10] ^ in2[10];
    assign G[55] = in1[9] & in2[9];
    assign P[55] = in1[9] ^ in2[9];
    assign G[56] = in1[8] & in2[8];
    assign P[56] = in1[8] ^ in2[8];
    assign G[57] = in1[7] & in2[7];
    assign P[57] = in1[7] ^ in2[7];
    assign G[58] = in1[6] & in2[6];
    assign P[58] = in1[6] ^ in2[6];
    assign G[59] = in1[5] & in2[5];
    assign P[59] = in1[5] ^ in2[5];
    assign G[60] = in1[4] & in2[4];
    assign P[60] = in1[4] ^ in2[4];
    assign G[61] = in1[3] & in2[3];
    assign P[61] = in1[3] ^ in2[3];
    assign G[62] = in1[2] & in2[2];
    assign P[62] = in1[2] ^ in2[2];
    assign G[63] = in1[1] & in2[1];
    assign P[63] = in1[1] ^ in2[1];
    assign G[64] = in1[0] & in2[0];
    assign P[64] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign cout = G[64] | (P[64] & C[64]);
    assign sum = P ^ C;
endmodule

module CLA_64(output [63:0] sum, output cout, input [63:0] in1, input [63:0] in2);

    wire[63:0] G;
    wire[63:0] C;
    wire[63:0] P;

    assign G[0] = in1[63] & in2[63];
    assign P[0] = in1[63] ^ in2[63];
    assign G[1] = in1[62] & in2[62];
    assign P[1] = in1[62] ^ in2[62];
    assign G[2] = in1[61] & in2[61];
    assign P[2] = in1[61] ^ in2[61];
    assign G[3] = in1[60] & in2[60];
    assign P[3] = in1[60] ^ in2[60];
    assign G[4] = in1[59] & in2[59];
    assign P[4] = in1[59] ^ in2[59];
    assign G[5] = in1[58] & in2[58];
    assign P[5] = in1[58] ^ in2[58];
    assign G[6] = in1[57] & in2[57];
    assign P[6] = in1[57] ^ in2[57];
    assign G[7] = in1[56] & in2[56];
    assign P[7] = in1[56] ^ in2[56];
    assign G[8] = in1[55] & in2[55];
    assign P[8] = in1[55] ^ in2[55];
    assign G[9] = in1[54] & in2[54];
    assign P[9] = in1[54] ^ in2[54];
    assign G[10] = in1[53] & in2[53];
    assign P[10] = in1[53] ^ in2[53];
    assign G[11] = in1[52] & in2[52];
    assign P[11] = in1[52] ^ in2[52];
    assign G[12] = in1[51] & in2[51];
    assign P[12] = in1[51] ^ in2[51];
    assign G[13] = in1[50] & in2[50];
    assign P[13] = in1[50] ^ in2[50];
    assign G[14] = in1[49] & in2[49];
    assign P[14] = in1[49] ^ in2[49];
    assign G[15] = in1[48] & in2[48];
    assign P[15] = in1[48] ^ in2[48];
    assign G[16] = in1[47] & in2[47];
    assign P[16] = in1[47] ^ in2[47];
    assign G[17] = in1[46] & in2[46];
    assign P[17] = in1[46] ^ in2[46];
    assign G[18] = in1[45] & in2[45];
    assign P[18] = in1[45] ^ in2[45];
    assign G[19] = in1[44] & in2[44];
    assign P[19] = in1[44] ^ in2[44];
    assign G[20] = in1[43] & in2[43];
    assign P[20] = in1[43] ^ in2[43];
    assign G[21] = in1[42] & in2[42];
    assign P[21] = in1[42] ^ in2[42];
    assign G[22] = in1[41] & in2[41];
    assign P[22] = in1[41] ^ in2[41];
    assign G[23] = in1[40] & in2[40];
    assign P[23] = in1[40] ^ in2[40];
    assign G[24] = in1[39] & in2[39];
    assign P[24] = in1[39] ^ in2[39];
    assign G[25] = in1[38] & in2[38];
    assign P[25] = in1[38] ^ in2[38];
    assign G[26] = in1[37] & in2[37];
    assign P[26] = in1[37] ^ in2[37];
    assign G[27] = in1[36] & in2[36];
    assign P[27] = in1[36] ^ in2[36];
    assign G[28] = in1[35] & in2[35];
    assign P[28] = in1[35] ^ in2[35];
    assign G[29] = in1[34] & in2[34];
    assign P[29] = in1[34] ^ in2[34];
    assign G[30] = in1[33] & in2[33];
    assign P[30] = in1[33] ^ in2[33];
    assign G[31] = in1[32] & in2[32];
    assign P[31] = in1[32] ^ in2[32];
    assign G[32] = in1[31] & in2[31];
    assign P[32] = in1[31] ^ in2[31];
    assign G[33] = in1[30] & in2[30];
    assign P[33] = in1[30] ^ in2[30];
    assign G[34] = in1[29] & in2[29];
    assign P[34] = in1[29] ^ in2[29];
    assign G[35] = in1[28] & in2[28];
    assign P[35] = in1[28] ^ in2[28];
    assign G[36] = in1[27] & in2[27];
    assign P[36] = in1[27] ^ in2[27];
    assign G[37] = in1[26] & in2[26];
    assign P[37] = in1[26] ^ in2[26];
    assign G[38] = in1[25] & in2[25];
    assign P[38] = in1[25] ^ in2[25];
    assign G[39] = in1[24] & in2[24];
    assign P[39] = in1[24] ^ in2[24];
    assign G[40] = in1[23] & in2[23];
    assign P[40] = in1[23] ^ in2[23];
    assign G[41] = in1[22] & in2[22];
    assign P[41] = in1[22] ^ in2[22];
    assign G[42] = in1[21] & in2[21];
    assign P[42] = in1[21] ^ in2[21];
    assign G[43] = in1[20] & in2[20];
    assign P[43] = in1[20] ^ in2[20];
    assign G[44] = in1[19] & in2[19];
    assign P[44] = in1[19] ^ in2[19];
    assign G[45] = in1[18] & in2[18];
    assign P[45] = in1[18] ^ in2[18];
    assign G[46] = in1[17] & in2[17];
    assign P[46] = in1[17] ^ in2[17];
    assign G[47] = in1[16] & in2[16];
    assign P[47] = in1[16] ^ in2[16];
    assign G[48] = in1[15] & in2[15];
    assign P[48] = in1[15] ^ in2[15];
    assign G[49] = in1[14] & in2[14];
    assign P[49] = in1[14] ^ in2[14];
    assign G[50] = in1[13] & in2[13];
    assign P[50] = in1[13] ^ in2[13];
    assign G[51] = in1[12] & in2[12];
    assign P[51] = in1[12] ^ in2[12];
    assign G[52] = in1[11] & in2[11];
    assign P[52] = in1[11] ^ in2[11];
    assign G[53] = in1[10] & in2[10];
    assign P[53] = in1[10] ^ in2[10];
    assign G[54] = in1[9] & in2[9];
    assign P[54] = in1[9] ^ in2[9];
    assign G[55] = in1[8] & in2[8];
    assign P[55] = in1[8] ^ in2[8];
    assign G[56] = in1[7] & in2[7];
    assign P[56] = in1[7] ^ in2[7];
    assign G[57] = in1[6] & in2[6];
    assign P[57] = in1[6] ^ in2[6];
    assign G[58] = in1[5] & in2[5];
    assign P[58] = in1[5] ^ in2[5];
    assign G[59] = in1[4] & in2[4];
    assign P[59] = in1[4] ^ in2[4];
    assign G[60] = in1[3] & in2[3];
    assign P[60] = in1[3] ^ in2[3];
    assign G[61] = in1[2] & in2[2];
    assign P[61] = in1[2] ^ in2[2];
    assign G[62] = in1[1] & in2[1];
    assign P[62] = in1[1] ^ in2[1];
    assign G[63] = in1[0] & in2[0];
    assign P[63] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign cout = G[63] | (P[63] & C[63]);
    assign sum = P ^ C;
endmodule

module CLA_63(output [62:0] sum, output cout, input [62:0] in1, input [62:0] in2);

    wire[62:0] G;
    wire[62:0] C;
    wire[62:0] P;

    assign G[0] = in1[62] & in2[62];
    assign P[0] = in1[62] ^ in2[62];
    assign G[1] = in1[61] & in2[61];
    assign P[1] = in1[61] ^ in2[61];
    assign G[2] = in1[60] & in2[60];
    assign P[2] = in1[60] ^ in2[60];
    assign G[3] = in1[59] & in2[59];
    assign P[3] = in1[59] ^ in2[59];
    assign G[4] = in1[58] & in2[58];
    assign P[4] = in1[58] ^ in2[58];
    assign G[5] = in1[57] & in2[57];
    assign P[5] = in1[57] ^ in2[57];
    assign G[6] = in1[56] & in2[56];
    assign P[6] = in1[56] ^ in2[56];
    assign G[7] = in1[55] & in2[55];
    assign P[7] = in1[55] ^ in2[55];
    assign G[8] = in1[54] & in2[54];
    assign P[8] = in1[54] ^ in2[54];
    assign G[9] = in1[53] & in2[53];
    assign P[9] = in1[53] ^ in2[53];
    assign G[10] = in1[52] & in2[52];
    assign P[10] = in1[52] ^ in2[52];
    assign G[11] = in1[51] & in2[51];
    assign P[11] = in1[51] ^ in2[51];
    assign G[12] = in1[50] & in2[50];
    assign P[12] = in1[50] ^ in2[50];
    assign G[13] = in1[49] & in2[49];
    assign P[13] = in1[49] ^ in2[49];
    assign G[14] = in1[48] & in2[48];
    assign P[14] = in1[48] ^ in2[48];
    assign G[15] = in1[47] & in2[47];
    assign P[15] = in1[47] ^ in2[47];
    assign G[16] = in1[46] & in2[46];
    assign P[16] = in1[46] ^ in2[46];
    assign G[17] = in1[45] & in2[45];
    assign P[17] = in1[45] ^ in2[45];
    assign G[18] = in1[44] & in2[44];
    assign P[18] = in1[44] ^ in2[44];
    assign G[19] = in1[43] & in2[43];
    assign P[19] = in1[43] ^ in2[43];
    assign G[20] = in1[42] & in2[42];
    assign P[20] = in1[42] ^ in2[42];
    assign G[21] = in1[41] & in2[41];
    assign P[21] = in1[41] ^ in2[41];
    assign G[22] = in1[40] & in2[40];
    assign P[22] = in1[40] ^ in2[40];
    assign G[23] = in1[39] & in2[39];
    assign P[23] = in1[39] ^ in2[39];
    assign G[24] = in1[38] & in2[38];
    assign P[24] = in1[38] ^ in2[38];
    assign G[25] = in1[37] & in2[37];
    assign P[25] = in1[37] ^ in2[37];
    assign G[26] = in1[36] & in2[36];
    assign P[26] = in1[36] ^ in2[36];
    assign G[27] = in1[35] & in2[35];
    assign P[27] = in1[35] ^ in2[35];
    assign G[28] = in1[34] & in2[34];
    assign P[28] = in1[34] ^ in2[34];
    assign G[29] = in1[33] & in2[33];
    assign P[29] = in1[33] ^ in2[33];
    assign G[30] = in1[32] & in2[32];
    assign P[30] = in1[32] ^ in2[32];
    assign G[31] = in1[31] & in2[31];
    assign P[31] = in1[31] ^ in2[31];
    assign G[32] = in1[30] & in2[30];
    assign P[32] = in1[30] ^ in2[30];
    assign G[33] = in1[29] & in2[29];
    assign P[33] = in1[29] ^ in2[29];
    assign G[34] = in1[28] & in2[28];
    assign P[34] = in1[28] ^ in2[28];
    assign G[35] = in1[27] & in2[27];
    assign P[35] = in1[27] ^ in2[27];
    assign G[36] = in1[26] & in2[26];
    assign P[36] = in1[26] ^ in2[26];
    assign G[37] = in1[25] & in2[25];
    assign P[37] = in1[25] ^ in2[25];
    assign G[38] = in1[24] & in2[24];
    assign P[38] = in1[24] ^ in2[24];
    assign G[39] = in1[23] & in2[23];
    assign P[39] = in1[23] ^ in2[23];
    assign G[40] = in1[22] & in2[22];
    assign P[40] = in1[22] ^ in2[22];
    assign G[41] = in1[21] & in2[21];
    assign P[41] = in1[21] ^ in2[21];
    assign G[42] = in1[20] & in2[20];
    assign P[42] = in1[20] ^ in2[20];
    assign G[43] = in1[19] & in2[19];
    assign P[43] = in1[19] ^ in2[19];
    assign G[44] = in1[18] & in2[18];
    assign P[44] = in1[18] ^ in2[18];
    assign G[45] = in1[17] & in2[17];
    assign P[45] = in1[17] ^ in2[17];
    assign G[46] = in1[16] & in2[16];
    assign P[46] = in1[16] ^ in2[16];
    assign G[47] = in1[15] & in2[15];
    assign P[47] = in1[15] ^ in2[15];
    assign G[48] = in1[14] & in2[14];
    assign P[48] = in1[14] ^ in2[14];
    assign G[49] = in1[13] & in2[13];
    assign P[49] = in1[13] ^ in2[13];
    assign G[50] = in1[12] & in2[12];
    assign P[50] = in1[12] ^ in2[12];
    assign G[51] = in1[11] & in2[11];
    assign P[51] = in1[11] ^ in2[11];
    assign G[52] = in1[10] & in2[10];
    assign P[52] = in1[10] ^ in2[10];
    assign G[53] = in1[9] & in2[9];
    assign P[53] = in1[9] ^ in2[9];
    assign G[54] = in1[8] & in2[8];
    assign P[54] = in1[8] ^ in2[8];
    assign G[55] = in1[7] & in2[7];
    assign P[55] = in1[7] ^ in2[7];
    assign G[56] = in1[6] & in2[6];
    assign P[56] = in1[6] ^ in2[6];
    assign G[57] = in1[5] & in2[5];
    assign P[57] = in1[5] ^ in2[5];
    assign G[58] = in1[4] & in2[4];
    assign P[58] = in1[4] ^ in2[4];
    assign G[59] = in1[3] & in2[3];
    assign P[59] = in1[3] ^ in2[3];
    assign G[60] = in1[2] & in2[2];
    assign P[60] = in1[2] ^ in2[2];
    assign G[61] = in1[1] & in2[1];
    assign P[61] = in1[1] ^ in2[1];
    assign G[62] = in1[0] & in2[0];
    assign P[62] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign cout = G[62] | (P[62] & C[62]);
    assign sum = P ^ C;
endmodule

module CLA_62(output [61:0] sum, output cout, input [61:0] in1, input [61:0] in2);

    wire[61:0] G;
    wire[61:0] C;
    wire[61:0] P;

    assign G[0] = in1[61] & in2[61];
    assign P[0] = in1[61] ^ in2[61];
    assign G[1] = in1[60] & in2[60];
    assign P[1] = in1[60] ^ in2[60];
    assign G[2] = in1[59] & in2[59];
    assign P[2] = in1[59] ^ in2[59];
    assign G[3] = in1[58] & in2[58];
    assign P[3] = in1[58] ^ in2[58];
    assign G[4] = in1[57] & in2[57];
    assign P[4] = in1[57] ^ in2[57];
    assign G[5] = in1[56] & in2[56];
    assign P[5] = in1[56] ^ in2[56];
    assign G[6] = in1[55] & in2[55];
    assign P[6] = in1[55] ^ in2[55];
    assign G[7] = in1[54] & in2[54];
    assign P[7] = in1[54] ^ in2[54];
    assign G[8] = in1[53] & in2[53];
    assign P[8] = in1[53] ^ in2[53];
    assign G[9] = in1[52] & in2[52];
    assign P[9] = in1[52] ^ in2[52];
    assign G[10] = in1[51] & in2[51];
    assign P[10] = in1[51] ^ in2[51];
    assign G[11] = in1[50] & in2[50];
    assign P[11] = in1[50] ^ in2[50];
    assign G[12] = in1[49] & in2[49];
    assign P[12] = in1[49] ^ in2[49];
    assign G[13] = in1[48] & in2[48];
    assign P[13] = in1[48] ^ in2[48];
    assign G[14] = in1[47] & in2[47];
    assign P[14] = in1[47] ^ in2[47];
    assign G[15] = in1[46] & in2[46];
    assign P[15] = in1[46] ^ in2[46];
    assign G[16] = in1[45] & in2[45];
    assign P[16] = in1[45] ^ in2[45];
    assign G[17] = in1[44] & in2[44];
    assign P[17] = in1[44] ^ in2[44];
    assign G[18] = in1[43] & in2[43];
    assign P[18] = in1[43] ^ in2[43];
    assign G[19] = in1[42] & in2[42];
    assign P[19] = in1[42] ^ in2[42];
    assign G[20] = in1[41] & in2[41];
    assign P[20] = in1[41] ^ in2[41];
    assign G[21] = in1[40] & in2[40];
    assign P[21] = in1[40] ^ in2[40];
    assign G[22] = in1[39] & in2[39];
    assign P[22] = in1[39] ^ in2[39];
    assign G[23] = in1[38] & in2[38];
    assign P[23] = in1[38] ^ in2[38];
    assign G[24] = in1[37] & in2[37];
    assign P[24] = in1[37] ^ in2[37];
    assign G[25] = in1[36] & in2[36];
    assign P[25] = in1[36] ^ in2[36];
    assign G[26] = in1[35] & in2[35];
    assign P[26] = in1[35] ^ in2[35];
    assign G[27] = in1[34] & in2[34];
    assign P[27] = in1[34] ^ in2[34];
    assign G[28] = in1[33] & in2[33];
    assign P[28] = in1[33] ^ in2[33];
    assign G[29] = in1[32] & in2[32];
    assign P[29] = in1[32] ^ in2[32];
    assign G[30] = in1[31] & in2[31];
    assign P[30] = in1[31] ^ in2[31];
    assign G[31] = in1[30] & in2[30];
    assign P[31] = in1[30] ^ in2[30];
    assign G[32] = in1[29] & in2[29];
    assign P[32] = in1[29] ^ in2[29];
    assign G[33] = in1[28] & in2[28];
    assign P[33] = in1[28] ^ in2[28];
    assign G[34] = in1[27] & in2[27];
    assign P[34] = in1[27] ^ in2[27];
    assign G[35] = in1[26] & in2[26];
    assign P[35] = in1[26] ^ in2[26];
    assign G[36] = in1[25] & in2[25];
    assign P[36] = in1[25] ^ in2[25];
    assign G[37] = in1[24] & in2[24];
    assign P[37] = in1[24] ^ in2[24];
    assign G[38] = in1[23] & in2[23];
    assign P[38] = in1[23] ^ in2[23];
    assign G[39] = in1[22] & in2[22];
    assign P[39] = in1[22] ^ in2[22];
    assign G[40] = in1[21] & in2[21];
    assign P[40] = in1[21] ^ in2[21];
    assign G[41] = in1[20] & in2[20];
    assign P[41] = in1[20] ^ in2[20];
    assign G[42] = in1[19] & in2[19];
    assign P[42] = in1[19] ^ in2[19];
    assign G[43] = in1[18] & in2[18];
    assign P[43] = in1[18] ^ in2[18];
    assign G[44] = in1[17] & in2[17];
    assign P[44] = in1[17] ^ in2[17];
    assign G[45] = in1[16] & in2[16];
    assign P[45] = in1[16] ^ in2[16];
    assign G[46] = in1[15] & in2[15];
    assign P[46] = in1[15] ^ in2[15];
    assign G[47] = in1[14] & in2[14];
    assign P[47] = in1[14] ^ in2[14];
    assign G[48] = in1[13] & in2[13];
    assign P[48] = in1[13] ^ in2[13];
    assign G[49] = in1[12] & in2[12];
    assign P[49] = in1[12] ^ in2[12];
    assign G[50] = in1[11] & in2[11];
    assign P[50] = in1[11] ^ in2[11];
    assign G[51] = in1[10] & in2[10];
    assign P[51] = in1[10] ^ in2[10];
    assign G[52] = in1[9] & in2[9];
    assign P[52] = in1[9] ^ in2[9];
    assign G[53] = in1[8] & in2[8];
    assign P[53] = in1[8] ^ in2[8];
    assign G[54] = in1[7] & in2[7];
    assign P[54] = in1[7] ^ in2[7];
    assign G[55] = in1[6] & in2[6];
    assign P[55] = in1[6] ^ in2[6];
    assign G[56] = in1[5] & in2[5];
    assign P[56] = in1[5] ^ in2[5];
    assign G[57] = in1[4] & in2[4];
    assign P[57] = in1[4] ^ in2[4];
    assign G[58] = in1[3] & in2[3];
    assign P[58] = in1[3] ^ in2[3];
    assign G[59] = in1[2] & in2[2];
    assign P[59] = in1[2] ^ in2[2];
    assign G[60] = in1[1] & in2[1];
    assign P[60] = in1[1] ^ in2[1];
    assign G[61] = in1[0] & in2[0];
    assign P[61] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign cout = G[61] | (P[61] & C[61]);
    assign sum = P ^ C;
endmodule

module CLA_61(output [60:0] sum, output cout, input [60:0] in1, input [60:0] in2);

    wire[60:0] G;
    wire[60:0] C;
    wire[60:0] P;

    assign G[0] = in1[60] & in2[60];
    assign P[0] = in1[60] ^ in2[60];
    assign G[1] = in1[59] & in2[59];
    assign P[1] = in1[59] ^ in2[59];
    assign G[2] = in1[58] & in2[58];
    assign P[2] = in1[58] ^ in2[58];
    assign G[3] = in1[57] & in2[57];
    assign P[3] = in1[57] ^ in2[57];
    assign G[4] = in1[56] & in2[56];
    assign P[4] = in1[56] ^ in2[56];
    assign G[5] = in1[55] & in2[55];
    assign P[5] = in1[55] ^ in2[55];
    assign G[6] = in1[54] & in2[54];
    assign P[6] = in1[54] ^ in2[54];
    assign G[7] = in1[53] & in2[53];
    assign P[7] = in1[53] ^ in2[53];
    assign G[8] = in1[52] & in2[52];
    assign P[8] = in1[52] ^ in2[52];
    assign G[9] = in1[51] & in2[51];
    assign P[9] = in1[51] ^ in2[51];
    assign G[10] = in1[50] & in2[50];
    assign P[10] = in1[50] ^ in2[50];
    assign G[11] = in1[49] & in2[49];
    assign P[11] = in1[49] ^ in2[49];
    assign G[12] = in1[48] & in2[48];
    assign P[12] = in1[48] ^ in2[48];
    assign G[13] = in1[47] & in2[47];
    assign P[13] = in1[47] ^ in2[47];
    assign G[14] = in1[46] & in2[46];
    assign P[14] = in1[46] ^ in2[46];
    assign G[15] = in1[45] & in2[45];
    assign P[15] = in1[45] ^ in2[45];
    assign G[16] = in1[44] & in2[44];
    assign P[16] = in1[44] ^ in2[44];
    assign G[17] = in1[43] & in2[43];
    assign P[17] = in1[43] ^ in2[43];
    assign G[18] = in1[42] & in2[42];
    assign P[18] = in1[42] ^ in2[42];
    assign G[19] = in1[41] & in2[41];
    assign P[19] = in1[41] ^ in2[41];
    assign G[20] = in1[40] & in2[40];
    assign P[20] = in1[40] ^ in2[40];
    assign G[21] = in1[39] & in2[39];
    assign P[21] = in1[39] ^ in2[39];
    assign G[22] = in1[38] & in2[38];
    assign P[22] = in1[38] ^ in2[38];
    assign G[23] = in1[37] & in2[37];
    assign P[23] = in1[37] ^ in2[37];
    assign G[24] = in1[36] & in2[36];
    assign P[24] = in1[36] ^ in2[36];
    assign G[25] = in1[35] & in2[35];
    assign P[25] = in1[35] ^ in2[35];
    assign G[26] = in1[34] & in2[34];
    assign P[26] = in1[34] ^ in2[34];
    assign G[27] = in1[33] & in2[33];
    assign P[27] = in1[33] ^ in2[33];
    assign G[28] = in1[32] & in2[32];
    assign P[28] = in1[32] ^ in2[32];
    assign G[29] = in1[31] & in2[31];
    assign P[29] = in1[31] ^ in2[31];
    assign G[30] = in1[30] & in2[30];
    assign P[30] = in1[30] ^ in2[30];
    assign G[31] = in1[29] & in2[29];
    assign P[31] = in1[29] ^ in2[29];
    assign G[32] = in1[28] & in2[28];
    assign P[32] = in1[28] ^ in2[28];
    assign G[33] = in1[27] & in2[27];
    assign P[33] = in1[27] ^ in2[27];
    assign G[34] = in1[26] & in2[26];
    assign P[34] = in1[26] ^ in2[26];
    assign G[35] = in1[25] & in2[25];
    assign P[35] = in1[25] ^ in2[25];
    assign G[36] = in1[24] & in2[24];
    assign P[36] = in1[24] ^ in2[24];
    assign G[37] = in1[23] & in2[23];
    assign P[37] = in1[23] ^ in2[23];
    assign G[38] = in1[22] & in2[22];
    assign P[38] = in1[22] ^ in2[22];
    assign G[39] = in1[21] & in2[21];
    assign P[39] = in1[21] ^ in2[21];
    assign G[40] = in1[20] & in2[20];
    assign P[40] = in1[20] ^ in2[20];
    assign G[41] = in1[19] & in2[19];
    assign P[41] = in1[19] ^ in2[19];
    assign G[42] = in1[18] & in2[18];
    assign P[42] = in1[18] ^ in2[18];
    assign G[43] = in1[17] & in2[17];
    assign P[43] = in1[17] ^ in2[17];
    assign G[44] = in1[16] & in2[16];
    assign P[44] = in1[16] ^ in2[16];
    assign G[45] = in1[15] & in2[15];
    assign P[45] = in1[15] ^ in2[15];
    assign G[46] = in1[14] & in2[14];
    assign P[46] = in1[14] ^ in2[14];
    assign G[47] = in1[13] & in2[13];
    assign P[47] = in1[13] ^ in2[13];
    assign G[48] = in1[12] & in2[12];
    assign P[48] = in1[12] ^ in2[12];
    assign G[49] = in1[11] & in2[11];
    assign P[49] = in1[11] ^ in2[11];
    assign G[50] = in1[10] & in2[10];
    assign P[50] = in1[10] ^ in2[10];
    assign G[51] = in1[9] & in2[9];
    assign P[51] = in1[9] ^ in2[9];
    assign G[52] = in1[8] & in2[8];
    assign P[52] = in1[8] ^ in2[8];
    assign G[53] = in1[7] & in2[7];
    assign P[53] = in1[7] ^ in2[7];
    assign G[54] = in1[6] & in2[6];
    assign P[54] = in1[6] ^ in2[6];
    assign G[55] = in1[5] & in2[5];
    assign P[55] = in1[5] ^ in2[5];
    assign G[56] = in1[4] & in2[4];
    assign P[56] = in1[4] ^ in2[4];
    assign G[57] = in1[3] & in2[3];
    assign P[57] = in1[3] ^ in2[3];
    assign G[58] = in1[2] & in2[2];
    assign P[58] = in1[2] ^ in2[2];
    assign G[59] = in1[1] & in2[1];
    assign P[59] = in1[1] ^ in2[1];
    assign G[60] = in1[0] & in2[0];
    assign P[60] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign cout = G[60] | (P[60] & C[60]);
    assign sum = P ^ C;
endmodule

module CLA_60(output [59:0] sum, output cout, input [59:0] in1, input [59:0] in2);

    wire[59:0] G;
    wire[59:0] C;
    wire[59:0] P;

    assign G[0] = in1[59] & in2[59];
    assign P[0] = in1[59] ^ in2[59];
    assign G[1] = in1[58] & in2[58];
    assign P[1] = in1[58] ^ in2[58];
    assign G[2] = in1[57] & in2[57];
    assign P[2] = in1[57] ^ in2[57];
    assign G[3] = in1[56] & in2[56];
    assign P[3] = in1[56] ^ in2[56];
    assign G[4] = in1[55] & in2[55];
    assign P[4] = in1[55] ^ in2[55];
    assign G[5] = in1[54] & in2[54];
    assign P[5] = in1[54] ^ in2[54];
    assign G[6] = in1[53] & in2[53];
    assign P[6] = in1[53] ^ in2[53];
    assign G[7] = in1[52] & in2[52];
    assign P[7] = in1[52] ^ in2[52];
    assign G[8] = in1[51] & in2[51];
    assign P[8] = in1[51] ^ in2[51];
    assign G[9] = in1[50] & in2[50];
    assign P[9] = in1[50] ^ in2[50];
    assign G[10] = in1[49] & in2[49];
    assign P[10] = in1[49] ^ in2[49];
    assign G[11] = in1[48] & in2[48];
    assign P[11] = in1[48] ^ in2[48];
    assign G[12] = in1[47] & in2[47];
    assign P[12] = in1[47] ^ in2[47];
    assign G[13] = in1[46] & in2[46];
    assign P[13] = in1[46] ^ in2[46];
    assign G[14] = in1[45] & in2[45];
    assign P[14] = in1[45] ^ in2[45];
    assign G[15] = in1[44] & in2[44];
    assign P[15] = in1[44] ^ in2[44];
    assign G[16] = in1[43] & in2[43];
    assign P[16] = in1[43] ^ in2[43];
    assign G[17] = in1[42] & in2[42];
    assign P[17] = in1[42] ^ in2[42];
    assign G[18] = in1[41] & in2[41];
    assign P[18] = in1[41] ^ in2[41];
    assign G[19] = in1[40] & in2[40];
    assign P[19] = in1[40] ^ in2[40];
    assign G[20] = in1[39] & in2[39];
    assign P[20] = in1[39] ^ in2[39];
    assign G[21] = in1[38] & in2[38];
    assign P[21] = in1[38] ^ in2[38];
    assign G[22] = in1[37] & in2[37];
    assign P[22] = in1[37] ^ in2[37];
    assign G[23] = in1[36] & in2[36];
    assign P[23] = in1[36] ^ in2[36];
    assign G[24] = in1[35] & in2[35];
    assign P[24] = in1[35] ^ in2[35];
    assign G[25] = in1[34] & in2[34];
    assign P[25] = in1[34] ^ in2[34];
    assign G[26] = in1[33] & in2[33];
    assign P[26] = in1[33] ^ in2[33];
    assign G[27] = in1[32] & in2[32];
    assign P[27] = in1[32] ^ in2[32];
    assign G[28] = in1[31] & in2[31];
    assign P[28] = in1[31] ^ in2[31];
    assign G[29] = in1[30] & in2[30];
    assign P[29] = in1[30] ^ in2[30];
    assign G[30] = in1[29] & in2[29];
    assign P[30] = in1[29] ^ in2[29];
    assign G[31] = in1[28] & in2[28];
    assign P[31] = in1[28] ^ in2[28];
    assign G[32] = in1[27] & in2[27];
    assign P[32] = in1[27] ^ in2[27];
    assign G[33] = in1[26] & in2[26];
    assign P[33] = in1[26] ^ in2[26];
    assign G[34] = in1[25] & in2[25];
    assign P[34] = in1[25] ^ in2[25];
    assign G[35] = in1[24] & in2[24];
    assign P[35] = in1[24] ^ in2[24];
    assign G[36] = in1[23] & in2[23];
    assign P[36] = in1[23] ^ in2[23];
    assign G[37] = in1[22] & in2[22];
    assign P[37] = in1[22] ^ in2[22];
    assign G[38] = in1[21] & in2[21];
    assign P[38] = in1[21] ^ in2[21];
    assign G[39] = in1[20] & in2[20];
    assign P[39] = in1[20] ^ in2[20];
    assign G[40] = in1[19] & in2[19];
    assign P[40] = in1[19] ^ in2[19];
    assign G[41] = in1[18] & in2[18];
    assign P[41] = in1[18] ^ in2[18];
    assign G[42] = in1[17] & in2[17];
    assign P[42] = in1[17] ^ in2[17];
    assign G[43] = in1[16] & in2[16];
    assign P[43] = in1[16] ^ in2[16];
    assign G[44] = in1[15] & in2[15];
    assign P[44] = in1[15] ^ in2[15];
    assign G[45] = in1[14] & in2[14];
    assign P[45] = in1[14] ^ in2[14];
    assign G[46] = in1[13] & in2[13];
    assign P[46] = in1[13] ^ in2[13];
    assign G[47] = in1[12] & in2[12];
    assign P[47] = in1[12] ^ in2[12];
    assign G[48] = in1[11] & in2[11];
    assign P[48] = in1[11] ^ in2[11];
    assign G[49] = in1[10] & in2[10];
    assign P[49] = in1[10] ^ in2[10];
    assign G[50] = in1[9] & in2[9];
    assign P[50] = in1[9] ^ in2[9];
    assign G[51] = in1[8] & in2[8];
    assign P[51] = in1[8] ^ in2[8];
    assign G[52] = in1[7] & in2[7];
    assign P[52] = in1[7] ^ in2[7];
    assign G[53] = in1[6] & in2[6];
    assign P[53] = in1[6] ^ in2[6];
    assign G[54] = in1[5] & in2[5];
    assign P[54] = in1[5] ^ in2[5];
    assign G[55] = in1[4] & in2[4];
    assign P[55] = in1[4] ^ in2[4];
    assign G[56] = in1[3] & in2[3];
    assign P[56] = in1[3] ^ in2[3];
    assign G[57] = in1[2] & in2[2];
    assign P[57] = in1[2] ^ in2[2];
    assign G[58] = in1[1] & in2[1];
    assign P[58] = in1[1] ^ in2[1];
    assign G[59] = in1[0] & in2[0];
    assign P[59] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign cout = G[59] | (P[59] & C[59]);
    assign sum = P ^ C;
endmodule

module CLA_59(output [58:0] sum, output cout, input [58:0] in1, input [58:0] in2);

    wire[58:0] G;
    wire[58:0] C;
    wire[58:0] P;

    assign G[0] = in1[58] & in2[58];
    assign P[0] = in1[58] ^ in2[58];
    assign G[1] = in1[57] & in2[57];
    assign P[1] = in1[57] ^ in2[57];
    assign G[2] = in1[56] & in2[56];
    assign P[2] = in1[56] ^ in2[56];
    assign G[3] = in1[55] & in2[55];
    assign P[3] = in1[55] ^ in2[55];
    assign G[4] = in1[54] & in2[54];
    assign P[4] = in1[54] ^ in2[54];
    assign G[5] = in1[53] & in2[53];
    assign P[5] = in1[53] ^ in2[53];
    assign G[6] = in1[52] & in2[52];
    assign P[6] = in1[52] ^ in2[52];
    assign G[7] = in1[51] & in2[51];
    assign P[7] = in1[51] ^ in2[51];
    assign G[8] = in1[50] & in2[50];
    assign P[8] = in1[50] ^ in2[50];
    assign G[9] = in1[49] & in2[49];
    assign P[9] = in1[49] ^ in2[49];
    assign G[10] = in1[48] & in2[48];
    assign P[10] = in1[48] ^ in2[48];
    assign G[11] = in1[47] & in2[47];
    assign P[11] = in1[47] ^ in2[47];
    assign G[12] = in1[46] & in2[46];
    assign P[12] = in1[46] ^ in2[46];
    assign G[13] = in1[45] & in2[45];
    assign P[13] = in1[45] ^ in2[45];
    assign G[14] = in1[44] & in2[44];
    assign P[14] = in1[44] ^ in2[44];
    assign G[15] = in1[43] & in2[43];
    assign P[15] = in1[43] ^ in2[43];
    assign G[16] = in1[42] & in2[42];
    assign P[16] = in1[42] ^ in2[42];
    assign G[17] = in1[41] & in2[41];
    assign P[17] = in1[41] ^ in2[41];
    assign G[18] = in1[40] & in2[40];
    assign P[18] = in1[40] ^ in2[40];
    assign G[19] = in1[39] & in2[39];
    assign P[19] = in1[39] ^ in2[39];
    assign G[20] = in1[38] & in2[38];
    assign P[20] = in1[38] ^ in2[38];
    assign G[21] = in1[37] & in2[37];
    assign P[21] = in1[37] ^ in2[37];
    assign G[22] = in1[36] & in2[36];
    assign P[22] = in1[36] ^ in2[36];
    assign G[23] = in1[35] & in2[35];
    assign P[23] = in1[35] ^ in2[35];
    assign G[24] = in1[34] & in2[34];
    assign P[24] = in1[34] ^ in2[34];
    assign G[25] = in1[33] & in2[33];
    assign P[25] = in1[33] ^ in2[33];
    assign G[26] = in1[32] & in2[32];
    assign P[26] = in1[32] ^ in2[32];
    assign G[27] = in1[31] & in2[31];
    assign P[27] = in1[31] ^ in2[31];
    assign G[28] = in1[30] & in2[30];
    assign P[28] = in1[30] ^ in2[30];
    assign G[29] = in1[29] & in2[29];
    assign P[29] = in1[29] ^ in2[29];
    assign G[30] = in1[28] & in2[28];
    assign P[30] = in1[28] ^ in2[28];
    assign G[31] = in1[27] & in2[27];
    assign P[31] = in1[27] ^ in2[27];
    assign G[32] = in1[26] & in2[26];
    assign P[32] = in1[26] ^ in2[26];
    assign G[33] = in1[25] & in2[25];
    assign P[33] = in1[25] ^ in2[25];
    assign G[34] = in1[24] & in2[24];
    assign P[34] = in1[24] ^ in2[24];
    assign G[35] = in1[23] & in2[23];
    assign P[35] = in1[23] ^ in2[23];
    assign G[36] = in1[22] & in2[22];
    assign P[36] = in1[22] ^ in2[22];
    assign G[37] = in1[21] & in2[21];
    assign P[37] = in1[21] ^ in2[21];
    assign G[38] = in1[20] & in2[20];
    assign P[38] = in1[20] ^ in2[20];
    assign G[39] = in1[19] & in2[19];
    assign P[39] = in1[19] ^ in2[19];
    assign G[40] = in1[18] & in2[18];
    assign P[40] = in1[18] ^ in2[18];
    assign G[41] = in1[17] & in2[17];
    assign P[41] = in1[17] ^ in2[17];
    assign G[42] = in1[16] & in2[16];
    assign P[42] = in1[16] ^ in2[16];
    assign G[43] = in1[15] & in2[15];
    assign P[43] = in1[15] ^ in2[15];
    assign G[44] = in1[14] & in2[14];
    assign P[44] = in1[14] ^ in2[14];
    assign G[45] = in1[13] & in2[13];
    assign P[45] = in1[13] ^ in2[13];
    assign G[46] = in1[12] & in2[12];
    assign P[46] = in1[12] ^ in2[12];
    assign G[47] = in1[11] & in2[11];
    assign P[47] = in1[11] ^ in2[11];
    assign G[48] = in1[10] & in2[10];
    assign P[48] = in1[10] ^ in2[10];
    assign G[49] = in1[9] & in2[9];
    assign P[49] = in1[9] ^ in2[9];
    assign G[50] = in1[8] & in2[8];
    assign P[50] = in1[8] ^ in2[8];
    assign G[51] = in1[7] & in2[7];
    assign P[51] = in1[7] ^ in2[7];
    assign G[52] = in1[6] & in2[6];
    assign P[52] = in1[6] ^ in2[6];
    assign G[53] = in1[5] & in2[5];
    assign P[53] = in1[5] ^ in2[5];
    assign G[54] = in1[4] & in2[4];
    assign P[54] = in1[4] ^ in2[4];
    assign G[55] = in1[3] & in2[3];
    assign P[55] = in1[3] ^ in2[3];
    assign G[56] = in1[2] & in2[2];
    assign P[56] = in1[2] ^ in2[2];
    assign G[57] = in1[1] & in2[1];
    assign P[57] = in1[1] ^ in2[1];
    assign G[58] = in1[0] & in2[0];
    assign P[58] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign cout = G[58] | (P[58] & C[58]);
    assign sum = P ^ C;
endmodule

module CLA_58(output [57:0] sum, output cout, input [57:0] in1, input [57:0] in2);

    wire[57:0] G;
    wire[57:0] C;
    wire[57:0] P;

    assign G[0] = in1[57] & in2[57];
    assign P[0] = in1[57] ^ in2[57];
    assign G[1] = in1[56] & in2[56];
    assign P[1] = in1[56] ^ in2[56];
    assign G[2] = in1[55] & in2[55];
    assign P[2] = in1[55] ^ in2[55];
    assign G[3] = in1[54] & in2[54];
    assign P[3] = in1[54] ^ in2[54];
    assign G[4] = in1[53] & in2[53];
    assign P[4] = in1[53] ^ in2[53];
    assign G[5] = in1[52] & in2[52];
    assign P[5] = in1[52] ^ in2[52];
    assign G[6] = in1[51] & in2[51];
    assign P[6] = in1[51] ^ in2[51];
    assign G[7] = in1[50] & in2[50];
    assign P[7] = in1[50] ^ in2[50];
    assign G[8] = in1[49] & in2[49];
    assign P[8] = in1[49] ^ in2[49];
    assign G[9] = in1[48] & in2[48];
    assign P[9] = in1[48] ^ in2[48];
    assign G[10] = in1[47] & in2[47];
    assign P[10] = in1[47] ^ in2[47];
    assign G[11] = in1[46] & in2[46];
    assign P[11] = in1[46] ^ in2[46];
    assign G[12] = in1[45] & in2[45];
    assign P[12] = in1[45] ^ in2[45];
    assign G[13] = in1[44] & in2[44];
    assign P[13] = in1[44] ^ in2[44];
    assign G[14] = in1[43] & in2[43];
    assign P[14] = in1[43] ^ in2[43];
    assign G[15] = in1[42] & in2[42];
    assign P[15] = in1[42] ^ in2[42];
    assign G[16] = in1[41] & in2[41];
    assign P[16] = in1[41] ^ in2[41];
    assign G[17] = in1[40] & in2[40];
    assign P[17] = in1[40] ^ in2[40];
    assign G[18] = in1[39] & in2[39];
    assign P[18] = in1[39] ^ in2[39];
    assign G[19] = in1[38] & in2[38];
    assign P[19] = in1[38] ^ in2[38];
    assign G[20] = in1[37] & in2[37];
    assign P[20] = in1[37] ^ in2[37];
    assign G[21] = in1[36] & in2[36];
    assign P[21] = in1[36] ^ in2[36];
    assign G[22] = in1[35] & in2[35];
    assign P[22] = in1[35] ^ in2[35];
    assign G[23] = in1[34] & in2[34];
    assign P[23] = in1[34] ^ in2[34];
    assign G[24] = in1[33] & in2[33];
    assign P[24] = in1[33] ^ in2[33];
    assign G[25] = in1[32] & in2[32];
    assign P[25] = in1[32] ^ in2[32];
    assign G[26] = in1[31] & in2[31];
    assign P[26] = in1[31] ^ in2[31];
    assign G[27] = in1[30] & in2[30];
    assign P[27] = in1[30] ^ in2[30];
    assign G[28] = in1[29] & in2[29];
    assign P[28] = in1[29] ^ in2[29];
    assign G[29] = in1[28] & in2[28];
    assign P[29] = in1[28] ^ in2[28];
    assign G[30] = in1[27] & in2[27];
    assign P[30] = in1[27] ^ in2[27];
    assign G[31] = in1[26] & in2[26];
    assign P[31] = in1[26] ^ in2[26];
    assign G[32] = in1[25] & in2[25];
    assign P[32] = in1[25] ^ in2[25];
    assign G[33] = in1[24] & in2[24];
    assign P[33] = in1[24] ^ in2[24];
    assign G[34] = in1[23] & in2[23];
    assign P[34] = in1[23] ^ in2[23];
    assign G[35] = in1[22] & in2[22];
    assign P[35] = in1[22] ^ in2[22];
    assign G[36] = in1[21] & in2[21];
    assign P[36] = in1[21] ^ in2[21];
    assign G[37] = in1[20] & in2[20];
    assign P[37] = in1[20] ^ in2[20];
    assign G[38] = in1[19] & in2[19];
    assign P[38] = in1[19] ^ in2[19];
    assign G[39] = in1[18] & in2[18];
    assign P[39] = in1[18] ^ in2[18];
    assign G[40] = in1[17] & in2[17];
    assign P[40] = in1[17] ^ in2[17];
    assign G[41] = in1[16] & in2[16];
    assign P[41] = in1[16] ^ in2[16];
    assign G[42] = in1[15] & in2[15];
    assign P[42] = in1[15] ^ in2[15];
    assign G[43] = in1[14] & in2[14];
    assign P[43] = in1[14] ^ in2[14];
    assign G[44] = in1[13] & in2[13];
    assign P[44] = in1[13] ^ in2[13];
    assign G[45] = in1[12] & in2[12];
    assign P[45] = in1[12] ^ in2[12];
    assign G[46] = in1[11] & in2[11];
    assign P[46] = in1[11] ^ in2[11];
    assign G[47] = in1[10] & in2[10];
    assign P[47] = in1[10] ^ in2[10];
    assign G[48] = in1[9] & in2[9];
    assign P[48] = in1[9] ^ in2[9];
    assign G[49] = in1[8] & in2[8];
    assign P[49] = in1[8] ^ in2[8];
    assign G[50] = in1[7] & in2[7];
    assign P[50] = in1[7] ^ in2[7];
    assign G[51] = in1[6] & in2[6];
    assign P[51] = in1[6] ^ in2[6];
    assign G[52] = in1[5] & in2[5];
    assign P[52] = in1[5] ^ in2[5];
    assign G[53] = in1[4] & in2[4];
    assign P[53] = in1[4] ^ in2[4];
    assign G[54] = in1[3] & in2[3];
    assign P[54] = in1[3] ^ in2[3];
    assign G[55] = in1[2] & in2[2];
    assign P[55] = in1[2] ^ in2[2];
    assign G[56] = in1[1] & in2[1];
    assign P[56] = in1[1] ^ in2[1];
    assign G[57] = in1[0] & in2[0];
    assign P[57] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign cout = G[57] | (P[57] & C[57]);
    assign sum = P ^ C;
endmodule

module CLA_57(output [56:0] sum, output cout, input [56:0] in1, input [56:0] in2);

    wire[56:0] G;
    wire[56:0] C;
    wire[56:0] P;

    assign G[0] = in1[56] & in2[56];
    assign P[0] = in1[56] ^ in2[56];
    assign G[1] = in1[55] & in2[55];
    assign P[1] = in1[55] ^ in2[55];
    assign G[2] = in1[54] & in2[54];
    assign P[2] = in1[54] ^ in2[54];
    assign G[3] = in1[53] & in2[53];
    assign P[3] = in1[53] ^ in2[53];
    assign G[4] = in1[52] & in2[52];
    assign P[4] = in1[52] ^ in2[52];
    assign G[5] = in1[51] & in2[51];
    assign P[5] = in1[51] ^ in2[51];
    assign G[6] = in1[50] & in2[50];
    assign P[6] = in1[50] ^ in2[50];
    assign G[7] = in1[49] & in2[49];
    assign P[7] = in1[49] ^ in2[49];
    assign G[8] = in1[48] & in2[48];
    assign P[8] = in1[48] ^ in2[48];
    assign G[9] = in1[47] & in2[47];
    assign P[9] = in1[47] ^ in2[47];
    assign G[10] = in1[46] & in2[46];
    assign P[10] = in1[46] ^ in2[46];
    assign G[11] = in1[45] & in2[45];
    assign P[11] = in1[45] ^ in2[45];
    assign G[12] = in1[44] & in2[44];
    assign P[12] = in1[44] ^ in2[44];
    assign G[13] = in1[43] & in2[43];
    assign P[13] = in1[43] ^ in2[43];
    assign G[14] = in1[42] & in2[42];
    assign P[14] = in1[42] ^ in2[42];
    assign G[15] = in1[41] & in2[41];
    assign P[15] = in1[41] ^ in2[41];
    assign G[16] = in1[40] & in2[40];
    assign P[16] = in1[40] ^ in2[40];
    assign G[17] = in1[39] & in2[39];
    assign P[17] = in1[39] ^ in2[39];
    assign G[18] = in1[38] & in2[38];
    assign P[18] = in1[38] ^ in2[38];
    assign G[19] = in1[37] & in2[37];
    assign P[19] = in1[37] ^ in2[37];
    assign G[20] = in1[36] & in2[36];
    assign P[20] = in1[36] ^ in2[36];
    assign G[21] = in1[35] & in2[35];
    assign P[21] = in1[35] ^ in2[35];
    assign G[22] = in1[34] & in2[34];
    assign P[22] = in1[34] ^ in2[34];
    assign G[23] = in1[33] & in2[33];
    assign P[23] = in1[33] ^ in2[33];
    assign G[24] = in1[32] & in2[32];
    assign P[24] = in1[32] ^ in2[32];
    assign G[25] = in1[31] & in2[31];
    assign P[25] = in1[31] ^ in2[31];
    assign G[26] = in1[30] & in2[30];
    assign P[26] = in1[30] ^ in2[30];
    assign G[27] = in1[29] & in2[29];
    assign P[27] = in1[29] ^ in2[29];
    assign G[28] = in1[28] & in2[28];
    assign P[28] = in1[28] ^ in2[28];
    assign G[29] = in1[27] & in2[27];
    assign P[29] = in1[27] ^ in2[27];
    assign G[30] = in1[26] & in2[26];
    assign P[30] = in1[26] ^ in2[26];
    assign G[31] = in1[25] & in2[25];
    assign P[31] = in1[25] ^ in2[25];
    assign G[32] = in1[24] & in2[24];
    assign P[32] = in1[24] ^ in2[24];
    assign G[33] = in1[23] & in2[23];
    assign P[33] = in1[23] ^ in2[23];
    assign G[34] = in1[22] & in2[22];
    assign P[34] = in1[22] ^ in2[22];
    assign G[35] = in1[21] & in2[21];
    assign P[35] = in1[21] ^ in2[21];
    assign G[36] = in1[20] & in2[20];
    assign P[36] = in1[20] ^ in2[20];
    assign G[37] = in1[19] & in2[19];
    assign P[37] = in1[19] ^ in2[19];
    assign G[38] = in1[18] & in2[18];
    assign P[38] = in1[18] ^ in2[18];
    assign G[39] = in1[17] & in2[17];
    assign P[39] = in1[17] ^ in2[17];
    assign G[40] = in1[16] & in2[16];
    assign P[40] = in1[16] ^ in2[16];
    assign G[41] = in1[15] & in2[15];
    assign P[41] = in1[15] ^ in2[15];
    assign G[42] = in1[14] & in2[14];
    assign P[42] = in1[14] ^ in2[14];
    assign G[43] = in1[13] & in2[13];
    assign P[43] = in1[13] ^ in2[13];
    assign G[44] = in1[12] & in2[12];
    assign P[44] = in1[12] ^ in2[12];
    assign G[45] = in1[11] & in2[11];
    assign P[45] = in1[11] ^ in2[11];
    assign G[46] = in1[10] & in2[10];
    assign P[46] = in1[10] ^ in2[10];
    assign G[47] = in1[9] & in2[9];
    assign P[47] = in1[9] ^ in2[9];
    assign G[48] = in1[8] & in2[8];
    assign P[48] = in1[8] ^ in2[8];
    assign G[49] = in1[7] & in2[7];
    assign P[49] = in1[7] ^ in2[7];
    assign G[50] = in1[6] & in2[6];
    assign P[50] = in1[6] ^ in2[6];
    assign G[51] = in1[5] & in2[5];
    assign P[51] = in1[5] ^ in2[5];
    assign G[52] = in1[4] & in2[4];
    assign P[52] = in1[4] ^ in2[4];
    assign G[53] = in1[3] & in2[3];
    assign P[53] = in1[3] ^ in2[3];
    assign G[54] = in1[2] & in2[2];
    assign P[54] = in1[2] ^ in2[2];
    assign G[55] = in1[1] & in2[1];
    assign P[55] = in1[1] ^ in2[1];
    assign G[56] = in1[0] & in2[0];
    assign P[56] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign cout = G[56] | (P[56] & C[56]);
    assign sum = P ^ C;
endmodule

module CLA_56(output [55:0] sum, output cout, input [55:0] in1, input [55:0] in2);

    wire[55:0] G;
    wire[55:0] C;
    wire[55:0] P;

    assign G[0] = in1[55] & in2[55];
    assign P[0] = in1[55] ^ in2[55];
    assign G[1] = in1[54] & in2[54];
    assign P[1] = in1[54] ^ in2[54];
    assign G[2] = in1[53] & in2[53];
    assign P[2] = in1[53] ^ in2[53];
    assign G[3] = in1[52] & in2[52];
    assign P[3] = in1[52] ^ in2[52];
    assign G[4] = in1[51] & in2[51];
    assign P[4] = in1[51] ^ in2[51];
    assign G[5] = in1[50] & in2[50];
    assign P[5] = in1[50] ^ in2[50];
    assign G[6] = in1[49] & in2[49];
    assign P[6] = in1[49] ^ in2[49];
    assign G[7] = in1[48] & in2[48];
    assign P[7] = in1[48] ^ in2[48];
    assign G[8] = in1[47] & in2[47];
    assign P[8] = in1[47] ^ in2[47];
    assign G[9] = in1[46] & in2[46];
    assign P[9] = in1[46] ^ in2[46];
    assign G[10] = in1[45] & in2[45];
    assign P[10] = in1[45] ^ in2[45];
    assign G[11] = in1[44] & in2[44];
    assign P[11] = in1[44] ^ in2[44];
    assign G[12] = in1[43] & in2[43];
    assign P[12] = in1[43] ^ in2[43];
    assign G[13] = in1[42] & in2[42];
    assign P[13] = in1[42] ^ in2[42];
    assign G[14] = in1[41] & in2[41];
    assign P[14] = in1[41] ^ in2[41];
    assign G[15] = in1[40] & in2[40];
    assign P[15] = in1[40] ^ in2[40];
    assign G[16] = in1[39] & in2[39];
    assign P[16] = in1[39] ^ in2[39];
    assign G[17] = in1[38] & in2[38];
    assign P[17] = in1[38] ^ in2[38];
    assign G[18] = in1[37] & in2[37];
    assign P[18] = in1[37] ^ in2[37];
    assign G[19] = in1[36] & in2[36];
    assign P[19] = in1[36] ^ in2[36];
    assign G[20] = in1[35] & in2[35];
    assign P[20] = in1[35] ^ in2[35];
    assign G[21] = in1[34] & in2[34];
    assign P[21] = in1[34] ^ in2[34];
    assign G[22] = in1[33] & in2[33];
    assign P[22] = in1[33] ^ in2[33];
    assign G[23] = in1[32] & in2[32];
    assign P[23] = in1[32] ^ in2[32];
    assign G[24] = in1[31] & in2[31];
    assign P[24] = in1[31] ^ in2[31];
    assign G[25] = in1[30] & in2[30];
    assign P[25] = in1[30] ^ in2[30];
    assign G[26] = in1[29] & in2[29];
    assign P[26] = in1[29] ^ in2[29];
    assign G[27] = in1[28] & in2[28];
    assign P[27] = in1[28] ^ in2[28];
    assign G[28] = in1[27] & in2[27];
    assign P[28] = in1[27] ^ in2[27];
    assign G[29] = in1[26] & in2[26];
    assign P[29] = in1[26] ^ in2[26];
    assign G[30] = in1[25] & in2[25];
    assign P[30] = in1[25] ^ in2[25];
    assign G[31] = in1[24] & in2[24];
    assign P[31] = in1[24] ^ in2[24];
    assign G[32] = in1[23] & in2[23];
    assign P[32] = in1[23] ^ in2[23];
    assign G[33] = in1[22] & in2[22];
    assign P[33] = in1[22] ^ in2[22];
    assign G[34] = in1[21] & in2[21];
    assign P[34] = in1[21] ^ in2[21];
    assign G[35] = in1[20] & in2[20];
    assign P[35] = in1[20] ^ in2[20];
    assign G[36] = in1[19] & in2[19];
    assign P[36] = in1[19] ^ in2[19];
    assign G[37] = in1[18] & in2[18];
    assign P[37] = in1[18] ^ in2[18];
    assign G[38] = in1[17] & in2[17];
    assign P[38] = in1[17] ^ in2[17];
    assign G[39] = in1[16] & in2[16];
    assign P[39] = in1[16] ^ in2[16];
    assign G[40] = in1[15] & in2[15];
    assign P[40] = in1[15] ^ in2[15];
    assign G[41] = in1[14] & in2[14];
    assign P[41] = in1[14] ^ in2[14];
    assign G[42] = in1[13] & in2[13];
    assign P[42] = in1[13] ^ in2[13];
    assign G[43] = in1[12] & in2[12];
    assign P[43] = in1[12] ^ in2[12];
    assign G[44] = in1[11] & in2[11];
    assign P[44] = in1[11] ^ in2[11];
    assign G[45] = in1[10] & in2[10];
    assign P[45] = in1[10] ^ in2[10];
    assign G[46] = in1[9] & in2[9];
    assign P[46] = in1[9] ^ in2[9];
    assign G[47] = in1[8] & in2[8];
    assign P[47] = in1[8] ^ in2[8];
    assign G[48] = in1[7] & in2[7];
    assign P[48] = in1[7] ^ in2[7];
    assign G[49] = in1[6] & in2[6];
    assign P[49] = in1[6] ^ in2[6];
    assign G[50] = in1[5] & in2[5];
    assign P[50] = in1[5] ^ in2[5];
    assign G[51] = in1[4] & in2[4];
    assign P[51] = in1[4] ^ in2[4];
    assign G[52] = in1[3] & in2[3];
    assign P[52] = in1[3] ^ in2[3];
    assign G[53] = in1[2] & in2[2];
    assign P[53] = in1[2] ^ in2[2];
    assign G[54] = in1[1] & in2[1];
    assign P[54] = in1[1] ^ in2[1];
    assign G[55] = in1[0] & in2[0];
    assign P[55] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign cout = G[55] | (P[55] & C[55]);
    assign sum = P ^ C;
endmodule

module CLA_55(output [54:0] sum, output cout, input [54:0] in1, input [54:0] in2);

    wire[54:0] G;
    wire[54:0] C;
    wire[54:0] P;

    assign G[0] = in1[54] & in2[54];
    assign P[0] = in1[54] ^ in2[54];
    assign G[1] = in1[53] & in2[53];
    assign P[1] = in1[53] ^ in2[53];
    assign G[2] = in1[52] & in2[52];
    assign P[2] = in1[52] ^ in2[52];
    assign G[3] = in1[51] & in2[51];
    assign P[3] = in1[51] ^ in2[51];
    assign G[4] = in1[50] & in2[50];
    assign P[4] = in1[50] ^ in2[50];
    assign G[5] = in1[49] & in2[49];
    assign P[5] = in1[49] ^ in2[49];
    assign G[6] = in1[48] & in2[48];
    assign P[6] = in1[48] ^ in2[48];
    assign G[7] = in1[47] & in2[47];
    assign P[7] = in1[47] ^ in2[47];
    assign G[8] = in1[46] & in2[46];
    assign P[8] = in1[46] ^ in2[46];
    assign G[9] = in1[45] & in2[45];
    assign P[9] = in1[45] ^ in2[45];
    assign G[10] = in1[44] & in2[44];
    assign P[10] = in1[44] ^ in2[44];
    assign G[11] = in1[43] & in2[43];
    assign P[11] = in1[43] ^ in2[43];
    assign G[12] = in1[42] & in2[42];
    assign P[12] = in1[42] ^ in2[42];
    assign G[13] = in1[41] & in2[41];
    assign P[13] = in1[41] ^ in2[41];
    assign G[14] = in1[40] & in2[40];
    assign P[14] = in1[40] ^ in2[40];
    assign G[15] = in1[39] & in2[39];
    assign P[15] = in1[39] ^ in2[39];
    assign G[16] = in1[38] & in2[38];
    assign P[16] = in1[38] ^ in2[38];
    assign G[17] = in1[37] & in2[37];
    assign P[17] = in1[37] ^ in2[37];
    assign G[18] = in1[36] & in2[36];
    assign P[18] = in1[36] ^ in2[36];
    assign G[19] = in1[35] & in2[35];
    assign P[19] = in1[35] ^ in2[35];
    assign G[20] = in1[34] & in2[34];
    assign P[20] = in1[34] ^ in2[34];
    assign G[21] = in1[33] & in2[33];
    assign P[21] = in1[33] ^ in2[33];
    assign G[22] = in1[32] & in2[32];
    assign P[22] = in1[32] ^ in2[32];
    assign G[23] = in1[31] & in2[31];
    assign P[23] = in1[31] ^ in2[31];
    assign G[24] = in1[30] & in2[30];
    assign P[24] = in1[30] ^ in2[30];
    assign G[25] = in1[29] & in2[29];
    assign P[25] = in1[29] ^ in2[29];
    assign G[26] = in1[28] & in2[28];
    assign P[26] = in1[28] ^ in2[28];
    assign G[27] = in1[27] & in2[27];
    assign P[27] = in1[27] ^ in2[27];
    assign G[28] = in1[26] & in2[26];
    assign P[28] = in1[26] ^ in2[26];
    assign G[29] = in1[25] & in2[25];
    assign P[29] = in1[25] ^ in2[25];
    assign G[30] = in1[24] & in2[24];
    assign P[30] = in1[24] ^ in2[24];
    assign G[31] = in1[23] & in2[23];
    assign P[31] = in1[23] ^ in2[23];
    assign G[32] = in1[22] & in2[22];
    assign P[32] = in1[22] ^ in2[22];
    assign G[33] = in1[21] & in2[21];
    assign P[33] = in1[21] ^ in2[21];
    assign G[34] = in1[20] & in2[20];
    assign P[34] = in1[20] ^ in2[20];
    assign G[35] = in1[19] & in2[19];
    assign P[35] = in1[19] ^ in2[19];
    assign G[36] = in1[18] & in2[18];
    assign P[36] = in1[18] ^ in2[18];
    assign G[37] = in1[17] & in2[17];
    assign P[37] = in1[17] ^ in2[17];
    assign G[38] = in1[16] & in2[16];
    assign P[38] = in1[16] ^ in2[16];
    assign G[39] = in1[15] & in2[15];
    assign P[39] = in1[15] ^ in2[15];
    assign G[40] = in1[14] & in2[14];
    assign P[40] = in1[14] ^ in2[14];
    assign G[41] = in1[13] & in2[13];
    assign P[41] = in1[13] ^ in2[13];
    assign G[42] = in1[12] & in2[12];
    assign P[42] = in1[12] ^ in2[12];
    assign G[43] = in1[11] & in2[11];
    assign P[43] = in1[11] ^ in2[11];
    assign G[44] = in1[10] & in2[10];
    assign P[44] = in1[10] ^ in2[10];
    assign G[45] = in1[9] & in2[9];
    assign P[45] = in1[9] ^ in2[9];
    assign G[46] = in1[8] & in2[8];
    assign P[46] = in1[8] ^ in2[8];
    assign G[47] = in1[7] & in2[7];
    assign P[47] = in1[7] ^ in2[7];
    assign G[48] = in1[6] & in2[6];
    assign P[48] = in1[6] ^ in2[6];
    assign G[49] = in1[5] & in2[5];
    assign P[49] = in1[5] ^ in2[5];
    assign G[50] = in1[4] & in2[4];
    assign P[50] = in1[4] ^ in2[4];
    assign G[51] = in1[3] & in2[3];
    assign P[51] = in1[3] ^ in2[3];
    assign G[52] = in1[2] & in2[2];
    assign P[52] = in1[2] ^ in2[2];
    assign G[53] = in1[1] & in2[1];
    assign P[53] = in1[1] ^ in2[1];
    assign G[54] = in1[0] & in2[0];
    assign P[54] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign cout = G[54] | (P[54] & C[54]);
    assign sum = P ^ C;
endmodule

module CLA_54(output [53:0] sum, output cout, input [53:0] in1, input [53:0] in2);

    wire[53:0] G;
    wire[53:0] C;
    wire[53:0] P;

    assign G[0] = in1[53] & in2[53];
    assign P[0] = in1[53] ^ in2[53];
    assign G[1] = in1[52] & in2[52];
    assign P[1] = in1[52] ^ in2[52];
    assign G[2] = in1[51] & in2[51];
    assign P[2] = in1[51] ^ in2[51];
    assign G[3] = in1[50] & in2[50];
    assign P[3] = in1[50] ^ in2[50];
    assign G[4] = in1[49] & in2[49];
    assign P[4] = in1[49] ^ in2[49];
    assign G[5] = in1[48] & in2[48];
    assign P[5] = in1[48] ^ in2[48];
    assign G[6] = in1[47] & in2[47];
    assign P[6] = in1[47] ^ in2[47];
    assign G[7] = in1[46] & in2[46];
    assign P[7] = in1[46] ^ in2[46];
    assign G[8] = in1[45] & in2[45];
    assign P[8] = in1[45] ^ in2[45];
    assign G[9] = in1[44] & in2[44];
    assign P[9] = in1[44] ^ in2[44];
    assign G[10] = in1[43] & in2[43];
    assign P[10] = in1[43] ^ in2[43];
    assign G[11] = in1[42] & in2[42];
    assign P[11] = in1[42] ^ in2[42];
    assign G[12] = in1[41] & in2[41];
    assign P[12] = in1[41] ^ in2[41];
    assign G[13] = in1[40] & in2[40];
    assign P[13] = in1[40] ^ in2[40];
    assign G[14] = in1[39] & in2[39];
    assign P[14] = in1[39] ^ in2[39];
    assign G[15] = in1[38] & in2[38];
    assign P[15] = in1[38] ^ in2[38];
    assign G[16] = in1[37] & in2[37];
    assign P[16] = in1[37] ^ in2[37];
    assign G[17] = in1[36] & in2[36];
    assign P[17] = in1[36] ^ in2[36];
    assign G[18] = in1[35] & in2[35];
    assign P[18] = in1[35] ^ in2[35];
    assign G[19] = in1[34] & in2[34];
    assign P[19] = in1[34] ^ in2[34];
    assign G[20] = in1[33] & in2[33];
    assign P[20] = in1[33] ^ in2[33];
    assign G[21] = in1[32] & in2[32];
    assign P[21] = in1[32] ^ in2[32];
    assign G[22] = in1[31] & in2[31];
    assign P[22] = in1[31] ^ in2[31];
    assign G[23] = in1[30] & in2[30];
    assign P[23] = in1[30] ^ in2[30];
    assign G[24] = in1[29] & in2[29];
    assign P[24] = in1[29] ^ in2[29];
    assign G[25] = in1[28] & in2[28];
    assign P[25] = in1[28] ^ in2[28];
    assign G[26] = in1[27] & in2[27];
    assign P[26] = in1[27] ^ in2[27];
    assign G[27] = in1[26] & in2[26];
    assign P[27] = in1[26] ^ in2[26];
    assign G[28] = in1[25] & in2[25];
    assign P[28] = in1[25] ^ in2[25];
    assign G[29] = in1[24] & in2[24];
    assign P[29] = in1[24] ^ in2[24];
    assign G[30] = in1[23] & in2[23];
    assign P[30] = in1[23] ^ in2[23];
    assign G[31] = in1[22] & in2[22];
    assign P[31] = in1[22] ^ in2[22];
    assign G[32] = in1[21] & in2[21];
    assign P[32] = in1[21] ^ in2[21];
    assign G[33] = in1[20] & in2[20];
    assign P[33] = in1[20] ^ in2[20];
    assign G[34] = in1[19] & in2[19];
    assign P[34] = in1[19] ^ in2[19];
    assign G[35] = in1[18] & in2[18];
    assign P[35] = in1[18] ^ in2[18];
    assign G[36] = in1[17] & in2[17];
    assign P[36] = in1[17] ^ in2[17];
    assign G[37] = in1[16] & in2[16];
    assign P[37] = in1[16] ^ in2[16];
    assign G[38] = in1[15] & in2[15];
    assign P[38] = in1[15] ^ in2[15];
    assign G[39] = in1[14] & in2[14];
    assign P[39] = in1[14] ^ in2[14];
    assign G[40] = in1[13] & in2[13];
    assign P[40] = in1[13] ^ in2[13];
    assign G[41] = in1[12] & in2[12];
    assign P[41] = in1[12] ^ in2[12];
    assign G[42] = in1[11] & in2[11];
    assign P[42] = in1[11] ^ in2[11];
    assign G[43] = in1[10] & in2[10];
    assign P[43] = in1[10] ^ in2[10];
    assign G[44] = in1[9] & in2[9];
    assign P[44] = in1[9] ^ in2[9];
    assign G[45] = in1[8] & in2[8];
    assign P[45] = in1[8] ^ in2[8];
    assign G[46] = in1[7] & in2[7];
    assign P[46] = in1[7] ^ in2[7];
    assign G[47] = in1[6] & in2[6];
    assign P[47] = in1[6] ^ in2[6];
    assign G[48] = in1[5] & in2[5];
    assign P[48] = in1[5] ^ in2[5];
    assign G[49] = in1[4] & in2[4];
    assign P[49] = in1[4] ^ in2[4];
    assign G[50] = in1[3] & in2[3];
    assign P[50] = in1[3] ^ in2[3];
    assign G[51] = in1[2] & in2[2];
    assign P[51] = in1[2] ^ in2[2];
    assign G[52] = in1[1] & in2[1];
    assign P[52] = in1[1] ^ in2[1];
    assign G[53] = in1[0] & in2[0];
    assign P[53] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign cout = G[53] | (P[53] & C[53]);
    assign sum = P ^ C;
endmodule

module CLA_53(output [52:0] sum, output cout, input [52:0] in1, input [52:0] in2);

    wire[52:0] G;
    wire[52:0] C;
    wire[52:0] P;

    assign G[0] = in1[52] & in2[52];
    assign P[0] = in1[52] ^ in2[52];
    assign G[1] = in1[51] & in2[51];
    assign P[1] = in1[51] ^ in2[51];
    assign G[2] = in1[50] & in2[50];
    assign P[2] = in1[50] ^ in2[50];
    assign G[3] = in1[49] & in2[49];
    assign P[3] = in1[49] ^ in2[49];
    assign G[4] = in1[48] & in2[48];
    assign P[4] = in1[48] ^ in2[48];
    assign G[5] = in1[47] & in2[47];
    assign P[5] = in1[47] ^ in2[47];
    assign G[6] = in1[46] & in2[46];
    assign P[6] = in1[46] ^ in2[46];
    assign G[7] = in1[45] & in2[45];
    assign P[7] = in1[45] ^ in2[45];
    assign G[8] = in1[44] & in2[44];
    assign P[8] = in1[44] ^ in2[44];
    assign G[9] = in1[43] & in2[43];
    assign P[9] = in1[43] ^ in2[43];
    assign G[10] = in1[42] & in2[42];
    assign P[10] = in1[42] ^ in2[42];
    assign G[11] = in1[41] & in2[41];
    assign P[11] = in1[41] ^ in2[41];
    assign G[12] = in1[40] & in2[40];
    assign P[12] = in1[40] ^ in2[40];
    assign G[13] = in1[39] & in2[39];
    assign P[13] = in1[39] ^ in2[39];
    assign G[14] = in1[38] & in2[38];
    assign P[14] = in1[38] ^ in2[38];
    assign G[15] = in1[37] & in2[37];
    assign P[15] = in1[37] ^ in2[37];
    assign G[16] = in1[36] & in2[36];
    assign P[16] = in1[36] ^ in2[36];
    assign G[17] = in1[35] & in2[35];
    assign P[17] = in1[35] ^ in2[35];
    assign G[18] = in1[34] & in2[34];
    assign P[18] = in1[34] ^ in2[34];
    assign G[19] = in1[33] & in2[33];
    assign P[19] = in1[33] ^ in2[33];
    assign G[20] = in1[32] & in2[32];
    assign P[20] = in1[32] ^ in2[32];
    assign G[21] = in1[31] & in2[31];
    assign P[21] = in1[31] ^ in2[31];
    assign G[22] = in1[30] & in2[30];
    assign P[22] = in1[30] ^ in2[30];
    assign G[23] = in1[29] & in2[29];
    assign P[23] = in1[29] ^ in2[29];
    assign G[24] = in1[28] & in2[28];
    assign P[24] = in1[28] ^ in2[28];
    assign G[25] = in1[27] & in2[27];
    assign P[25] = in1[27] ^ in2[27];
    assign G[26] = in1[26] & in2[26];
    assign P[26] = in1[26] ^ in2[26];
    assign G[27] = in1[25] & in2[25];
    assign P[27] = in1[25] ^ in2[25];
    assign G[28] = in1[24] & in2[24];
    assign P[28] = in1[24] ^ in2[24];
    assign G[29] = in1[23] & in2[23];
    assign P[29] = in1[23] ^ in2[23];
    assign G[30] = in1[22] & in2[22];
    assign P[30] = in1[22] ^ in2[22];
    assign G[31] = in1[21] & in2[21];
    assign P[31] = in1[21] ^ in2[21];
    assign G[32] = in1[20] & in2[20];
    assign P[32] = in1[20] ^ in2[20];
    assign G[33] = in1[19] & in2[19];
    assign P[33] = in1[19] ^ in2[19];
    assign G[34] = in1[18] & in2[18];
    assign P[34] = in1[18] ^ in2[18];
    assign G[35] = in1[17] & in2[17];
    assign P[35] = in1[17] ^ in2[17];
    assign G[36] = in1[16] & in2[16];
    assign P[36] = in1[16] ^ in2[16];
    assign G[37] = in1[15] & in2[15];
    assign P[37] = in1[15] ^ in2[15];
    assign G[38] = in1[14] & in2[14];
    assign P[38] = in1[14] ^ in2[14];
    assign G[39] = in1[13] & in2[13];
    assign P[39] = in1[13] ^ in2[13];
    assign G[40] = in1[12] & in2[12];
    assign P[40] = in1[12] ^ in2[12];
    assign G[41] = in1[11] & in2[11];
    assign P[41] = in1[11] ^ in2[11];
    assign G[42] = in1[10] & in2[10];
    assign P[42] = in1[10] ^ in2[10];
    assign G[43] = in1[9] & in2[9];
    assign P[43] = in1[9] ^ in2[9];
    assign G[44] = in1[8] & in2[8];
    assign P[44] = in1[8] ^ in2[8];
    assign G[45] = in1[7] & in2[7];
    assign P[45] = in1[7] ^ in2[7];
    assign G[46] = in1[6] & in2[6];
    assign P[46] = in1[6] ^ in2[6];
    assign G[47] = in1[5] & in2[5];
    assign P[47] = in1[5] ^ in2[5];
    assign G[48] = in1[4] & in2[4];
    assign P[48] = in1[4] ^ in2[4];
    assign G[49] = in1[3] & in2[3];
    assign P[49] = in1[3] ^ in2[3];
    assign G[50] = in1[2] & in2[2];
    assign P[50] = in1[2] ^ in2[2];
    assign G[51] = in1[1] & in2[1];
    assign P[51] = in1[1] ^ in2[1];
    assign G[52] = in1[0] & in2[0];
    assign P[52] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign cout = G[52] | (P[52] & C[52]);
    assign sum = P ^ C;
endmodule

module CLA_52(output [51:0] sum, output cout, input [51:0] in1, input [51:0] in2);

    wire[51:0] G;
    wire[51:0] C;
    wire[51:0] P;

    assign G[0] = in1[51] & in2[51];
    assign P[0] = in1[51] ^ in2[51];
    assign G[1] = in1[50] & in2[50];
    assign P[1] = in1[50] ^ in2[50];
    assign G[2] = in1[49] & in2[49];
    assign P[2] = in1[49] ^ in2[49];
    assign G[3] = in1[48] & in2[48];
    assign P[3] = in1[48] ^ in2[48];
    assign G[4] = in1[47] & in2[47];
    assign P[4] = in1[47] ^ in2[47];
    assign G[5] = in1[46] & in2[46];
    assign P[5] = in1[46] ^ in2[46];
    assign G[6] = in1[45] & in2[45];
    assign P[6] = in1[45] ^ in2[45];
    assign G[7] = in1[44] & in2[44];
    assign P[7] = in1[44] ^ in2[44];
    assign G[8] = in1[43] & in2[43];
    assign P[8] = in1[43] ^ in2[43];
    assign G[9] = in1[42] & in2[42];
    assign P[9] = in1[42] ^ in2[42];
    assign G[10] = in1[41] & in2[41];
    assign P[10] = in1[41] ^ in2[41];
    assign G[11] = in1[40] & in2[40];
    assign P[11] = in1[40] ^ in2[40];
    assign G[12] = in1[39] & in2[39];
    assign P[12] = in1[39] ^ in2[39];
    assign G[13] = in1[38] & in2[38];
    assign P[13] = in1[38] ^ in2[38];
    assign G[14] = in1[37] & in2[37];
    assign P[14] = in1[37] ^ in2[37];
    assign G[15] = in1[36] & in2[36];
    assign P[15] = in1[36] ^ in2[36];
    assign G[16] = in1[35] & in2[35];
    assign P[16] = in1[35] ^ in2[35];
    assign G[17] = in1[34] & in2[34];
    assign P[17] = in1[34] ^ in2[34];
    assign G[18] = in1[33] & in2[33];
    assign P[18] = in1[33] ^ in2[33];
    assign G[19] = in1[32] & in2[32];
    assign P[19] = in1[32] ^ in2[32];
    assign G[20] = in1[31] & in2[31];
    assign P[20] = in1[31] ^ in2[31];
    assign G[21] = in1[30] & in2[30];
    assign P[21] = in1[30] ^ in2[30];
    assign G[22] = in1[29] & in2[29];
    assign P[22] = in1[29] ^ in2[29];
    assign G[23] = in1[28] & in2[28];
    assign P[23] = in1[28] ^ in2[28];
    assign G[24] = in1[27] & in2[27];
    assign P[24] = in1[27] ^ in2[27];
    assign G[25] = in1[26] & in2[26];
    assign P[25] = in1[26] ^ in2[26];
    assign G[26] = in1[25] & in2[25];
    assign P[26] = in1[25] ^ in2[25];
    assign G[27] = in1[24] & in2[24];
    assign P[27] = in1[24] ^ in2[24];
    assign G[28] = in1[23] & in2[23];
    assign P[28] = in1[23] ^ in2[23];
    assign G[29] = in1[22] & in2[22];
    assign P[29] = in1[22] ^ in2[22];
    assign G[30] = in1[21] & in2[21];
    assign P[30] = in1[21] ^ in2[21];
    assign G[31] = in1[20] & in2[20];
    assign P[31] = in1[20] ^ in2[20];
    assign G[32] = in1[19] & in2[19];
    assign P[32] = in1[19] ^ in2[19];
    assign G[33] = in1[18] & in2[18];
    assign P[33] = in1[18] ^ in2[18];
    assign G[34] = in1[17] & in2[17];
    assign P[34] = in1[17] ^ in2[17];
    assign G[35] = in1[16] & in2[16];
    assign P[35] = in1[16] ^ in2[16];
    assign G[36] = in1[15] & in2[15];
    assign P[36] = in1[15] ^ in2[15];
    assign G[37] = in1[14] & in2[14];
    assign P[37] = in1[14] ^ in2[14];
    assign G[38] = in1[13] & in2[13];
    assign P[38] = in1[13] ^ in2[13];
    assign G[39] = in1[12] & in2[12];
    assign P[39] = in1[12] ^ in2[12];
    assign G[40] = in1[11] & in2[11];
    assign P[40] = in1[11] ^ in2[11];
    assign G[41] = in1[10] & in2[10];
    assign P[41] = in1[10] ^ in2[10];
    assign G[42] = in1[9] & in2[9];
    assign P[42] = in1[9] ^ in2[9];
    assign G[43] = in1[8] & in2[8];
    assign P[43] = in1[8] ^ in2[8];
    assign G[44] = in1[7] & in2[7];
    assign P[44] = in1[7] ^ in2[7];
    assign G[45] = in1[6] & in2[6];
    assign P[45] = in1[6] ^ in2[6];
    assign G[46] = in1[5] & in2[5];
    assign P[46] = in1[5] ^ in2[5];
    assign G[47] = in1[4] & in2[4];
    assign P[47] = in1[4] ^ in2[4];
    assign G[48] = in1[3] & in2[3];
    assign P[48] = in1[3] ^ in2[3];
    assign G[49] = in1[2] & in2[2];
    assign P[49] = in1[2] ^ in2[2];
    assign G[50] = in1[1] & in2[1];
    assign P[50] = in1[1] ^ in2[1];
    assign G[51] = in1[0] & in2[0];
    assign P[51] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign cout = G[51] | (P[51] & C[51]);
    assign sum = P ^ C;
endmodule

module CLA_51(output [50:0] sum, output cout, input [50:0] in1, input [50:0] in2);

    wire[50:0] G;
    wire[50:0] C;
    wire[50:0] P;

    assign G[0] = in1[50] & in2[50];
    assign P[0] = in1[50] ^ in2[50];
    assign G[1] = in1[49] & in2[49];
    assign P[1] = in1[49] ^ in2[49];
    assign G[2] = in1[48] & in2[48];
    assign P[2] = in1[48] ^ in2[48];
    assign G[3] = in1[47] & in2[47];
    assign P[3] = in1[47] ^ in2[47];
    assign G[4] = in1[46] & in2[46];
    assign P[4] = in1[46] ^ in2[46];
    assign G[5] = in1[45] & in2[45];
    assign P[5] = in1[45] ^ in2[45];
    assign G[6] = in1[44] & in2[44];
    assign P[6] = in1[44] ^ in2[44];
    assign G[7] = in1[43] & in2[43];
    assign P[7] = in1[43] ^ in2[43];
    assign G[8] = in1[42] & in2[42];
    assign P[8] = in1[42] ^ in2[42];
    assign G[9] = in1[41] & in2[41];
    assign P[9] = in1[41] ^ in2[41];
    assign G[10] = in1[40] & in2[40];
    assign P[10] = in1[40] ^ in2[40];
    assign G[11] = in1[39] & in2[39];
    assign P[11] = in1[39] ^ in2[39];
    assign G[12] = in1[38] & in2[38];
    assign P[12] = in1[38] ^ in2[38];
    assign G[13] = in1[37] & in2[37];
    assign P[13] = in1[37] ^ in2[37];
    assign G[14] = in1[36] & in2[36];
    assign P[14] = in1[36] ^ in2[36];
    assign G[15] = in1[35] & in2[35];
    assign P[15] = in1[35] ^ in2[35];
    assign G[16] = in1[34] & in2[34];
    assign P[16] = in1[34] ^ in2[34];
    assign G[17] = in1[33] & in2[33];
    assign P[17] = in1[33] ^ in2[33];
    assign G[18] = in1[32] & in2[32];
    assign P[18] = in1[32] ^ in2[32];
    assign G[19] = in1[31] & in2[31];
    assign P[19] = in1[31] ^ in2[31];
    assign G[20] = in1[30] & in2[30];
    assign P[20] = in1[30] ^ in2[30];
    assign G[21] = in1[29] & in2[29];
    assign P[21] = in1[29] ^ in2[29];
    assign G[22] = in1[28] & in2[28];
    assign P[22] = in1[28] ^ in2[28];
    assign G[23] = in1[27] & in2[27];
    assign P[23] = in1[27] ^ in2[27];
    assign G[24] = in1[26] & in2[26];
    assign P[24] = in1[26] ^ in2[26];
    assign G[25] = in1[25] & in2[25];
    assign P[25] = in1[25] ^ in2[25];
    assign G[26] = in1[24] & in2[24];
    assign P[26] = in1[24] ^ in2[24];
    assign G[27] = in1[23] & in2[23];
    assign P[27] = in1[23] ^ in2[23];
    assign G[28] = in1[22] & in2[22];
    assign P[28] = in1[22] ^ in2[22];
    assign G[29] = in1[21] & in2[21];
    assign P[29] = in1[21] ^ in2[21];
    assign G[30] = in1[20] & in2[20];
    assign P[30] = in1[20] ^ in2[20];
    assign G[31] = in1[19] & in2[19];
    assign P[31] = in1[19] ^ in2[19];
    assign G[32] = in1[18] & in2[18];
    assign P[32] = in1[18] ^ in2[18];
    assign G[33] = in1[17] & in2[17];
    assign P[33] = in1[17] ^ in2[17];
    assign G[34] = in1[16] & in2[16];
    assign P[34] = in1[16] ^ in2[16];
    assign G[35] = in1[15] & in2[15];
    assign P[35] = in1[15] ^ in2[15];
    assign G[36] = in1[14] & in2[14];
    assign P[36] = in1[14] ^ in2[14];
    assign G[37] = in1[13] & in2[13];
    assign P[37] = in1[13] ^ in2[13];
    assign G[38] = in1[12] & in2[12];
    assign P[38] = in1[12] ^ in2[12];
    assign G[39] = in1[11] & in2[11];
    assign P[39] = in1[11] ^ in2[11];
    assign G[40] = in1[10] & in2[10];
    assign P[40] = in1[10] ^ in2[10];
    assign G[41] = in1[9] & in2[9];
    assign P[41] = in1[9] ^ in2[9];
    assign G[42] = in1[8] & in2[8];
    assign P[42] = in1[8] ^ in2[8];
    assign G[43] = in1[7] & in2[7];
    assign P[43] = in1[7] ^ in2[7];
    assign G[44] = in1[6] & in2[6];
    assign P[44] = in1[6] ^ in2[6];
    assign G[45] = in1[5] & in2[5];
    assign P[45] = in1[5] ^ in2[5];
    assign G[46] = in1[4] & in2[4];
    assign P[46] = in1[4] ^ in2[4];
    assign G[47] = in1[3] & in2[3];
    assign P[47] = in1[3] ^ in2[3];
    assign G[48] = in1[2] & in2[2];
    assign P[48] = in1[2] ^ in2[2];
    assign G[49] = in1[1] & in2[1];
    assign P[49] = in1[1] ^ in2[1];
    assign G[50] = in1[0] & in2[0];
    assign P[50] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign cout = G[50] | (P[50] & C[50]);
    assign sum = P ^ C;
endmodule

module CLA_50(output [49:0] sum, output cout, input [49:0] in1, input [49:0] in2);

    wire[49:0] G;
    wire[49:0] C;
    wire[49:0] P;

    assign G[0] = in1[49] & in2[49];
    assign P[0] = in1[49] ^ in2[49];
    assign G[1] = in1[48] & in2[48];
    assign P[1] = in1[48] ^ in2[48];
    assign G[2] = in1[47] & in2[47];
    assign P[2] = in1[47] ^ in2[47];
    assign G[3] = in1[46] & in2[46];
    assign P[3] = in1[46] ^ in2[46];
    assign G[4] = in1[45] & in2[45];
    assign P[4] = in1[45] ^ in2[45];
    assign G[5] = in1[44] & in2[44];
    assign P[5] = in1[44] ^ in2[44];
    assign G[6] = in1[43] & in2[43];
    assign P[6] = in1[43] ^ in2[43];
    assign G[7] = in1[42] & in2[42];
    assign P[7] = in1[42] ^ in2[42];
    assign G[8] = in1[41] & in2[41];
    assign P[8] = in1[41] ^ in2[41];
    assign G[9] = in1[40] & in2[40];
    assign P[9] = in1[40] ^ in2[40];
    assign G[10] = in1[39] & in2[39];
    assign P[10] = in1[39] ^ in2[39];
    assign G[11] = in1[38] & in2[38];
    assign P[11] = in1[38] ^ in2[38];
    assign G[12] = in1[37] & in2[37];
    assign P[12] = in1[37] ^ in2[37];
    assign G[13] = in1[36] & in2[36];
    assign P[13] = in1[36] ^ in2[36];
    assign G[14] = in1[35] & in2[35];
    assign P[14] = in1[35] ^ in2[35];
    assign G[15] = in1[34] & in2[34];
    assign P[15] = in1[34] ^ in2[34];
    assign G[16] = in1[33] & in2[33];
    assign P[16] = in1[33] ^ in2[33];
    assign G[17] = in1[32] & in2[32];
    assign P[17] = in1[32] ^ in2[32];
    assign G[18] = in1[31] & in2[31];
    assign P[18] = in1[31] ^ in2[31];
    assign G[19] = in1[30] & in2[30];
    assign P[19] = in1[30] ^ in2[30];
    assign G[20] = in1[29] & in2[29];
    assign P[20] = in1[29] ^ in2[29];
    assign G[21] = in1[28] & in2[28];
    assign P[21] = in1[28] ^ in2[28];
    assign G[22] = in1[27] & in2[27];
    assign P[22] = in1[27] ^ in2[27];
    assign G[23] = in1[26] & in2[26];
    assign P[23] = in1[26] ^ in2[26];
    assign G[24] = in1[25] & in2[25];
    assign P[24] = in1[25] ^ in2[25];
    assign G[25] = in1[24] & in2[24];
    assign P[25] = in1[24] ^ in2[24];
    assign G[26] = in1[23] & in2[23];
    assign P[26] = in1[23] ^ in2[23];
    assign G[27] = in1[22] & in2[22];
    assign P[27] = in1[22] ^ in2[22];
    assign G[28] = in1[21] & in2[21];
    assign P[28] = in1[21] ^ in2[21];
    assign G[29] = in1[20] & in2[20];
    assign P[29] = in1[20] ^ in2[20];
    assign G[30] = in1[19] & in2[19];
    assign P[30] = in1[19] ^ in2[19];
    assign G[31] = in1[18] & in2[18];
    assign P[31] = in1[18] ^ in2[18];
    assign G[32] = in1[17] & in2[17];
    assign P[32] = in1[17] ^ in2[17];
    assign G[33] = in1[16] & in2[16];
    assign P[33] = in1[16] ^ in2[16];
    assign G[34] = in1[15] & in2[15];
    assign P[34] = in1[15] ^ in2[15];
    assign G[35] = in1[14] & in2[14];
    assign P[35] = in1[14] ^ in2[14];
    assign G[36] = in1[13] & in2[13];
    assign P[36] = in1[13] ^ in2[13];
    assign G[37] = in1[12] & in2[12];
    assign P[37] = in1[12] ^ in2[12];
    assign G[38] = in1[11] & in2[11];
    assign P[38] = in1[11] ^ in2[11];
    assign G[39] = in1[10] & in2[10];
    assign P[39] = in1[10] ^ in2[10];
    assign G[40] = in1[9] & in2[9];
    assign P[40] = in1[9] ^ in2[9];
    assign G[41] = in1[8] & in2[8];
    assign P[41] = in1[8] ^ in2[8];
    assign G[42] = in1[7] & in2[7];
    assign P[42] = in1[7] ^ in2[7];
    assign G[43] = in1[6] & in2[6];
    assign P[43] = in1[6] ^ in2[6];
    assign G[44] = in1[5] & in2[5];
    assign P[44] = in1[5] ^ in2[5];
    assign G[45] = in1[4] & in2[4];
    assign P[45] = in1[4] ^ in2[4];
    assign G[46] = in1[3] & in2[3];
    assign P[46] = in1[3] ^ in2[3];
    assign G[47] = in1[2] & in2[2];
    assign P[47] = in1[2] ^ in2[2];
    assign G[48] = in1[1] & in2[1];
    assign P[48] = in1[1] ^ in2[1];
    assign G[49] = in1[0] & in2[0];
    assign P[49] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign cout = G[49] | (P[49] & C[49]);
    assign sum = P ^ C;
endmodule

module CLA_49(output [48:0] sum, output cout, input [48:0] in1, input [48:0] in2);

    wire[48:0] G;
    wire[48:0] C;
    wire[48:0] P;

    assign G[0] = in1[48] & in2[48];
    assign P[0] = in1[48] ^ in2[48];
    assign G[1] = in1[47] & in2[47];
    assign P[1] = in1[47] ^ in2[47];
    assign G[2] = in1[46] & in2[46];
    assign P[2] = in1[46] ^ in2[46];
    assign G[3] = in1[45] & in2[45];
    assign P[3] = in1[45] ^ in2[45];
    assign G[4] = in1[44] & in2[44];
    assign P[4] = in1[44] ^ in2[44];
    assign G[5] = in1[43] & in2[43];
    assign P[5] = in1[43] ^ in2[43];
    assign G[6] = in1[42] & in2[42];
    assign P[6] = in1[42] ^ in2[42];
    assign G[7] = in1[41] & in2[41];
    assign P[7] = in1[41] ^ in2[41];
    assign G[8] = in1[40] & in2[40];
    assign P[8] = in1[40] ^ in2[40];
    assign G[9] = in1[39] & in2[39];
    assign P[9] = in1[39] ^ in2[39];
    assign G[10] = in1[38] & in2[38];
    assign P[10] = in1[38] ^ in2[38];
    assign G[11] = in1[37] & in2[37];
    assign P[11] = in1[37] ^ in2[37];
    assign G[12] = in1[36] & in2[36];
    assign P[12] = in1[36] ^ in2[36];
    assign G[13] = in1[35] & in2[35];
    assign P[13] = in1[35] ^ in2[35];
    assign G[14] = in1[34] & in2[34];
    assign P[14] = in1[34] ^ in2[34];
    assign G[15] = in1[33] & in2[33];
    assign P[15] = in1[33] ^ in2[33];
    assign G[16] = in1[32] & in2[32];
    assign P[16] = in1[32] ^ in2[32];
    assign G[17] = in1[31] & in2[31];
    assign P[17] = in1[31] ^ in2[31];
    assign G[18] = in1[30] & in2[30];
    assign P[18] = in1[30] ^ in2[30];
    assign G[19] = in1[29] & in2[29];
    assign P[19] = in1[29] ^ in2[29];
    assign G[20] = in1[28] & in2[28];
    assign P[20] = in1[28] ^ in2[28];
    assign G[21] = in1[27] & in2[27];
    assign P[21] = in1[27] ^ in2[27];
    assign G[22] = in1[26] & in2[26];
    assign P[22] = in1[26] ^ in2[26];
    assign G[23] = in1[25] & in2[25];
    assign P[23] = in1[25] ^ in2[25];
    assign G[24] = in1[24] & in2[24];
    assign P[24] = in1[24] ^ in2[24];
    assign G[25] = in1[23] & in2[23];
    assign P[25] = in1[23] ^ in2[23];
    assign G[26] = in1[22] & in2[22];
    assign P[26] = in1[22] ^ in2[22];
    assign G[27] = in1[21] & in2[21];
    assign P[27] = in1[21] ^ in2[21];
    assign G[28] = in1[20] & in2[20];
    assign P[28] = in1[20] ^ in2[20];
    assign G[29] = in1[19] & in2[19];
    assign P[29] = in1[19] ^ in2[19];
    assign G[30] = in1[18] & in2[18];
    assign P[30] = in1[18] ^ in2[18];
    assign G[31] = in1[17] & in2[17];
    assign P[31] = in1[17] ^ in2[17];
    assign G[32] = in1[16] & in2[16];
    assign P[32] = in1[16] ^ in2[16];
    assign G[33] = in1[15] & in2[15];
    assign P[33] = in1[15] ^ in2[15];
    assign G[34] = in1[14] & in2[14];
    assign P[34] = in1[14] ^ in2[14];
    assign G[35] = in1[13] & in2[13];
    assign P[35] = in1[13] ^ in2[13];
    assign G[36] = in1[12] & in2[12];
    assign P[36] = in1[12] ^ in2[12];
    assign G[37] = in1[11] & in2[11];
    assign P[37] = in1[11] ^ in2[11];
    assign G[38] = in1[10] & in2[10];
    assign P[38] = in1[10] ^ in2[10];
    assign G[39] = in1[9] & in2[9];
    assign P[39] = in1[9] ^ in2[9];
    assign G[40] = in1[8] & in2[8];
    assign P[40] = in1[8] ^ in2[8];
    assign G[41] = in1[7] & in2[7];
    assign P[41] = in1[7] ^ in2[7];
    assign G[42] = in1[6] & in2[6];
    assign P[42] = in1[6] ^ in2[6];
    assign G[43] = in1[5] & in2[5];
    assign P[43] = in1[5] ^ in2[5];
    assign G[44] = in1[4] & in2[4];
    assign P[44] = in1[4] ^ in2[4];
    assign G[45] = in1[3] & in2[3];
    assign P[45] = in1[3] ^ in2[3];
    assign G[46] = in1[2] & in2[2];
    assign P[46] = in1[2] ^ in2[2];
    assign G[47] = in1[1] & in2[1];
    assign P[47] = in1[1] ^ in2[1];
    assign G[48] = in1[0] & in2[0];
    assign P[48] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign cout = G[48] | (P[48] & C[48]);
    assign sum = P ^ C;
endmodule

module CLA_48(output [47:0] sum, output cout, input [47:0] in1, input [47:0] in2);

    wire[47:0] G;
    wire[47:0] C;
    wire[47:0] P;

    assign G[0] = in1[47] & in2[47];
    assign P[0] = in1[47] ^ in2[47];
    assign G[1] = in1[46] & in2[46];
    assign P[1] = in1[46] ^ in2[46];
    assign G[2] = in1[45] & in2[45];
    assign P[2] = in1[45] ^ in2[45];
    assign G[3] = in1[44] & in2[44];
    assign P[3] = in1[44] ^ in2[44];
    assign G[4] = in1[43] & in2[43];
    assign P[4] = in1[43] ^ in2[43];
    assign G[5] = in1[42] & in2[42];
    assign P[5] = in1[42] ^ in2[42];
    assign G[6] = in1[41] & in2[41];
    assign P[6] = in1[41] ^ in2[41];
    assign G[7] = in1[40] & in2[40];
    assign P[7] = in1[40] ^ in2[40];
    assign G[8] = in1[39] & in2[39];
    assign P[8] = in1[39] ^ in2[39];
    assign G[9] = in1[38] & in2[38];
    assign P[9] = in1[38] ^ in2[38];
    assign G[10] = in1[37] & in2[37];
    assign P[10] = in1[37] ^ in2[37];
    assign G[11] = in1[36] & in2[36];
    assign P[11] = in1[36] ^ in2[36];
    assign G[12] = in1[35] & in2[35];
    assign P[12] = in1[35] ^ in2[35];
    assign G[13] = in1[34] & in2[34];
    assign P[13] = in1[34] ^ in2[34];
    assign G[14] = in1[33] & in2[33];
    assign P[14] = in1[33] ^ in2[33];
    assign G[15] = in1[32] & in2[32];
    assign P[15] = in1[32] ^ in2[32];
    assign G[16] = in1[31] & in2[31];
    assign P[16] = in1[31] ^ in2[31];
    assign G[17] = in1[30] & in2[30];
    assign P[17] = in1[30] ^ in2[30];
    assign G[18] = in1[29] & in2[29];
    assign P[18] = in1[29] ^ in2[29];
    assign G[19] = in1[28] & in2[28];
    assign P[19] = in1[28] ^ in2[28];
    assign G[20] = in1[27] & in2[27];
    assign P[20] = in1[27] ^ in2[27];
    assign G[21] = in1[26] & in2[26];
    assign P[21] = in1[26] ^ in2[26];
    assign G[22] = in1[25] & in2[25];
    assign P[22] = in1[25] ^ in2[25];
    assign G[23] = in1[24] & in2[24];
    assign P[23] = in1[24] ^ in2[24];
    assign G[24] = in1[23] & in2[23];
    assign P[24] = in1[23] ^ in2[23];
    assign G[25] = in1[22] & in2[22];
    assign P[25] = in1[22] ^ in2[22];
    assign G[26] = in1[21] & in2[21];
    assign P[26] = in1[21] ^ in2[21];
    assign G[27] = in1[20] & in2[20];
    assign P[27] = in1[20] ^ in2[20];
    assign G[28] = in1[19] & in2[19];
    assign P[28] = in1[19] ^ in2[19];
    assign G[29] = in1[18] & in2[18];
    assign P[29] = in1[18] ^ in2[18];
    assign G[30] = in1[17] & in2[17];
    assign P[30] = in1[17] ^ in2[17];
    assign G[31] = in1[16] & in2[16];
    assign P[31] = in1[16] ^ in2[16];
    assign G[32] = in1[15] & in2[15];
    assign P[32] = in1[15] ^ in2[15];
    assign G[33] = in1[14] & in2[14];
    assign P[33] = in1[14] ^ in2[14];
    assign G[34] = in1[13] & in2[13];
    assign P[34] = in1[13] ^ in2[13];
    assign G[35] = in1[12] & in2[12];
    assign P[35] = in1[12] ^ in2[12];
    assign G[36] = in1[11] & in2[11];
    assign P[36] = in1[11] ^ in2[11];
    assign G[37] = in1[10] & in2[10];
    assign P[37] = in1[10] ^ in2[10];
    assign G[38] = in1[9] & in2[9];
    assign P[38] = in1[9] ^ in2[9];
    assign G[39] = in1[8] & in2[8];
    assign P[39] = in1[8] ^ in2[8];
    assign G[40] = in1[7] & in2[7];
    assign P[40] = in1[7] ^ in2[7];
    assign G[41] = in1[6] & in2[6];
    assign P[41] = in1[6] ^ in2[6];
    assign G[42] = in1[5] & in2[5];
    assign P[42] = in1[5] ^ in2[5];
    assign G[43] = in1[4] & in2[4];
    assign P[43] = in1[4] ^ in2[4];
    assign G[44] = in1[3] & in2[3];
    assign P[44] = in1[3] ^ in2[3];
    assign G[45] = in1[2] & in2[2];
    assign P[45] = in1[2] ^ in2[2];
    assign G[46] = in1[1] & in2[1];
    assign P[46] = in1[1] ^ in2[1];
    assign G[47] = in1[0] & in2[0];
    assign P[47] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign cout = G[47] | (P[47] & C[47]);
    assign sum = P ^ C;
endmodule

module CLA_47(output [46:0] sum, output cout, input [46:0] in1, input [46:0] in2);

    wire[46:0] G;
    wire[46:0] C;
    wire[46:0] P;

    assign G[0] = in1[46] & in2[46];
    assign P[0] = in1[46] ^ in2[46];
    assign G[1] = in1[45] & in2[45];
    assign P[1] = in1[45] ^ in2[45];
    assign G[2] = in1[44] & in2[44];
    assign P[2] = in1[44] ^ in2[44];
    assign G[3] = in1[43] & in2[43];
    assign P[3] = in1[43] ^ in2[43];
    assign G[4] = in1[42] & in2[42];
    assign P[4] = in1[42] ^ in2[42];
    assign G[5] = in1[41] & in2[41];
    assign P[5] = in1[41] ^ in2[41];
    assign G[6] = in1[40] & in2[40];
    assign P[6] = in1[40] ^ in2[40];
    assign G[7] = in1[39] & in2[39];
    assign P[7] = in1[39] ^ in2[39];
    assign G[8] = in1[38] & in2[38];
    assign P[8] = in1[38] ^ in2[38];
    assign G[9] = in1[37] & in2[37];
    assign P[9] = in1[37] ^ in2[37];
    assign G[10] = in1[36] & in2[36];
    assign P[10] = in1[36] ^ in2[36];
    assign G[11] = in1[35] & in2[35];
    assign P[11] = in1[35] ^ in2[35];
    assign G[12] = in1[34] & in2[34];
    assign P[12] = in1[34] ^ in2[34];
    assign G[13] = in1[33] & in2[33];
    assign P[13] = in1[33] ^ in2[33];
    assign G[14] = in1[32] & in2[32];
    assign P[14] = in1[32] ^ in2[32];
    assign G[15] = in1[31] & in2[31];
    assign P[15] = in1[31] ^ in2[31];
    assign G[16] = in1[30] & in2[30];
    assign P[16] = in1[30] ^ in2[30];
    assign G[17] = in1[29] & in2[29];
    assign P[17] = in1[29] ^ in2[29];
    assign G[18] = in1[28] & in2[28];
    assign P[18] = in1[28] ^ in2[28];
    assign G[19] = in1[27] & in2[27];
    assign P[19] = in1[27] ^ in2[27];
    assign G[20] = in1[26] & in2[26];
    assign P[20] = in1[26] ^ in2[26];
    assign G[21] = in1[25] & in2[25];
    assign P[21] = in1[25] ^ in2[25];
    assign G[22] = in1[24] & in2[24];
    assign P[22] = in1[24] ^ in2[24];
    assign G[23] = in1[23] & in2[23];
    assign P[23] = in1[23] ^ in2[23];
    assign G[24] = in1[22] & in2[22];
    assign P[24] = in1[22] ^ in2[22];
    assign G[25] = in1[21] & in2[21];
    assign P[25] = in1[21] ^ in2[21];
    assign G[26] = in1[20] & in2[20];
    assign P[26] = in1[20] ^ in2[20];
    assign G[27] = in1[19] & in2[19];
    assign P[27] = in1[19] ^ in2[19];
    assign G[28] = in1[18] & in2[18];
    assign P[28] = in1[18] ^ in2[18];
    assign G[29] = in1[17] & in2[17];
    assign P[29] = in1[17] ^ in2[17];
    assign G[30] = in1[16] & in2[16];
    assign P[30] = in1[16] ^ in2[16];
    assign G[31] = in1[15] & in2[15];
    assign P[31] = in1[15] ^ in2[15];
    assign G[32] = in1[14] & in2[14];
    assign P[32] = in1[14] ^ in2[14];
    assign G[33] = in1[13] & in2[13];
    assign P[33] = in1[13] ^ in2[13];
    assign G[34] = in1[12] & in2[12];
    assign P[34] = in1[12] ^ in2[12];
    assign G[35] = in1[11] & in2[11];
    assign P[35] = in1[11] ^ in2[11];
    assign G[36] = in1[10] & in2[10];
    assign P[36] = in1[10] ^ in2[10];
    assign G[37] = in1[9] & in2[9];
    assign P[37] = in1[9] ^ in2[9];
    assign G[38] = in1[8] & in2[8];
    assign P[38] = in1[8] ^ in2[8];
    assign G[39] = in1[7] & in2[7];
    assign P[39] = in1[7] ^ in2[7];
    assign G[40] = in1[6] & in2[6];
    assign P[40] = in1[6] ^ in2[6];
    assign G[41] = in1[5] & in2[5];
    assign P[41] = in1[5] ^ in2[5];
    assign G[42] = in1[4] & in2[4];
    assign P[42] = in1[4] ^ in2[4];
    assign G[43] = in1[3] & in2[3];
    assign P[43] = in1[3] ^ in2[3];
    assign G[44] = in1[2] & in2[2];
    assign P[44] = in1[2] ^ in2[2];
    assign G[45] = in1[1] & in2[1];
    assign P[45] = in1[1] ^ in2[1];
    assign G[46] = in1[0] & in2[0];
    assign P[46] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign cout = G[46] | (P[46] & C[46]);
    assign sum = P ^ C;
endmodule

module CLA_46(output [45:0] sum, output cout, input [45:0] in1, input [45:0] in2);

    wire[45:0] G;
    wire[45:0] C;
    wire[45:0] P;

    assign G[0] = in1[45] & in2[45];
    assign P[0] = in1[45] ^ in2[45];
    assign G[1] = in1[44] & in2[44];
    assign P[1] = in1[44] ^ in2[44];
    assign G[2] = in1[43] & in2[43];
    assign P[2] = in1[43] ^ in2[43];
    assign G[3] = in1[42] & in2[42];
    assign P[3] = in1[42] ^ in2[42];
    assign G[4] = in1[41] & in2[41];
    assign P[4] = in1[41] ^ in2[41];
    assign G[5] = in1[40] & in2[40];
    assign P[5] = in1[40] ^ in2[40];
    assign G[6] = in1[39] & in2[39];
    assign P[6] = in1[39] ^ in2[39];
    assign G[7] = in1[38] & in2[38];
    assign P[7] = in1[38] ^ in2[38];
    assign G[8] = in1[37] & in2[37];
    assign P[8] = in1[37] ^ in2[37];
    assign G[9] = in1[36] & in2[36];
    assign P[9] = in1[36] ^ in2[36];
    assign G[10] = in1[35] & in2[35];
    assign P[10] = in1[35] ^ in2[35];
    assign G[11] = in1[34] & in2[34];
    assign P[11] = in1[34] ^ in2[34];
    assign G[12] = in1[33] & in2[33];
    assign P[12] = in1[33] ^ in2[33];
    assign G[13] = in1[32] & in2[32];
    assign P[13] = in1[32] ^ in2[32];
    assign G[14] = in1[31] & in2[31];
    assign P[14] = in1[31] ^ in2[31];
    assign G[15] = in1[30] & in2[30];
    assign P[15] = in1[30] ^ in2[30];
    assign G[16] = in1[29] & in2[29];
    assign P[16] = in1[29] ^ in2[29];
    assign G[17] = in1[28] & in2[28];
    assign P[17] = in1[28] ^ in2[28];
    assign G[18] = in1[27] & in2[27];
    assign P[18] = in1[27] ^ in2[27];
    assign G[19] = in1[26] & in2[26];
    assign P[19] = in1[26] ^ in2[26];
    assign G[20] = in1[25] & in2[25];
    assign P[20] = in1[25] ^ in2[25];
    assign G[21] = in1[24] & in2[24];
    assign P[21] = in1[24] ^ in2[24];
    assign G[22] = in1[23] & in2[23];
    assign P[22] = in1[23] ^ in2[23];
    assign G[23] = in1[22] & in2[22];
    assign P[23] = in1[22] ^ in2[22];
    assign G[24] = in1[21] & in2[21];
    assign P[24] = in1[21] ^ in2[21];
    assign G[25] = in1[20] & in2[20];
    assign P[25] = in1[20] ^ in2[20];
    assign G[26] = in1[19] & in2[19];
    assign P[26] = in1[19] ^ in2[19];
    assign G[27] = in1[18] & in2[18];
    assign P[27] = in1[18] ^ in2[18];
    assign G[28] = in1[17] & in2[17];
    assign P[28] = in1[17] ^ in2[17];
    assign G[29] = in1[16] & in2[16];
    assign P[29] = in1[16] ^ in2[16];
    assign G[30] = in1[15] & in2[15];
    assign P[30] = in1[15] ^ in2[15];
    assign G[31] = in1[14] & in2[14];
    assign P[31] = in1[14] ^ in2[14];
    assign G[32] = in1[13] & in2[13];
    assign P[32] = in1[13] ^ in2[13];
    assign G[33] = in1[12] & in2[12];
    assign P[33] = in1[12] ^ in2[12];
    assign G[34] = in1[11] & in2[11];
    assign P[34] = in1[11] ^ in2[11];
    assign G[35] = in1[10] & in2[10];
    assign P[35] = in1[10] ^ in2[10];
    assign G[36] = in1[9] & in2[9];
    assign P[36] = in1[9] ^ in2[9];
    assign G[37] = in1[8] & in2[8];
    assign P[37] = in1[8] ^ in2[8];
    assign G[38] = in1[7] & in2[7];
    assign P[38] = in1[7] ^ in2[7];
    assign G[39] = in1[6] & in2[6];
    assign P[39] = in1[6] ^ in2[6];
    assign G[40] = in1[5] & in2[5];
    assign P[40] = in1[5] ^ in2[5];
    assign G[41] = in1[4] & in2[4];
    assign P[41] = in1[4] ^ in2[4];
    assign G[42] = in1[3] & in2[3];
    assign P[42] = in1[3] ^ in2[3];
    assign G[43] = in1[2] & in2[2];
    assign P[43] = in1[2] ^ in2[2];
    assign G[44] = in1[1] & in2[1];
    assign P[44] = in1[1] ^ in2[1];
    assign G[45] = in1[0] & in2[0];
    assign P[45] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign cout = G[45] | (P[45] & C[45]);
    assign sum = P ^ C;
endmodule

module CLA_45(output [44:0] sum, output cout, input [44:0] in1, input [44:0] in2);

    wire[44:0] G;
    wire[44:0] C;
    wire[44:0] P;

    assign G[0] = in1[44] & in2[44];
    assign P[0] = in1[44] ^ in2[44];
    assign G[1] = in1[43] & in2[43];
    assign P[1] = in1[43] ^ in2[43];
    assign G[2] = in1[42] & in2[42];
    assign P[2] = in1[42] ^ in2[42];
    assign G[3] = in1[41] & in2[41];
    assign P[3] = in1[41] ^ in2[41];
    assign G[4] = in1[40] & in2[40];
    assign P[4] = in1[40] ^ in2[40];
    assign G[5] = in1[39] & in2[39];
    assign P[5] = in1[39] ^ in2[39];
    assign G[6] = in1[38] & in2[38];
    assign P[6] = in1[38] ^ in2[38];
    assign G[7] = in1[37] & in2[37];
    assign P[7] = in1[37] ^ in2[37];
    assign G[8] = in1[36] & in2[36];
    assign P[8] = in1[36] ^ in2[36];
    assign G[9] = in1[35] & in2[35];
    assign P[9] = in1[35] ^ in2[35];
    assign G[10] = in1[34] & in2[34];
    assign P[10] = in1[34] ^ in2[34];
    assign G[11] = in1[33] & in2[33];
    assign P[11] = in1[33] ^ in2[33];
    assign G[12] = in1[32] & in2[32];
    assign P[12] = in1[32] ^ in2[32];
    assign G[13] = in1[31] & in2[31];
    assign P[13] = in1[31] ^ in2[31];
    assign G[14] = in1[30] & in2[30];
    assign P[14] = in1[30] ^ in2[30];
    assign G[15] = in1[29] & in2[29];
    assign P[15] = in1[29] ^ in2[29];
    assign G[16] = in1[28] & in2[28];
    assign P[16] = in1[28] ^ in2[28];
    assign G[17] = in1[27] & in2[27];
    assign P[17] = in1[27] ^ in2[27];
    assign G[18] = in1[26] & in2[26];
    assign P[18] = in1[26] ^ in2[26];
    assign G[19] = in1[25] & in2[25];
    assign P[19] = in1[25] ^ in2[25];
    assign G[20] = in1[24] & in2[24];
    assign P[20] = in1[24] ^ in2[24];
    assign G[21] = in1[23] & in2[23];
    assign P[21] = in1[23] ^ in2[23];
    assign G[22] = in1[22] & in2[22];
    assign P[22] = in1[22] ^ in2[22];
    assign G[23] = in1[21] & in2[21];
    assign P[23] = in1[21] ^ in2[21];
    assign G[24] = in1[20] & in2[20];
    assign P[24] = in1[20] ^ in2[20];
    assign G[25] = in1[19] & in2[19];
    assign P[25] = in1[19] ^ in2[19];
    assign G[26] = in1[18] & in2[18];
    assign P[26] = in1[18] ^ in2[18];
    assign G[27] = in1[17] & in2[17];
    assign P[27] = in1[17] ^ in2[17];
    assign G[28] = in1[16] & in2[16];
    assign P[28] = in1[16] ^ in2[16];
    assign G[29] = in1[15] & in2[15];
    assign P[29] = in1[15] ^ in2[15];
    assign G[30] = in1[14] & in2[14];
    assign P[30] = in1[14] ^ in2[14];
    assign G[31] = in1[13] & in2[13];
    assign P[31] = in1[13] ^ in2[13];
    assign G[32] = in1[12] & in2[12];
    assign P[32] = in1[12] ^ in2[12];
    assign G[33] = in1[11] & in2[11];
    assign P[33] = in1[11] ^ in2[11];
    assign G[34] = in1[10] & in2[10];
    assign P[34] = in1[10] ^ in2[10];
    assign G[35] = in1[9] & in2[9];
    assign P[35] = in1[9] ^ in2[9];
    assign G[36] = in1[8] & in2[8];
    assign P[36] = in1[8] ^ in2[8];
    assign G[37] = in1[7] & in2[7];
    assign P[37] = in1[7] ^ in2[7];
    assign G[38] = in1[6] & in2[6];
    assign P[38] = in1[6] ^ in2[6];
    assign G[39] = in1[5] & in2[5];
    assign P[39] = in1[5] ^ in2[5];
    assign G[40] = in1[4] & in2[4];
    assign P[40] = in1[4] ^ in2[4];
    assign G[41] = in1[3] & in2[3];
    assign P[41] = in1[3] ^ in2[3];
    assign G[42] = in1[2] & in2[2];
    assign P[42] = in1[2] ^ in2[2];
    assign G[43] = in1[1] & in2[1];
    assign P[43] = in1[1] ^ in2[1];
    assign G[44] = in1[0] & in2[0];
    assign P[44] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign cout = G[44] | (P[44] & C[44]);
    assign sum = P ^ C;
endmodule

module CLA_44(output [43:0] sum, output cout, input [43:0] in1, input [43:0] in2);

    wire[43:0] G;
    wire[43:0] C;
    wire[43:0] P;

    assign G[0] = in1[43] & in2[43];
    assign P[0] = in1[43] ^ in2[43];
    assign G[1] = in1[42] & in2[42];
    assign P[1] = in1[42] ^ in2[42];
    assign G[2] = in1[41] & in2[41];
    assign P[2] = in1[41] ^ in2[41];
    assign G[3] = in1[40] & in2[40];
    assign P[3] = in1[40] ^ in2[40];
    assign G[4] = in1[39] & in2[39];
    assign P[4] = in1[39] ^ in2[39];
    assign G[5] = in1[38] & in2[38];
    assign P[5] = in1[38] ^ in2[38];
    assign G[6] = in1[37] & in2[37];
    assign P[6] = in1[37] ^ in2[37];
    assign G[7] = in1[36] & in2[36];
    assign P[7] = in1[36] ^ in2[36];
    assign G[8] = in1[35] & in2[35];
    assign P[8] = in1[35] ^ in2[35];
    assign G[9] = in1[34] & in2[34];
    assign P[9] = in1[34] ^ in2[34];
    assign G[10] = in1[33] & in2[33];
    assign P[10] = in1[33] ^ in2[33];
    assign G[11] = in1[32] & in2[32];
    assign P[11] = in1[32] ^ in2[32];
    assign G[12] = in1[31] & in2[31];
    assign P[12] = in1[31] ^ in2[31];
    assign G[13] = in1[30] & in2[30];
    assign P[13] = in1[30] ^ in2[30];
    assign G[14] = in1[29] & in2[29];
    assign P[14] = in1[29] ^ in2[29];
    assign G[15] = in1[28] & in2[28];
    assign P[15] = in1[28] ^ in2[28];
    assign G[16] = in1[27] & in2[27];
    assign P[16] = in1[27] ^ in2[27];
    assign G[17] = in1[26] & in2[26];
    assign P[17] = in1[26] ^ in2[26];
    assign G[18] = in1[25] & in2[25];
    assign P[18] = in1[25] ^ in2[25];
    assign G[19] = in1[24] & in2[24];
    assign P[19] = in1[24] ^ in2[24];
    assign G[20] = in1[23] & in2[23];
    assign P[20] = in1[23] ^ in2[23];
    assign G[21] = in1[22] & in2[22];
    assign P[21] = in1[22] ^ in2[22];
    assign G[22] = in1[21] & in2[21];
    assign P[22] = in1[21] ^ in2[21];
    assign G[23] = in1[20] & in2[20];
    assign P[23] = in1[20] ^ in2[20];
    assign G[24] = in1[19] & in2[19];
    assign P[24] = in1[19] ^ in2[19];
    assign G[25] = in1[18] & in2[18];
    assign P[25] = in1[18] ^ in2[18];
    assign G[26] = in1[17] & in2[17];
    assign P[26] = in1[17] ^ in2[17];
    assign G[27] = in1[16] & in2[16];
    assign P[27] = in1[16] ^ in2[16];
    assign G[28] = in1[15] & in2[15];
    assign P[28] = in1[15] ^ in2[15];
    assign G[29] = in1[14] & in2[14];
    assign P[29] = in1[14] ^ in2[14];
    assign G[30] = in1[13] & in2[13];
    assign P[30] = in1[13] ^ in2[13];
    assign G[31] = in1[12] & in2[12];
    assign P[31] = in1[12] ^ in2[12];
    assign G[32] = in1[11] & in2[11];
    assign P[32] = in1[11] ^ in2[11];
    assign G[33] = in1[10] & in2[10];
    assign P[33] = in1[10] ^ in2[10];
    assign G[34] = in1[9] & in2[9];
    assign P[34] = in1[9] ^ in2[9];
    assign G[35] = in1[8] & in2[8];
    assign P[35] = in1[8] ^ in2[8];
    assign G[36] = in1[7] & in2[7];
    assign P[36] = in1[7] ^ in2[7];
    assign G[37] = in1[6] & in2[6];
    assign P[37] = in1[6] ^ in2[6];
    assign G[38] = in1[5] & in2[5];
    assign P[38] = in1[5] ^ in2[5];
    assign G[39] = in1[4] & in2[4];
    assign P[39] = in1[4] ^ in2[4];
    assign G[40] = in1[3] & in2[3];
    assign P[40] = in1[3] ^ in2[3];
    assign G[41] = in1[2] & in2[2];
    assign P[41] = in1[2] ^ in2[2];
    assign G[42] = in1[1] & in2[1];
    assign P[42] = in1[1] ^ in2[1];
    assign G[43] = in1[0] & in2[0];
    assign P[43] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign cout = G[43] | (P[43] & C[43]);
    assign sum = P ^ C;
endmodule

module CLA_43(output [42:0] sum, output cout, input [42:0] in1, input [42:0] in2);

    wire[42:0] G;
    wire[42:0] C;
    wire[42:0] P;

    assign G[0] = in1[42] & in2[42];
    assign P[0] = in1[42] ^ in2[42];
    assign G[1] = in1[41] & in2[41];
    assign P[1] = in1[41] ^ in2[41];
    assign G[2] = in1[40] & in2[40];
    assign P[2] = in1[40] ^ in2[40];
    assign G[3] = in1[39] & in2[39];
    assign P[3] = in1[39] ^ in2[39];
    assign G[4] = in1[38] & in2[38];
    assign P[4] = in1[38] ^ in2[38];
    assign G[5] = in1[37] & in2[37];
    assign P[5] = in1[37] ^ in2[37];
    assign G[6] = in1[36] & in2[36];
    assign P[6] = in1[36] ^ in2[36];
    assign G[7] = in1[35] & in2[35];
    assign P[7] = in1[35] ^ in2[35];
    assign G[8] = in1[34] & in2[34];
    assign P[8] = in1[34] ^ in2[34];
    assign G[9] = in1[33] & in2[33];
    assign P[9] = in1[33] ^ in2[33];
    assign G[10] = in1[32] & in2[32];
    assign P[10] = in1[32] ^ in2[32];
    assign G[11] = in1[31] & in2[31];
    assign P[11] = in1[31] ^ in2[31];
    assign G[12] = in1[30] & in2[30];
    assign P[12] = in1[30] ^ in2[30];
    assign G[13] = in1[29] & in2[29];
    assign P[13] = in1[29] ^ in2[29];
    assign G[14] = in1[28] & in2[28];
    assign P[14] = in1[28] ^ in2[28];
    assign G[15] = in1[27] & in2[27];
    assign P[15] = in1[27] ^ in2[27];
    assign G[16] = in1[26] & in2[26];
    assign P[16] = in1[26] ^ in2[26];
    assign G[17] = in1[25] & in2[25];
    assign P[17] = in1[25] ^ in2[25];
    assign G[18] = in1[24] & in2[24];
    assign P[18] = in1[24] ^ in2[24];
    assign G[19] = in1[23] & in2[23];
    assign P[19] = in1[23] ^ in2[23];
    assign G[20] = in1[22] & in2[22];
    assign P[20] = in1[22] ^ in2[22];
    assign G[21] = in1[21] & in2[21];
    assign P[21] = in1[21] ^ in2[21];
    assign G[22] = in1[20] & in2[20];
    assign P[22] = in1[20] ^ in2[20];
    assign G[23] = in1[19] & in2[19];
    assign P[23] = in1[19] ^ in2[19];
    assign G[24] = in1[18] & in2[18];
    assign P[24] = in1[18] ^ in2[18];
    assign G[25] = in1[17] & in2[17];
    assign P[25] = in1[17] ^ in2[17];
    assign G[26] = in1[16] & in2[16];
    assign P[26] = in1[16] ^ in2[16];
    assign G[27] = in1[15] & in2[15];
    assign P[27] = in1[15] ^ in2[15];
    assign G[28] = in1[14] & in2[14];
    assign P[28] = in1[14] ^ in2[14];
    assign G[29] = in1[13] & in2[13];
    assign P[29] = in1[13] ^ in2[13];
    assign G[30] = in1[12] & in2[12];
    assign P[30] = in1[12] ^ in2[12];
    assign G[31] = in1[11] & in2[11];
    assign P[31] = in1[11] ^ in2[11];
    assign G[32] = in1[10] & in2[10];
    assign P[32] = in1[10] ^ in2[10];
    assign G[33] = in1[9] & in2[9];
    assign P[33] = in1[9] ^ in2[9];
    assign G[34] = in1[8] & in2[8];
    assign P[34] = in1[8] ^ in2[8];
    assign G[35] = in1[7] & in2[7];
    assign P[35] = in1[7] ^ in2[7];
    assign G[36] = in1[6] & in2[6];
    assign P[36] = in1[6] ^ in2[6];
    assign G[37] = in1[5] & in2[5];
    assign P[37] = in1[5] ^ in2[5];
    assign G[38] = in1[4] & in2[4];
    assign P[38] = in1[4] ^ in2[4];
    assign G[39] = in1[3] & in2[3];
    assign P[39] = in1[3] ^ in2[3];
    assign G[40] = in1[2] & in2[2];
    assign P[40] = in1[2] ^ in2[2];
    assign G[41] = in1[1] & in2[1];
    assign P[41] = in1[1] ^ in2[1];
    assign G[42] = in1[0] & in2[0];
    assign P[42] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign cout = G[42] | (P[42] & C[42]);
    assign sum = P ^ C;
endmodule

module CLA_42(output [41:0] sum, output cout, input [41:0] in1, input [41:0] in2);

    wire[41:0] G;
    wire[41:0] C;
    wire[41:0] P;

    assign G[0] = in1[41] & in2[41];
    assign P[0] = in1[41] ^ in2[41];
    assign G[1] = in1[40] & in2[40];
    assign P[1] = in1[40] ^ in2[40];
    assign G[2] = in1[39] & in2[39];
    assign P[2] = in1[39] ^ in2[39];
    assign G[3] = in1[38] & in2[38];
    assign P[3] = in1[38] ^ in2[38];
    assign G[4] = in1[37] & in2[37];
    assign P[4] = in1[37] ^ in2[37];
    assign G[5] = in1[36] & in2[36];
    assign P[5] = in1[36] ^ in2[36];
    assign G[6] = in1[35] & in2[35];
    assign P[6] = in1[35] ^ in2[35];
    assign G[7] = in1[34] & in2[34];
    assign P[7] = in1[34] ^ in2[34];
    assign G[8] = in1[33] & in2[33];
    assign P[8] = in1[33] ^ in2[33];
    assign G[9] = in1[32] & in2[32];
    assign P[9] = in1[32] ^ in2[32];
    assign G[10] = in1[31] & in2[31];
    assign P[10] = in1[31] ^ in2[31];
    assign G[11] = in1[30] & in2[30];
    assign P[11] = in1[30] ^ in2[30];
    assign G[12] = in1[29] & in2[29];
    assign P[12] = in1[29] ^ in2[29];
    assign G[13] = in1[28] & in2[28];
    assign P[13] = in1[28] ^ in2[28];
    assign G[14] = in1[27] & in2[27];
    assign P[14] = in1[27] ^ in2[27];
    assign G[15] = in1[26] & in2[26];
    assign P[15] = in1[26] ^ in2[26];
    assign G[16] = in1[25] & in2[25];
    assign P[16] = in1[25] ^ in2[25];
    assign G[17] = in1[24] & in2[24];
    assign P[17] = in1[24] ^ in2[24];
    assign G[18] = in1[23] & in2[23];
    assign P[18] = in1[23] ^ in2[23];
    assign G[19] = in1[22] & in2[22];
    assign P[19] = in1[22] ^ in2[22];
    assign G[20] = in1[21] & in2[21];
    assign P[20] = in1[21] ^ in2[21];
    assign G[21] = in1[20] & in2[20];
    assign P[21] = in1[20] ^ in2[20];
    assign G[22] = in1[19] & in2[19];
    assign P[22] = in1[19] ^ in2[19];
    assign G[23] = in1[18] & in2[18];
    assign P[23] = in1[18] ^ in2[18];
    assign G[24] = in1[17] & in2[17];
    assign P[24] = in1[17] ^ in2[17];
    assign G[25] = in1[16] & in2[16];
    assign P[25] = in1[16] ^ in2[16];
    assign G[26] = in1[15] & in2[15];
    assign P[26] = in1[15] ^ in2[15];
    assign G[27] = in1[14] & in2[14];
    assign P[27] = in1[14] ^ in2[14];
    assign G[28] = in1[13] & in2[13];
    assign P[28] = in1[13] ^ in2[13];
    assign G[29] = in1[12] & in2[12];
    assign P[29] = in1[12] ^ in2[12];
    assign G[30] = in1[11] & in2[11];
    assign P[30] = in1[11] ^ in2[11];
    assign G[31] = in1[10] & in2[10];
    assign P[31] = in1[10] ^ in2[10];
    assign G[32] = in1[9] & in2[9];
    assign P[32] = in1[9] ^ in2[9];
    assign G[33] = in1[8] & in2[8];
    assign P[33] = in1[8] ^ in2[8];
    assign G[34] = in1[7] & in2[7];
    assign P[34] = in1[7] ^ in2[7];
    assign G[35] = in1[6] & in2[6];
    assign P[35] = in1[6] ^ in2[6];
    assign G[36] = in1[5] & in2[5];
    assign P[36] = in1[5] ^ in2[5];
    assign G[37] = in1[4] & in2[4];
    assign P[37] = in1[4] ^ in2[4];
    assign G[38] = in1[3] & in2[3];
    assign P[38] = in1[3] ^ in2[3];
    assign G[39] = in1[2] & in2[2];
    assign P[39] = in1[2] ^ in2[2];
    assign G[40] = in1[1] & in2[1];
    assign P[40] = in1[1] ^ in2[1];
    assign G[41] = in1[0] & in2[0];
    assign P[41] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign cout = G[41] | (P[41] & C[41]);
    assign sum = P ^ C;
endmodule

module CLA_41(output [40:0] sum, output cout, input [40:0] in1, input [40:0] in2);

    wire[40:0] G;
    wire[40:0] C;
    wire[40:0] P;

    assign G[0] = in1[40] & in2[40];
    assign P[0] = in1[40] ^ in2[40];
    assign G[1] = in1[39] & in2[39];
    assign P[1] = in1[39] ^ in2[39];
    assign G[2] = in1[38] & in2[38];
    assign P[2] = in1[38] ^ in2[38];
    assign G[3] = in1[37] & in2[37];
    assign P[3] = in1[37] ^ in2[37];
    assign G[4] = in1[36] & in2[36];
    assign P[4] = in1[36] ^ in2[36];
    assign G[5] = in1[35] & in2[35];
    assign P[5] = in1[35] ^ in2[35];
    assign G[6] = in1[34] & in2[34];
    assign P[6] = in1[34] ^ in2[34];
    assign G[7] = in1[33] & in2[33];
    assign P[7] = in1[33] ^ in2[33];
    assign G[8] = in1[32] & in2[32];
    assign P[8] = in1[32] ^ in2[32];
    assign G[9] = in1[31] & in2[31];
    assign P[9] = in1[31] ^ in2[31];
    assign G[10] = in1[30] & in2[30];
    assign P[10] = in1[30] ^ in2[30];
    assign G[11] = in1[29] & in2[29];
    assign P[11] = in1[29] ^ in2[29];
    assign G[12] = in1[28] & in2[28];
    assign P[12] = in1[28] ^ in2[28];
    assign G[13] = in1[27] & in2[27];
    assign P[13] = in1[27] ^ in2[27];
    assign G[14] = in1[26] & in2[26];
    assign P[14] = in1[26] ^ in2[26];
    assign G[15] = in1[25] & in2[25];
    assign P[15] = in1[25] ^ in2[25];
    assign G[16] = in1[24] & in2[24];
    assign P[16] = in1[24] ^ in2[24];
    assign G[17] = in1[23] & in2[23];
    assign P[17] = in1[23] ^ in2[23];
    assign G[18] = in1[22] & in2[22];
    assign P[18] = in1[22] ^ in2[22];
    assign G[19] = in1[21] & in2[21];
    assign P[19] = in1[21] ^ in2[21];
    assign G[20] = in1[20] & in2[20];
    assign P[20] = in1[20] ^ in2[20];
    assign G[21] = in1[19] & in2[19];
    assign P[21] = in1[19] ^ in2[19];
    assign G[22] = in1[18] & in2[18];
    assign P[22] = in1[18] ^ in2[18];
    assign G[23] = in1[17] & in2[17];
    assign P[23] = in1[17] ^ in2[17];
    assign G[24] = in1[16] & in2[16];
    assign P[24] = in1[16] ^ in2[16];
    assign G[25] = in1[15] & in2[15];
    assign P[25] = in1[15] ^ in2[15];
    assign G[26] = in1[14] & in2[14];
    assign P[26] = in1[14] ^ in2[14];
    assign G[27] = in1[13] & in2[13];
    assign P[27] = in1[13] ^ in2[13];
    assign G[28] = in1[12] & in2[12];
    assign P[28] = in1[12] ^ in2[12];
    assign G[29] = in1[11] & in2[11];
    assign P[29] = in1[11] ^ in2[11];
    assign G[30] = in1[10] & in2[10];
    assign P[30] = in1[10] ^ in2[10];
    assign G[31] = in1[9] & in2[9];
    assign P[31] = in1[9] ^ in2[9];
    assign G[32] = in1[8] & in2[8];
    assign P[32] = in1[8] ^ in2[8];
    assign G[33] = in1[7] & in2[7];
    assign P[33] = in1[7] ^ in2[7];
    assign G[34] = in1[6] & in2[6];
    assign P[34] = in1[6] ^ in2[6];
    assign G[35] = in1[5] & in2[5];
    assign P[35] = in1[5] ^ in2[5];
    assign G[36] = in1[4] & in2[4];
    assign P[36] = in1[4] ^ in2[4];
    assign G[37] = in1[3] & in2[3];
    assign P[37] = in1[3] ^ in2[3];
    assign G[38] = in1[2] & in2[2];
    assign P[38] = in1[2] ^ in2[2];
    assign G[39] = in1[1] & in2[1];
    assign P[39] = in1[1] ^ in2[1];
    assign G[40] = in1[0] & in2[0];
    assign P[40] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign cout = G[40] | (P[40] & C[40]);
    assign sum = P ^ C;
endmodule

module CLA_40(output [39:0] sum, output cout, input [39:0] in1, input [39:0] in2);

    wire[39:0] G;
    wire[39:0] C;
    wire[39:0] P;

    assign G[0] = in1[39] & in2[39];
    assign P[0] = in1[39] ^ in2[39];
    assign G[1] = in1[38] & in2[38];
    assign P[1] = in1[38] ^ in2[38];
    assign G[2] = in1[37] & in2[37];
    assign P[2] = in1[37] ^ in2[37];
    assign G[3] = in1[36] & in2[36];
    assign P[3] = in1[36] ^ in2[36];
    assign G[4] = in1[35] & in2[35];
    assign P[4] = in1[35] ^ in2[35];
    assign G[5] = in1[34] & in2[34];
    assign P[5] = in1[34] ^ in2[34];
    assign G[6] = in1[33] & in2[33];
    assign P[6] = in1[33] ^ in2[33];
    assign G[7] = in1[32] & in2[32];
    assign P[7] = in1[32] ^ in2[32];
    assign G[8] = in1[31] & in2[31];
    assign P[8] = in1[31] ^ in2[31];
    assign G[9] = in1[30] & in2[30];
    assign P[9] = in1[30] ^ in2[30];
    assign G[10] = in1[29] & in2[29];
    assign P[10] = in1[29] ^ in2[29];
    assign G[11] = in1[28] & in2[28];
    assign P[11] = in1[28] ^ in2[28];
    assign G[12] = in1[27] & in2[27];
    assign P[12] = in1[27] ^ in2[27];
    assign G[13] = in1[26] & in2[26];
    assign P[13] = in1[26] ^ in2[26];
    assign G[14] = in1[25] & in2[25];
    assign P[14] = in1[25] ^ in2[25];
    assign G[15] = in1[24] & in2[24];
    assign P[15] = in1[24] ^ in2[24];
    assign G[16] = in1[23] & in2[23];
    assign P[16] = in1[23] ^ in2[23];
    assign G[17] = in1[22] & in2[22];
    assign P[17] = in1[22] ^ in2[22];
    assign G[18] = in1[21] & in2[21];
    assign P[18] = in1[21] ^ in2[21];
    assign G[19] = in1[20] & in2[20];
    assign P[19] = in1[20] ^ in2[20];
    assign G[20] = in1[19] & in2[19];
    assign P[20] = in1[19] ^ in2[19];
    assign G[21] = in1[18] & in2[18];
    assign P[21] = in1[18] ^ in2[18];
    assign G[22] = in1[17] & in2[17];
    assign P[22] = in1[17] ^ in2[17];
    assign G[23] = in1[16] & in2[16];
    assign P[23] = in1[16] ^ in2[16];
    assign G[24] = in1[15] & in2[15];
    assign P[24] = in1[15] ^ in2[15];
    assign G[25] = in1[14] & in2[14];
    assign P[25] = in1[14] ^ in2[14];
    assign G[26] = in1[13] & in2[13];
    assign P[26] = in1[13] ^ in2[13];
    assign G[27] = in1[12] & in2[12];
    assign P[27] = in1[12] ^ in2[12];
    assign G[28] = in1[11] & in2[11];
    assign P[28] = in1[11] ^ in2[11];
    assign G[29] = in1[10] & in2[10];
    assign P[29] = in1[10] ^ in2[10];
    assign G[30] = in1[9] & in2[9];
    assign P[30] = in1[9] ^ in2[9];
    assign G[31] = in1[8] & in2[8];
    assign P[31] = in1[8] ^ in2[8];
    assign G[32] = in1[7] & in2[7];
    assign P[32] = in1[7] ^ in2[7];
    assign G[33] = in1[6] & in2[6];
    assign P[33] = in1[6] ^ in2[6];
    assign G[34] = in1[5] & in2[5];
    assign P[34] = in1[5] ^ in2[5];
    assign G[35] = in1[4] & in2[4];
    assign P[35] = in1[4] ^ in2[4];
    assign G[36] = in1[3] & in2[3];
    assign P[36] = in1[3] ^ in2[3];
    assign G[37] = in1[2] & in2[2];
    assign P[37] = in1[2] ^ in2[2];
    assign G[38] = in1[1] & in2[1];
    assign P[38] = in1[1] ^ in2[1];
    assign G[39] = in1[0] & in2[0];
    assign P[39] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign cout = G[39] | (P[39] & C[39]);
    assign sum = P ^ C;
endmodule

module CLA_39(output [38:0] sum, output cout, input [38:0] in1, input [38:0] in2);

    wire[38:0] G;
    wire[38:0] C;
    wire[38:0] P;

    assign G[0] = in1[38] & in2[38];
    assign P[0] = in1[38] ^ in2[38];
    assign G[1] = in1[37] & in2[37];
    assign P[1] = in1[37] ^ in2[37];
    assign G[2] = in1[36] & in2[36];
    assign P[2] = in1[36] ^ in2[36];
    assign G[3] = in1[35] & in2[35];
    assign P[3] = in1[35] ^ in2[35];
    assign G[4] = in1[34] & in2[34];
    assign P[4] = in1[34] ^ in2[34];
    assign G[5] = in1[33] & in2[33];
    assign P[5] = in1[33] ^ in2[33];
    assign G[6] = in1[32] & in2[32];
    assign P[6] = in1[32] ^ in2[32];
    assign G[7] = in1[31] & in2[31];
    assign P[7] = in1[31] ^ in2[31];
    assign G[8] = in1[30] & in2[30];
    assign P[8] = in1[30] ^ in2[30];
    assign G[9] = in1[29] & in2[29];
    assign P[9] = in1[29] ^ in2[29];
    assign G[10] = in1[28] & in2[28];
    assign P[10] = in1[28] ^ in2[28];
    assign G[11] = in1[27] & in2[27];
    assign P[11] = in1[27] ^ in2[27];
    assign G[12] = in1[26] & in2[26];
    assign P[12] = in1[26] ^ in2[26];
    assign G[13] = in1[25] & in2[25];
    assign P[13] = in1[25] ^ in2[25];
    assign G[14] = in1[24] & in2[24];
    assign P[14] = in1[24] ^ in2[24];
    assign G[15] = in1[23] & in2[23];
    assign P[15] = in1[23] ^ in2[23];
    assign G[16] = in1[22] & in2[22];
    assign P[16] = in1[22] ^ in2[22];
    assign G[17] = in1[21] & in2[21];
    assign P[17] = in1[21] ^ in2[21];
    assign G[18] = in1[20] & in2[20];
    assign P[18] = in1[20] ^ in2[20];
    assign G[19] = in1[19] & in2[19];
    assign P[19] = in1[19] ^ in2[19];
    assign G[20] = in1[18] & in2[18];
    assign P[20] = in1[18] ^ in2[18];
    assign G[21] = in1[17] & in2[17];
    assign P[21] = in1[17] ^ in2[17];
    assign G[22] = in1[16] & in2[16];
    assign P[22] = in1[16] ^ in2[16];
    assign G[23] = in1[15] & in2[15];
    assign P[23] = in1[15] ^ in2[15];
    assign G[24] = in1[14] & in2[14];
    assign P[24] = in1[14] ^ in2[14];
    assign G[25] = in1[13] & in2[13];
    assign P[25] = in1[13] ^ in2[13];
    assign G[26] = in1[12] & in2[12];
    assign P[26] = in1[12] ^ in2[12];
    assign G[27] = in1[11] & in2[11];
    assign P[27] = in1[11] ^ in2[11];
    assign G[28] = in1[10] & in2[10];
    assign P[28] = in1[10] ^ in2[10];
    assign G[29] = in1[9] & in2[9];
    assign P[29] = in1[9] ^ in2[9];
    assign G[30] = in1[8] & in2[8];
    assign P[30] = in1[8] ^ in2[8];
    assign G[31] = in1[7] & in2[7];
    assign P[31] = in1[7] ^ in2[7];
    assign G[32] = in1[6] & in2[6];
    assign P[32] = in1[6] ^ in2[6];
    assign G[33] = in1[5] & in2[5];
    assign P[33] = in1[5] ^ in2[5];
    assign G[34] = in1[4] & in2[4];
    assign P[34] = in1[4] ^ in2[4];
    assign G[35] = in1[3] & in2[3];
    assign P[35] = in1[3] ^ in2[3];
    assign G[36] = in1[2] & in2[2];
    assign P[36] = in1[2] ^ in2[2];
    assign G[37] = in1[1] & in2[1];
    assign P[37] = in1[1] ^ in2[1];
    assign G[38] = in1[0] & in2[0];
    assign P[38] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign cout = G[38] | (P[38] & C[38]);
    assign sum = P ^ C;
endmodule

module CLA_38(output [37:0] sum, output cout, input [37:0] in1, input [37:0] in2);

    wire[37:0] G;
    wire[37:0] C;
    wire[37:0] P;

    assign G[0] = in1[37] & in2[37];
    assign P[0] = in1[37] ^ in2[37];
    assign G[1] = in1[36] & in2[36];
    assign P[1] = in1[36] ^ in2[36];
    assign G[2] = in1[35] & in2[35];
    assign P[2] = in1[35] ^ in2[35];
    assign G[3] = in1[34] & in2[34];
    assign P[3] = in1[34] ^ in2[34];
    assign G[4] = in1[33] & in2[33];
    assign P[4] = in1[33] ^ in2[33];
    assign G[5] = in1[32] & in2[32];
    assign P[5] = in1[32] ^ in2[32];
    assign G[6] = in1[31] & in2[31];
    assign P[6] = in1[31] ^ in2[31];
    assign G[7] = in1[30] & in2[30];
    assign P[7] = in1[30] ^ in2[30];
    assign G[8] = in1[29] & in2[29];
    assign P[8] = in1[29] ^ in2[29];
    assign G[9] = in1[28] & in2[28];
    assign P[9] = in1[28] ^ in2[28];
    assign G[10] = in1[27] & in2[27];
    assign P[10] = in1[27] ^ in2[27];
    assign G[11] = in1[26] & in2[26];
    assign P[11] = in1[26] ^ in2[26];
    assign G[12] = in1[25] & in2[25];
    assign P[12] = in1[25] ^ in2[25];
    assign G[13] = in1[24] & in2[24];
    assign P[13] = in1[24] ^ in2[24];
    assign G[14] = in1[23] & in2[23];
    assign P[14] = in1[23] ^ in2[23];
    assign G[15] = in1[22] & in2[22];
    assign P[15] = in1[22] ^ in2[22];
    assign G[16] = in1[21] & in2[21];
    assign P[16] = in1[21] ^ in2[21];
    assign G[17] = in1[20] & in2[20];
    assign P[17] = in1[20] ^ in2[20];
    assign G[18] = in1[19] & in2[19];
    assign P[18] = in1[19] ^ in2[19];
    assign G[19] = in1[18] & in2[18];
    assign P[19] = in1[18] ^ in2[18];
    assign G[20] = in1[17] & in2[17];
    assign P[20] = in1[17] ^ in2[17];
    assign G[21] = in1[16] & in2[16];
    assign P[21] = in1[16] ^ in2[16];
    assign G[22] = in1[15] & in2[15];
    assign P[22] = in1[15] ^ in2[15];
    assign G[23] = in1[14] & in2[14];
    assign P[23] = in1[14] ^ in2[14];
    assign G[24] = in1[13] & in2[13];
    assign P[24] = in1[13] ^ in2[13];
    assign G[25] = in1[12] & in2[12];
    assign P[25] = in1[12] ^ in2[12];
    assign G[26] = in1[11] & in2[11];
    assign P[26] = in1[11] ^ in2[11];
    assign G[27] = in1[10] & in2[10];
    assign P[27] = in1[10] ^ in2[10];
    assign G[28] = in1[9] & in2[9];
    assign P[28] = in1[9] ^ in2[9];
    assign G[29] = in1[8] & in2[8];
    assign P[29] = in1[8] ^ in2[8];
    assign G[30] = in1[7] & in2[7];
    assign P[30] = in1[7] ^ in2[7];
    assign G[31] = in1[6] & in2[6];
    assign P[31] = in1[6] ^ in2[6];
    assign G[32] = in1[5] & in2[5];
    assign P[32] = in1[5] ^ in2[5];
    assign G[33] = in1[4] & in2[4];
    assign P[33] = in1[4] ^ in2[4];
    assign G[34] = in1[3] & in2[3];
    assign P[34] = in1[3] ^ in2[3];
    assign G[35] = in1[2] & in2[2];
    assign P[35] = in1[2] ^ in2[2];
    assign G[36] = in1[1] & in2[1];
    assign P[36] = in1[1] ^ in2[1];
    assign G[37] = in1[0] & in2[0];
    assign P[37] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign cout = G[37] | (P[37] & C[37]);
    assign sum = P ^ C;
endmodule

module CLA_37(output [36:0] sum, output cout, input [36:0] in1, input [36:0] in2);

    wire[36:0] G;
    wire[36:0] C;
    wire[36:0] P;

    assign G[0] = in1[36] & in2[36];
    assign P[0] = in1[36] ^ in2[36];
    assign G[1] = in1[35] & in2[35];
    assign P[1] = in1[35] ^ in2[35];
    assign G[2] = in1[34] & in2[34];
    assign P[2] = in1[34] ^ in2[34];
    assign G[3] = in1[33] & in2[33];
    assign P[3] = in1[33] ^ in2[33];
    assign G[4] = in1[32] & in2[32];
    assign P[4] = in1[32] ^ in2[32];
    assign G[5] = in1[31] & in2[31];
    assign P[5] = in1[31] ^ in2[31];
    assign G[6] = in1[30] & in2[30];
    assign P[6] = in1[30] ^ in2[30];
    assign G[7] = in1[29] & in2[29];
    assign P[7] = in1[29] ^ in2[29];
    assign G[8] = in1[28] & in2[28];
    assign P[8] = in1[28] ^ in2[28];
    assign G[9] = in1[27] & in2[27];
    assign P[9] = in1[27] ^ in2[27];
    assign G[10] = in1[26] & in2[26];
    assign P[10] = in1[26] ^ in2[26];
    assign G[11] = in1[25] & in2[25];
    assign P[11] = in1[25] ^ in2[25];
    assign G[12] = in1[24] & in2[24];
    assign P[12] = in1[24] ^ in2[24];
    assign G[13] = in1[23] & in2[23];
    assign P[13] = in1[23] ^ in2[23];
    assign G[14] = in1[22] & in2[22];
    assign P[14] = in1[22] ^ in2[22];
    assign G[15] = in1[21] & in2[21];
    assign P[15] = in1[21] ^ in2[21];
    assign G[16] = in1[20] & in2[20];
    assign P[16] = in1[20] ^ in2[20];
    assign G[17] = in1[19] & in2[19];
    assign P[17] = in1[19] ^ in2[19];
    assign G[18] = in1[18] & in2[18];
    assign P[18] = in1[18] ^ in2[18];
    assign G[19] = in1[17] & in2[17];
    assign P[19] = in1[17] ^ in2[17];
    assign G[20] = in1[16] & in2[16];
    assign P[20] = in1[16] ^ in2[16];
    assign G[21] = in1[15] & in2[15];
    assign P[21] = in1[15] ^ in2[15];
    assign G[22] = in1[14] & in2[14];
    assign P[22] = in1[14] ^ in2[14];
    assign G[23] = in1[13] & in2[13];
    assign P[23] = in1[13] ^ in2[13];
    assign G[24] = in1[12] & in2[12];
    assign P[24] = in1[12] ^ in2[12];
    assign G[25] = in1[11] & in2[11];
    assign P[25] = in1[11] ^ in2[11];
    assign G[26] = in1[10] & in2[10];
    assign P[26] = in1[10] ^ in2[10];
    assign G[27] = in1[9] & in2[9];
    assign P[27] = in1[9] ^ in2[9];
    assign G[28] = in1[8] & in2[8];
    assign P[28] = in1[8] ^ in2[8];
    assign G[29] = in1[7] & in2[7];
    assign P[29] = in1[7] ^ in2[7];
    assign G[30] = in1[6] & in2[6];
    assign P[30] = in1[6] ^ in2[6];
    assign G[31] = in1[5] & in2[5];
    assign P[31] = in1[5] ^ in2[5];
    assign G[32] = in1[4] & in2[4];
    assign P[32] = in1[4] ^ in2[4];
    assign G[33] = in1[3] & in2[3];
    assign P[33] = in1[3] ^ in2[3];
    assign G[34] = in1[2] & in2[2];
    assign P[34] = in1[2] ^ in2[2];
    assign G[35] = in1[1] & in2[1];
    assign P[35] = in1[1] ^ in2[1];
    assign G[36] = in1[0] & in2[0];
    assign P[36] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign cout = G[36] | (P[36] & C[36]);
    assign sum = P ^ C;
endmodule

module CLA_36(output [35:0] sum, output cout, input [35:0] in1, input [35:0] in2);

    wire[35:0] G;
    wire[35:0] C;
    wire[35:0] P;

    assign G[0] = in1[35] & in2[35];
    assign P[0] = in1[35] ^ in2[35];
    assign G[1] = in1[34] & in2[34];
    assign P[1] = in1[34] ^ in2[34];
    assign G[2] = in1[33] & in2[33];
    assign P[2] = in1[33] ^ in2[33];
    assign G[3] = in1[32] & in2[32];
    assign P[3] = in1[32] ^ in2[32];
    assign G[4] = in1[31] & in2[31];
    assign P[4] = in1[31] ^ in2[31];
    assign G[5] = in1[30] & in2[30];
    assign P[5] = in1[30] ^ in2[30];
    assign G[6] = in1[29] & in2[29];
    assign P[6] = in1[29] ^ in2[29];
    assign G[7] = in1[28] & in2[28];
    assign P[7] = in1[28] ^ in2[28];
    assign G[8] = in1[27] & in2[27];
    assign P[8] = in1[27] ^ in2[27];
    assign G[9] = in1[26] & in2[26];
    assign P[9] = in1[26] ^ in2[26];
    assign G[10] = in1[25] & in2[25];
    assign P[10] = in1[25] ^ in2[25];
    assign G[11] = in1[24] & in2[24];
    assign P[11] = in1[24] ^ in2[24];
    assign G[12] = in1[23] & in2[23];
    assign P[12] = in1[23] ^ in2[23];
    assign G[13] = in1[22] & in2[22];
    assign P[13] = in1[22] ^ in2[22];
    assign G[14] = in1[21] & in2[21];
    assign P[14] = in1[21] ^ in2[21];
    assign G[15] = in1[20] & in2[20];
    assign P[15] = in1[20] ^ in2[20];
    assign G[16] = in1[19] & in2[19];
    assign P[16] = in1[19] ^ in2[19];
    assign G[17] = in1[18] & in2[18];
    assign P[17] = in1[18] ^ in2[18];
    assign G[18] = in1[17] & in2[17];
    assign P[18] = in1[17] ^ in2[17];
    assign G[19] = in1[16] & in2[16];
    assign P[19] = in1[16] ^ in2[16];
    assign G[20] = in1[15] & in2[15];
    assign P[20] = in1[15] ^ in2[15];
    assign G[21] = in1[14] & in2[14];
    assign P[21] = in1[14] ^ in2[14];
    assign G[22] = in1[13] & in2[13];
    assign P[22] = in1[13] ^ in2[13];
    assign G[23] = in1[12] & in2[12];
    assign P[23] = in1[12] ^ in2[12];
    assign G[24] = in1[11] & in2[11];
    assign P[24] = in1[11] ^ in2[11];
    assign G[25] = in1[10] & in2[10];
    assign P[25] = in1[10] ^ in2[10];
    assign G[26] = in1[9] & in2[9];
    assign P[26] = in1[9] ^ in2[9];
    assign G[27] = in1[8] & in2[8];
    assign P[27] = in1[8] ^ in2[8];
    assign G[28] = in1[7] & in2[7];
    assign P[28] = in1[7] ^ in2[7];
    assign G[29] = in1[6] & in2[6];
    assign P[29] = in1[6] ^ in2[6];
    assign G[30] = in1[5] & in2[5];
    assign P[30] = in1[5] ^ in2[5];
    assign G[31] = in1[4] & in2[4];
    assign P[31] = in1[4] ^ in2[4];
    assign G[32] = in1[3] & in2[3];
    assign P[32] = in1[3] ^ in2[3];
    assign G[33] = in1[2] & in2[2];
    assign P[33] = in1[2] ^ in2[2];
    assign G[34] = in1[1] & in2[1];
    assign P[34] = in1[1] ^ in2[1];
    assign G[35] = in1[0] & in2[0];
    assign P[35] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign cout = G[35] | (P[35] & C[35]);
    assign sum = P ^ C;
endmodule

module CLA_35(output [34:0] sum, output cout, input [34:0] in1, input [34:0] in2);

    wire[34:0] G;
    wire[34:0] C;
    wire[34:0] P;

    assign G[0] = in1[34] & in2[34];
    assign P[0] = in1[34] ^ in2[34];
    assign G[1] = in1[33] & in2[33];
    assign P[1] = in1[33] ^ in2[33];
    assign G[2] = in1[32] & in2[32];
    assign P[2] = in1[32] ^ in2[32];
    assign G[3] = in1[31] & in2[31];
    assign P[3] = in1[31] ^ in2[31];
    assign G[4] = in1[30] & in2[30];
    assign P[4] = in1[30] ^ in2[30];
    assign G[5] = in1[29] & in2[29];
    assign P[5] = in1[29] ^ in2[29];
    assign G[6] = in1[28] & in2[28];
    assign P[6] = in1[28] ^ in2[28];
    assign G[7] = in1[27] & in2[27];
    assign P[7] = in1[27] ^ in2[27];
    assign G[8] = in1[26] & in2[26];
    assign P[8] = in1[26] ^ in2[26];
    assign G[9] = in1[25] & in2[25];
    assign P[9] = in1[25] ^ in2[25];
    assign G[10] = in1[24] & in2[24];
    assign P[10] = in1[24] ^ in2[24];
    assign G[11] = in1[23] & in2[23];
    assign P[11] = in1[23] ^ in2[23];
    assign G[12] = in1[22] & in2[22];
    assign P[12] = in1[22] ^ in2[22];
    assign G[13] = in1[21] & in2[21];
    assign P[13] = in1[21] ^ in2[21];
    assign G[14] = in1[20] & in2[20];
    assign P[14] = in1[20] ^ in2[20];
    assign G[15] = in1[19] & in2[19];
    assign P[15] = in1[19] ^ in2[19];
    assign G[16] = in1[18] & in2[18];
    assign P[16] = in1[18] ^ in2[18];
    assign G[17] = in1[17] & in2[17];
    assign P[17] = in1[17] ^ in2[17];
    assign G[18] = in1[16] & in2[16];
    assign P[18] = in1[16] ^ in2[16];
    assign G[19] = in1[15] & in2[15];
    assign P[19] = in1[15] ^ in2[15];
    assign G[20] = in1[14] & in2[14];
    assign P[20] = in1[14] ^ in2[14];
    assign G[21] = in1[13] & in2[13];
    assign P[21] = in1[13] ^ in2[13];
    assign G[22] = in1[12] & in2[12];
    assign P[22] = in1[12] ^ in2[12];
    assign G[23] = in1[11] & in2[11];
    assign P[23] = in1[11] ^ in2[11];
    assign G[24] = in1[10] & in2[10];
    assign P[24] = in1[10] ^ in2[10];
    assign G[25] = in1[9] & in2[9];
    assign P[25] = in1[9] ^ in2[9];
    assign G[26] = in1[8] & in2[8];
    assign P[26] = in1[8] ^ in2[8];
    assign G[27] = in1[7] & in2[7];
    assign P[27] = in1[7] ^ in2[7];
    assign G[28] = in1[6] & in2[6];
    assign P[28] = in1[6] ^ in2[6];
    assign G[29] = in1[5] & in2[5];
    assign P[29] = in1[5] ^ in2[5];
    assign G[30] = in1[4] & in2[4];
    assign P[30] = in1[4] ^ in2[4];
    assign G[31] = in1[3] & in2[3];
    assign P[31] = in1[3] ^ in2[3];
    assign G[32] = in1[2] & in2[2];
    assign P[32] = in1[2] ^ in2[2];
    assign G[33] = in1[1] & in2[1];
    assign P[33] = in1[1] ^ in2[1];
    assign G[34] = in1[0] & in2[0];
    assign P[34] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign cout = G[34] | (P[34] & C[34]);
    assign sum = P ^ C;
endmodule

module CLA_34(output [33:0] sum, output cout, input [33:0] in1, input [33:0] in2);

    wire[33:0] G;
    wire[33:0] C;
    wire[33:0] P;

    assign G[0] = in1[33] & in2[33];
    assign P[0] = in1[33] ^ in2[33];
    assign G[1] = in1[32] & in2[32];
    assign P[1] = in1[32] ^ in2[32];
    assign G[2] = in1[31] & in2[31];
    assign P[2] = in1[31] ^ in2[31];
    assign G[3] = in1[30] & in2[30];
    assign P[3] = in1[30] ^ in2[30];
    assign G[4] = in1[29] & in2[29];
    assign P[4] = in1[29] ^ in2[29];
    assign G[5] = in1[28] & in2[28];
    assign P[5] = in1[28] ^ in2[28];
    assign G[6] = in1[27] & in2[27];
    assign P[6] = in1[27] ^ in2[27];
    assign G[7] = in1[26] & in2[26];
    assign P[7] = in1[26] ^ in2[26];
    assign G[8] = in1[25] & in2[25];
    assign P[8] = in1[25] ^ in2[25];
    assign G[9] = in1[24] & in2[24];
    assign P[9] = in1[24] ^ in2[24];
    assign G[10] = in1[23] & in2[23];
    assign P[10] = in1[23] ^ in2[23];
    assign G[11] = in1[22] & in2[22];
    assign P[11] = in1[22] ^ in2[22];
    assign G[12] = in1[21] & in2[21];
    assign P[12] = in1[21] ^ in2[21];
    assign G[13] = in1[20] & in2[20];
    assign P[13] = in1[20] ^ in2[20];
    assign G[14] = in1[19] & in2[19];
    assign P[14] = in1[19] ^ in2[19];
    assign G[15] = in1[18] & in2[18];
    assign P[15] = in1[18] ^ in2[18];
    assign G[16] = in1[17] & in2[17];
    assign P[16] = in1[17] ^ in2[17];
    assign G[17] = in1[16] & in2[16];
    assign P[17] = in1[16] ^ in2[16];
    assign G[18] = in1[15] & in2[15];
    assign P[18] = in1[15] ^ in2[15];
    assign G[19] = in1[14] & in2[14];
    assign P[19] = in1[14] ^ in2[14];
    assign G[20] = in1[13] & in2[13];
    assign P[20] = in1[13] ^ in2[13];
    assign G[21] = in1[12] & in2[12];
    assign P[21] = in1[12] ^ in2[12];
    assign G[22] = in1[11] & in2[11];
    assign P[22] = in1[11] ^ in2[11];
    assign G[23] = in1[10] & in2[10];
    assign P[23] = in1[10] ^ in2[10];
    assign G[24] = in1[9] & in2[9];
    assign P[24] = in1[9] ^ in2[9];
    assign G[25] = in1[8] & in2[8];
    assign P[25] = in1[8] ^ in2[8];
    assign G[26] = in1[7] & in2[7];
    assign P[26] = in1[7] ^ in2[7];
    assign G[27] = in1[6] & in2[6];
    assign P[27] = in1[6] ^ in2[6];
    assign G[28] = in1[5] & in2[5];
    assign P[28] = in1[5] ^ in2[5];
    assign G[29] = in1[4] & in2[4];
    assign P[29] = in1[4] ^ in2[4];
    assign G[30] = in1[3] & in2[3];
    assign P[30] = in1[3] ^ in2[3];
    assign G[31] = in1[2] & in2[2];
    assign P[31] = in1[2] ^ in2[2];
    assign G[32] = in1[1] & in2[1];
    assign P[32] = in1[1] ^ in2[1];
    assign G[33] = in1[0] & in2[0];
    assign P[33] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign cout = G[33] | (P[33] & C[33]);
    assign sum = P ^ C;
endmodule

module CLA_33(output [32:0] sum, output cout, input [32:0] in1, input [32:0] in2);

    wire[32:0] G;
    wire[32:0] C;
    wire[32:0] P;

    assign G[0] = in1[32] & in2[32];
    assign P[0] = in1[32] ^ in2[32];
    assign G[1] = in1[31] & in2[31];
    assign P[1] = in1[31] ^ in2[31];
    assign G[2] = in1[30] & in2[30];
    assign P[2] = in1[30] ^ in2[30];
    assign G[3] = in1[29] & in2[29];
    assign P[3] = in1[29] ^ in2[29];
    assign G[4] = in1[28] & in2[28];
    assign P[4] = in1[28] ^ in2[28];
    assign G[5] = in1[27] & in2[27];
    assign P[5] = in1[27] ^ in2[27];
    assign G[6] = in1[26] & in2[26];
    assign P[6] = in1[26] ^ in2[26];
    assign G[7] = in1[25] & in2[25];
    assign P[7] = in1[25] ^ in2[25];
    assign G[8] = in1[24] & in2[24];
    assign P[8] = in1[24] ^ in2[24];
    assign G[9] = in1[23] & in2[23];
    assign P[9] = in1[23] ^ in2[23];
    assign G[10] = in1[22] & in2[22];
    assign P[10] = in1[22] ^ in2[22];
    assign G[11] = in1[21] & in2[21];
    assign P[11] = in1[21] ^ in2[21];
    assign G[12] = in1[20] & in2[20];
    assign P[12] = in1[20] ^ in2[20];
    assign G[13] = in1[19] & in2[19];
    assign P[13] = in1[19] ^ in2[19];
    assign G[14] = in1[18] & in2[18];
    assign P[14] = in1[18] ^ in2[18];
    assign G[15] = in1[17] & in2[17];
    assign P[15] = in1[17] ^ in2[17];
    assign G[16] = in1[16] & in2[16];
    assign P[16] = in1[16] ^ in2[16];
    assign G[17] = in1[15] & in2[15];
    assign P[17] = in1[15] ^ in2[15];
    assign G[18] = in1[14] & in2[14];
    assign P[18] = in1[14] ^ in2[14];
    assign G[19] = in1[13] & in2[13];
    assign P[19] = in1[13] ^ in2[13];
    assign G[20] = in1[12] & in2[12];
    assign P[20] = in1[12] ^ in2[12];
    assign G[21] = in1[11] & in2[11];
    assign P[21] = in1[11] ^ in2[11];
    assign G[22] = in1[10] & in2[10];
    assign P[22] = in1[10] ^ in2[10];
    assign G[23] = in1[9] & in2[9];
    assign P[23] = in1[9] ^ in2[9];
    assign G[24] = in1[8] & in2[8];
    assign P[24] = in1[8] ^ in2[8];
    assign G[25] = in1[7] & in2[7];
    assign P[25] = in1[7] ^ in2[7];
    assign G[26] = in1[6] & in2[6];
    assign P[26] = in1[6] ^ in2[6];
    assign G[27] = in1[5] & in2[5];
    assign P[27] = in1[5] ^ in2[5];
    assign G[28] = in1[4] & in2[4];
    assign P[28] = in1[4] ^ in2[4];
    assign G[29] = in1[3] & in2[3];
    assign P[29] = in1[3] ^ in2[3];
    assign G[30] = in1[2] & in2[2];
    assign P[30] = in1[2] ^ in2[2];
    assign G[31] = in1[1] & in2[1];
    assign P[31] = in1[1] ^ in2[1];
    assign G[32] = in1[0] & in2[0];
    assign P[32] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign cout = G[32] | (P[32] & C[32]);
    assign sum = P ^ C;
endmodule

module CLA_32(output [31:0] sum, output cout, input [31:0] in1, input [31:0] in2);

    wire[31:0] G;
    wire[31:0] C;
    wire[31:0] P;

    assign G[0] = in1[31] & in2[31];
    assign P[0] = in1[31] ^ in2[31];
    assign G[1] = in1[30] & in2[30];
    assign P[1] = in1[30] ^ in2[30];
    assign G[2] = in1[29] & in2[29];
    assign P[2] = in1[29] ^ in2[29];
    assign G[3] = in1[28] & in2[28];
    assign P[3] = in1[28] ^ in2[28];
    assign G[4] = in1[27] & in2[27];
    assign P[4] = in1[27] ^ in2[27];
    assign G[5] = in1[26] & in2[26];
    assign P[5] = in1[26] ^ in2[26];
    assign G[6] = in1[25] & in2[25];
    assign P[6] = in1[25] ^ in2[25];
    assign G[7] = in1[24] & in2[24];
    assign P[7] = in1[24] ^ in2[24];
    assign G[8] = in1[23] & in2[23];
    assign P[8] = in1[23] ^ in2[23];
    assign G[9] = in1[22] & in2[22];
    assign P[9] = in1[22] ^ in2[22];
    assign G[10] = in1[21] & in2[21];
    assign P[10] = in1[21] ^ in2[21];
    assign G[11] = in1[20] & in2[20];
    assign P[11] = in1[20] ^ in2[20];
    assign G[12] = in1[19] & in2[19];
    assign P[12] = in1[19] ^ in2[19];
    assign G[13] = in1[18] & in2[18];
    assign P[13] = in1[18] ^ in2[18];
    assign G[14] = in1[17] & in2[17];
    assign P[14] = in1[17] ^ in2[17];
    assign G[15] = in1[16] & in2[16];
    assign P[15] = in1[16] ^ in2[16];
    assign G[16] = in1[15] & in2[15];
    assign P[16] = in1[15] ^ in2[15];
    assign G[17] = in1[14] & in2[14];
    assign P[17] = in1[14] ^ in2[14];
    assign G[18] = in1[13] & in2[13];
    assign P[18] = in1[13] ^ in2[13];
    assign G[19] = in1[12] & in2[12];
    assign P[19] = in1[12] ^ in2[12];
    assign G[20] = in1[11] & in2[11];
    assign P[20] = in1[11] ^ in2[11];
    assign G[21] = in1[10] & in2[10];
    assign P[21] = in1[10] ^ in2[10];
    assign G[22] = in1[9] & in2[9];
    assign P[22] = in1[9] ^ in2[9];
    assign G[23] = in1[8] & in2[8];
    assign P[23] = in1[8] ^ in2[8];
    assign G[24] = in1[7] & in2[7];
    assign P[24] = in1[7] ^ in2[7];
    assign G[25] = in1[6] & in2[6];
    assign P[25] = in1[6] ^ in2[6];
    assign G[26] = in1[5] & in2[5];
    assign P[26] = in1[5] ^ in2[5];
    assign G[27] = in1[4] & in2[4];
    assign P[27] = in1[4] ^ in2[4];
    assign G[28] = in1[3] & in2[3];
    assign P[28] = in1[3] ^ in2[3];
    assign G[29] = in1[2] & in2[2];
    assign P[29] = in1[2] ^ in2[2];
    assign G[30] = in1[1] & in2[1];
    assign P[30] = in1[1] ^ in2[1];
    assign G[31] = in1[0] & in2[0];
    assign P[31] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign cout = G[31] | (P[31] & C[31]);
    assign sum = P ^ C;
endmodule

module CLA_31(output [30:0] sum, output cout, input [30:0] in1, input [30:0] in2);

    wire[30:0] G;
    wire[30:0] C;
    wire[30:0] P;

    assign G[0] = in1[30] & in2[30];
    assign P[0] = in1[30] ^ in2[30];
    assign G[1] = in1[29] & in2[29];
    assign P[1] = in1[29] ^ in2[29];
    assign G[2] = in1[28] & in2[28];
    assign P[2] = in1[28] ^ in2[28];
    assign G[3] = in1[27] & in2[27];
    assign P[3] = in1[27] ^ in2[27];
    assign G[4] = in1[26] & in2[26];
    assign P[4] = in1[26] ^ in2[26];
    assign G[5] = in1[25] & in2[25];
    assign P[5] = in1[25] ^ in2[25];
    assign G[6] = in1[24] & in2[24];
    assign P[6] = in1[24] ^ in2[24];
    assign G[7] = in1[23] & in2[23];
    assign P[7] = in1[23] ^ in2[23];
    assign G[8] = in1[22] & in2[22];
    assign P[8] = in1[22] ^ in2[22];
    assign G[9] = in1[21] & in2[21];
    assign P[9] = in1[21] ^ in2[21];
    assign G[10] = in1[20] & in2[20];
    assign P[10] = in1[20] ^ in2[20];
    assign G[11] = in1[19] & in2[19];
    assign P[11] = in1[19] ^ in2[19];
    assign G[12] = in1[18] & in2[18];
    assign P[12] = in1[18] ^ in2[18];
    assign G[13] = in1[17] & in2[17];
    assign P[13] = in1[17] ^ in2[17];
    assign G[14] = in1[16] & in2[16];
    assign P[14] = in1[16] ^ in2[16];
    assign G[15] = in1[15] & in2[15];
    assign P[15] = in1[15] ^ in2[15];
    assign G[16] = in1[14] & in2[14];
    assign P[16] = in1[14] ^ in2[14];
    assign G[17] = in1[13] & in2[13];
    assign P[17] = in1[13] ^ in2[13];
    assign G[18] = in1[12] & in2[12];
    assign P[18] = in1[12] ^ in2[12];
    assign G[19] = in1[11] & in2[11];
    assign P[19] = in1[11] ^ in2[11];
    assign G[20] = in1[10] & in2[10];
    assign P[20] = in1[10] ^ in2[10];
    assign G[21] = in1[9] & in2[9];
    assign P[21] = in1[9] ^ in2[9];
    assign G[22] = in1[8] & in2[8];
    assign P[22] = in1[8] ^ in2[8];
    assign G[23] = in1[7] & in2[7];
    assign P[23] = in1[7] ^ in2[7];
    assign G[24] = in1[6] & in2[6];
    assign P[24] = in1[6] ^ in2[6];
    assign G[25] = in1[5] & in2[5];
    assign P[25] = in1[5] ^ in2[5];
    assign G[26] = in1[4] & in2[4];
    assign P[26] = in1[4] ^ in2[4];
    assign G[27] = in1[3] & in2[3];
    assign P[27] = in1[3] ^ in2[3];
    assign G[28] = in1[2] & in2[2];
    assign P[28] = in1[2] ^ in2[2];
    assign G[29] = in1[1] & in2[1];
    assign P[29] = in1[1] ^ in2[1];
    assign G[30] = in1[0] & in2[0];
    assign P[30] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign cout = G[30] | (P[30] & C[30]);
    assign sum = P ^ C;
endmodule

module CLA_30(output [29:0] sum, output cout, input [29:0] in1, input [29:0] in2);

    wire[29:0] G;
    wire[29:0] C;
    wire[29:0] P;

    assign G[0] = in1[29] & in2[29];
    assign P[0] = in1[29] ^ in2[29];
    assign G[1] = in1[28] & in2[28];
    assign P[1] = in1[28] ^ in2[28];
    assign G[2] = in1[27] & in2[27];
    assign P[2] = in1[27] ^ in2[27];
    assign G[3] = in1[26] & in2[26];
    assign P[3] = in1[26] ^ in2[26];
    assign G[4] = in1[25] & in2[25];
    assign P[4] = in1[25] ^ in2[25];
    assign G[5] = in1[24] & in2[24];
    assign P[5] = in1[24] ^ in2[24];
    assign G[6] = in1[23] & in2[23];
    assign P[6] = in1[23] ^ in2[23];
    assign G[7] = in1[22] & in2[22];
    assign P[7] = in1[22] ^ in2[22];
    assign G[8] = in1[21] & in2[21];
    assign P[8] = in1[21] ^ in2[21];
    assign G[9] = in1[20] & in2[20];
    assign P[9] = in1[20] ^ in2[20];
    assign G[10] = in1[19] & in2[19];
    assign P[10] = in1[19] ^ in2[19];
    assign G[11] = in1[18] & in2[18];
    assign P[11] = in1[18] ^ in2[18];
    assign G[12] = in1[17] & in2[17];
    assign P[12] = in1[17] ^ in2[17];
    assign G[13] = in1[16] & in2[16];
    assign P[13] = in1[16] ^ in2[16];
    assign G[14] = in1[15] & in2[15];
    assign P[14] = in1[15] ^ in2[15];
    assign G[15] = in1[14] & in2[14];
    assign P[15] = in1[14] ^ in2[14];
    assign G[16] = in1[13] & in2[13];
    assign P[16] = in1[13] ^ in2[13];
    assign G[17] = in1[12] & in2[12];
    assign P[17] = in1[12] ^ in2[12];
    assign G[18] = in1[11] & in2[11];
    assign P[18] = in1[11] ^ in2[11];
    assign G[19] = in1[10] & in2[10];
    assign P[19] = in1[10] ^ in2[10];
    assign G[20] = in1[9] & in2[9];
    assign P[20] = in1[9] ^ in2[9];
    assign G[21] = in1[8] & in2[8];
    assign P[21] = in1[8] ^ in2[8];
    assign G[22] = in1[7] & in2[7];
    assign P[22] = in1[7] ^ in2[7];
    assign G[23] = in1[6] & in2[6];
    assign P[23] = in1[6] ^ in2[6];
    assign G[24] = in1[5] & in2[5];
    assign P[24] = in1[5] ^ in2[5];
    assign G[25] = in1[4] & in2[4];
    assign P[25] = in1[4] ^ in2[4];
    assign G[26] = in1[3] & in2[3];
    assign P[26] = in1[3] ^ in2[3];
    assign G[27] = in1[2] & in2[2];
    assign P[27] = in1[2] ^ in2[2];
    assign G[28] = in1[1] & in2[1];
    assign P[28] = in1[1] ^ in2[1];
    assign G[29] = in1[0] & in2[0];
    assign P[29] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign cout = G[29] | (P[29] & C[29]);
    assign sum = P ^ C;
endmodule

module CLA_29(output [28:0] sum, output cout, input [28:0] in1, input [28:0] in2);

    wire[28:0] G;
    wire[28:0] C;
    wire[28:0] P;

    assign G[0] = in1[28] & in2[28];
    assign P[0] = in1[28] ^ in2[28];
    assign G[1] = in1[27] & in2[27];
    assign P[1] = in1[27] ^ in2[27];
    assign G[2] = in1[26] & in2[26];
    assign P[2] = in1[26] ^ in2[26];
    assign G[3] = in1[25] & in2[25];
    assign P[3] = in1[25] ^ in2[25];
    assign G[4] = in1[24] & in2[24];
    assign P[4] = in1[24] ^ in2[24];
    assign G[5] = in1[23] & in2[23];
    assign P[5] = in1[23] ^ in2[23];
    assign G[6] = in1[22] & in2[22];
    assign P[6] = in1[22] ^ in2[22];
    assign G[7] = in1[21] & in2[21];
    assign P[7] = in1[21] ^ in2[21];
    assign G[8] = in1[20] & in2[20];
    assign P[8] = in1[20] ^ in2[20];
    assign G[9] = in1[19] & in2[19];
    assign P[9] = in1[19] ^ in2[19];
    assign G[10] = in1[18] & in2[18];
    assign P[10] = in1[18] ^ in2[18];
    assign G[11] = in1[17] & in2[17];
    assign P[11] = in1[17] ^ in2[17];
    assign G[12] = in1[16] & in2[16];
    assign P[12] = in1[16] ^ in2[16];
    assign G[13] = in1[15] & in2[15];
    assign P[13] = in1[15] ^ in2[15];
    assign G[14] = in1[14] & in2[14];
    assign P[14] = in1[14] ^ in2[14];
    assign G[15] = in1[13] & in2[13];
    assign P[15] = in1[13] ^ in2[13];
    assign G[16] = in1[12] & in2[12];
    assign P[16] = in1[12] ^ in2[12];
    assign G[17] = in1[11] & in2[11];
    assign P[17] = in1[11] ^ in2[11];
    assign G[18] = in1[10] & in2[10];
    assign P[18] = in1[10] ^ in2[10];
    assign G[19] = in1[9] & in2[9];
    assign P[19] = in1[9] ^ in2[9];
    assign G[20] = in1[8] & in2[8];
    assign P[20] = in1[8] ^ in2[8];
    assign G[21] = in1[7] & in2[7];
    assign P[21] = in1[7] ^ in2[7];
    assign G[22] = in1[6] & in2[6];
    assign P[22] = in1[6] ^ in2[6];
    assign G[23] = in1[5] & in2[5];
    assign P[23] = in1[5] ^ in2[5];
    assign G[24] = in1[4] & in2[4];
    assign P[24] = in1[4] ^ in2[4];
    assign G[25] = in1[3] & in2[3];
    assign P[25] = in1[3] ^ in2[3];
    assign G[26] = in1[2] & in2[2];
    assign P[26] = in1[2] ^ in2[2];
    assign G[27] = in1[1] & in2[1];
    assign P[27] = in1[1] ^ in2[1];
    assign G[28] = in1[0] & in2[0];
    assign P[28] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign cout = G[28] | (P[28] & C[28]);
    assign sum = P ^ C;
endmodule

module CLA_28(output [27:0] sum, output cout, input [27:0] in1, input [27:0] in2);

    wire[27:0] G;
    wire[27:0] C;
    wire[27:0] P;

    assign G[0] = in1[27] & in2[27];
    assign P[0] = in1[27] ^ in2[27];
    assign G[1] = in1[26] & in2[26];
    assign P[1] = in1[26] ^ in2[26];
    assign G[2] = in1[25] & in2[25];
    assign P[2] = in1[25] ^ in2[25];
    assign G[3] = in1[24] & in2[24];
    assign P[3] = in1[24] ^ in2[24];
    assign G[4] = in1[23] & in2[23];
    assign P[4] = in1[23] ^ in2[23];
    assign G[5] = in1[22] & in2[22];
    assign P[5] = in1[22] ^ in2[22];
    assign G[6] = in1[21] & in2[21];
    assign P[6] = in1[21] ^ in2[21];
    assign G[7] = in1[20] & in2[20];
    assign P[7] = in1[20] ^ in2[20];
    assign G[8] = in1[19] & in2[19];
    assign P[8] = in1[19] ^ in2[19];
    assign G[9] = in1[18] & in2[18];
    assign P[9] = in1[18] ^ in2[18];
    assign G[10] = in1[17] & in2[17];
    assign P[10] = in1[17] ^ in2[17];
    assign G[11] = in1[16] & in2[16];
    assign P[11] = in1[16] ^ in2[16];
    assign G[12] = in1[15] & in2[15];
    assign P[12] = in1[15] ^ in2[15];
    assign G[13] = in1[14] & in2[14];
    assign P[13] = in1[14] ^ in2[14];
    assign G[14] = in1[13] & in2[13];
    assign P[14] = in1[13] ^ in2[13];
    assign G[15] = in1[12] & in2[12];
    assign P[15] = in1[12] ^ in2[12];
    assign G[16] = in1[11] & in2[11];
    assign P[16] = in1[11] ^ in2[11];
    assign G[17] = in1[10] & in2[10];
    assign P[17] = in1[10] ^ in2[10];
    assign G[18] = in1[9] & in2[9];
    assign P[18] = in1[9] ^ in2[9];
    assign G[19] = in1[8] & in2[8];
    assign P[19] = in1[8] ^ in2[8];
    assign G[20] = in1[7] & in2[7];
    assign P[20] = in1[7] ^ in2[7];
    assign G[21] = in1[6] & in2[6];
    assign P[21] = in1[6] ^ in2[6];
    assign G[22] = in1[5] & in2[5];
    assign P[22] = in1[5] ^ in2[5];
    assign G[23] = in1[4] & in2[4];
    assign P[23] = in1[4] ^ in2[4];
    assign G[24] = in1[3] & in2[3];
    assign P[24] = in1[3] ^ in2[3];
    assign G[25] = in1[2] & in2[2];
    assign P[25] = in1[2] ^ in2[2];
    assign G[26] = in1[1] & in2[1];
    assign P[26] = in1[1] ^ in2[1];
    assign G[27] = in1[0] & in2[0];
    assign P[27] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign cout = G[27] | (P[27] & C[27]);
    assign sum = P ^ C;
endmodule

module CLA_27(output [26:0] sum, output cout, input [26:0] in1, input [26:0] in2);

    wire[26:0] G;
    wire[26:0] C;
    wire[26:0] P;

    assign G[0] = in1[26] & in2[26];
    assign P[0] = in1[26] ^ in2[26];
    assign G[1] = in1[25] & in2[25];
    assign P[1] = in1[25] ^ in2[25];
    assign G[2] = in1[24] & in2[24];
    assign P[2] = in1[24] ^ in2[24];
    assign G[3] = in1[23] & in2[23];
    assign P[3] = in1[23] ^ in2[23];
    assign G[4] = in1[22] & in2[22];
    assign P[4] = in1[22] ^ in2[22];
    assign G[5] = in1[21] & in2[21];
    assign P[5] = in1[21] ^ in2[21];
    assign G[6] = in1[20] & in2[20];
    assign P[6] = in1[20] ^ in2[20];
    assign G[7] = in1[19] & in2[19];
    assign P[7] = in1[19] ^ in2[19];
    assign G[8] = in1[18] & in2[18];
    assign P[8] = in1[18] ^ in2[18];
    assign G[9] = in1[17] & in2[17];
    assign P[9] = in1[17] ^ in2[17];
    assign G[10] = in1[16] & in2[16];
    assign P[10] = in1[16] ^ in2[16];
    assign G[11] = in1[15] & in2[15];
    assign P[11] = in1[15] ^ in2[15];
    assign G[12] = in1[14] & in2[14];
    assign P[12] = in1[14] ^ in2[14];
    assign G[13] = in1[13] & in2[13];
    assign P[13] = in1[13] ^ in2[13];
    assign G[14] = in1[12] & in2[12];
    assign P[14] = in1[12] ^ in2[12];
    assign G[15] = in1[11] & in2[11];
    assign P[15] = in1[11] ^ in2[11];
    assign G[16] = in1[10] & in2[10];
    assign P[16] = in1[10] ^ in2[10];
    assign G[17] = in1[9] & in2[9];
    assign P[17] = in1[9] ^ in2[9];
    assign G[18] = in1[8] & in2[8];
    assign P[18] = in1[8] ^ in2[8];
    assign G[19] = in1[7] & in2[7];
    assign P[19] = in1[7] ^ in2[7];
    assign G[20] = in1[6] & in2[6];
    assign P[20] = in1[6] ^ in2[6];
    assign G[21] = in1[5] & in2[5];
    assign P[21] = in1[5] ^ in2[5];
    assign G[22] = in1[4] & in2[4];
    assign P[22] = in1[4] ^ in2[4];
    assign G[23] = in1[3] & in2[3];
    assign P[23] = in1[3] ^ in2[3];
    assign G[24] = in1[2] & in2[2];
    assign P[24] = in1[2] ^ in2[2];
    assign G[25] = in1[1] & in2[1];
    assign P[25] = in1[1] ^ in2[1];
    assign G[26] = in1[0] & in2[0];
    assign P[26] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign cout = G[26] | (P[26] & C[26]);
    assign sum = P ^ C;
endmodule

module CLA_26(output [25:0] sum, output cout, input [25:0] in1, input [25:0] in2);

    wire[25:0] G;
    wire[25:0] C;
    wire[25:0] P;

    assign G[0] = in1[25] & in2[25];
    assign P[0] = in1[25] ^ in2[25];
    assign G[1] = in1[24] & in2[24];
    assign P[1] = in1[24] ^ in2[24];
    assign G[2] = in1[23] & in2[23];
    assign P[2] = in1[23] ^ in2[23];
    assign G[3] = in1[22] & in2[22];
    assign P[3] = in1[22] ^ in2[22];
    assign G[4] = in1[21] & in2[21];
    assign P[4] = in1[21] ^ in2[21];
    assign G[5] = in1[20] & in2[20];
    assign P[5] = in1[20] ^ in2[20];
    assign G[6] = in1[19] & in2[19];
    assign P[6] = in1[19] ^ in2[19];
    assign G[7] = in1[18] & in2[18];
    assign P[7] = in1[18] ^ in2[18];
    assign G[8] = in1[17] & in2[17];
    assign P[8] = in1[17] ^ in2[17];
    assign G[9] = in1[16] & in2[16];
    assign P[9] = in1[16] ^ in2[16];
    assign G[10] = in1[15] & in2[15];
    assign P[10] = in1[15] ^ in2[15];
    assign G[11] = in1[14] & in2[14];
    assign P[11] = in1[14] ^ in2[14];
    assign G[12] = in1[13] & in2[13];
    assign P[12] = in1[13] ^ in2[13];
    assign G[13] = in1[12] & in2[12];
    assign P[13] = in1[12] ^ in2[12];
    assign G[14] = in1[11] & in2[11];
    assign P[14] = in1[11] ^ in2[11];
    assign G[15] = in1[10] & in2[10];
    assign P[15] = in1[10] ^ in2[10];
    assign G[16] = in1[9] & in2[9];
    assign P[16] = in1[9] ^ in2[9];
    assign G[17] = in1[8] & in2[8];
    assign P[17] = in1[8] ^ in2[8];
    assign G[18] = in1[7] & in2[7];
    assign P[18] = in1[7] ^ in2[7];
    assign G[19] = in1[6] & in2[6];
    assign P[19] = in1[6] ^ in2[6];
    assign G[20] = in1[5] & in2[5];
    assign P[20] = in1[5] ^ in2[5];
    assign G[21] = in1[4] & in2[4];
    assign P[21] = in1[4] ^ in2[4];
    assign G[22] = in1[3] & in2[3];
    assign P[22] = in1[3] ^ in2[3];
    assign G[23] = in1[2] & in2[2];
    assign P[23] = in1[2] ^ in2[2];
    assign G[24] = in1[1] & in2[1];
    assign P[24] = in1[1] ^ in2[1];
    assign G[25] = in1[0] & in2[0];
    assign P[25] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign cout = G[25] | (P[25] & C[25]);
    assign sum = P ^ C;
endmodule

module CLA_25(output [24:0] sum, output cout, input [24:0] in1, input [24:0] in2);

    wire[24:0] G;
    wire[24:0] C;
    wire[24:0] P;

    assign G[0] = in1[24] & in2[24];
    assign P[0] = in1[24] ^ in2[24];
    assign G[1] = in1[23] & in2[23];
    assign P[1] = in1[23] ^ in2[23];
    assign G[2] = in1[22] & in2[22];
    assign P[2] = in1[22] ^ in2[22];
    assign G[3] = in1[21] & in2[21];
    assign P[3] = in1[21] ^ in2[21];
    assign G[4] = in1[20] & in2[20];
    assign P[4] = in1[20] ^ in2[20];
    assign G[5] = in1[19] & in2[19];
    assign P[5] = in1[19] ^ in2[19];
    assign G[6] = in1[18] & in2[18];
    assign P[6] = in1[18] ^ in2[18];
    assign G[7] = in1[17] & in2[17];
    assign P[7] = in1[17] ^ in2[17];
    assign G[8] = in1[16] & in2[16];
    assign P[8] = in1[16] ^ in2[16];
    assign G[9] = in1[15] & in2[15];
    assign P[9] = in1[15] ^ in2[15];
    assign G[10] = in1[14] & in2[14];
    assign P[10] = in1[14] ^ in2[14];
    assign G[11] = in1[13] & in2[13];
    assign P[11] = in1[13] ^ in2[13];
    assign G[12] = in1[12] & in2[12];
    assign P[12] = in1[12] ^ in2[12];
    assign G[13] = in1[11] & in2[11];
    assign P[13] = in1[11] ^ in2[11];
    assign G[14] = in1[10] & in2[10];
    assign P[14] = in1[10] ^ in2[10];
    assign G[15] = in1[9] & in2[9];
    assign P[15] = in1[9] ^ in2[9];
    assign G[16] = in1[8] & in2[8];
    assign P[16] = in1[8] ^ in2[8];
    assign G[17] = in1[7] & in2[7];
    assign P[17] = in1[7] ^ in2[7];
    assign G[18] = in1[6] & in2[6];
    assign P[18] = in1[6] ^ in2[6];
    assign G[19] = in1[5] & in2[5];
    assign P[19] = in1[5] ^ in2[5];
    assign G[20] = in1[4] & in2[4];
    assign P[20] = in1[4] ^ in2[4];
    assign G[21] = in1[3] & in2[3];
    assign P[21] = in1[3] ^ in2[3];
    assign G[22] = in1[2] & in2[2];
    assign P[22] = in1[2] ^ in2[2];
    assign G[23] = in1[1] & in2[1];
    assign P[23] = in1[1] ^ in2[1];
    assign G[24] = in1[0] & in2[0];
    assign P[24] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign cout = G[24] | (P[24] & C[24]);
    assign sum = P ^ C;
endmodule

module CLA_24(output [23:0] sum, output cout, input [23:0] in1, input [23:0] in2);

    wire[23:0] G;
    wire[23:0] C;
    wire[23:0] P;

    assign G[0] = in1[23] & in2[23];
    assign P[0] = in1[23] ^ in2[23];
    assign G[1] = in1[22] & in2[22];
    assign P[1] = in1[22] ^ in2[22];
    assign G[2] = in1[21] & in2[21];
    assign P[2] = in1[21] ^ in2[21];
    assign G[3] = in1[20] & in2[20];
    assign P[3] = in1[20] ^ in2[20];
    assign G[4] = in1[19] & in2[19];
    assign P[4] = in1[19] ^ in2[19];
    assign G[5] = in1[18] & in2[18];
    assign P[5] = in1[18] ^ in2[18];
    assign G[6] = in1[17] & in2[17];
    assign P[6] = in1[17] ^ in2[17];
    assign G[7] = in1[16] & in2[16];
    assign P[7] = in1[16] ^ in2[16];
    assign G[8] = in1[15] & in2[15];
    assign P[8] = in1[15] ^ in2[15];
    assign G[9] = in1[14] & in2[14];
    assign P[9] = in1[14] ^ in2[14];
    assign G[10] = in1[13] & in2[13];
    assign P[10] = in1[13] ^ in2[13];
    assign G[11] = in1[12] & in2[12];
    assign P[11] = in1[12] ^ in2[12];
    assign G[12] = in1[11] & in2[11];
    assign P[12] = in1[11] ^ in2[11];
    assign G[13] = in1[10] & in2[10];
    assign P[13] = in1[10] ^ in2[10];
    assign G[14] = in1[9] & in2[9];
    assign P[14] = in1[9] ^ in2[9];
    assign G[15] = in1[8] & in2[8];
    assign P[15] = in1[8] ^ in2[8];
    assign G[16] = in1[7] & in2[7];
    assign P[16] = in1[7] ^ in2[7];
    assign G[17] = in1[6] & in2[6];
    assign P[17] = in1[6] ^ in2[6];
    assign G[18] = in1[5] & in2[5];
    assign P[18] = in1[5] ^ in2[5];
    assign G[19] = in1[4] & in2[4];
    assign P[19] = in1[4] ^ in2[4];
    assign G[20] = in1[3] & in2[3];
    assign P[20] = in1[3] ^ in2[3];
    assign G[21] = in1[2] & in2[2];
    assign P[21] = in1[2] ^ in2[2];
    assign G[22] = in1[1] & in2[1];
    assign P[22] = in1[1] ^ in2[1];
    assign G[23] = in1[0] & in2[0];
    assign P[23] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign cout = G[23] | (P[23] & C[23]);
    assign sum = P ^ C;
endmodule

module CLA_23(output [22:0] sum, output cout, input [22:0] in1, input [22:0] in2);

    wire[22:0] G;
    wire[22:0] C;
    wire[22:0] P;

    assign G[0] = in1[22] & in2[22];
    assign P[0] = in1[22] ^ in2[22];
    assign G[1] = in1[21] & in2[21];
    assign P[1] = in1[21] ^ in2[21];
    assign G[2] = in1[20] & in2[20];
    assign P[2] = in1[20] ^ in2[20];
    assign G[3] = in1[19] & in2[19];
    assign P[3] = in1[19] ^ in2[19];
    assign G[4] = in1[18] & in2[18];
    assign P[4] = in1[18] ^ in2[18];
    assign G[5] = in1[17] & in2[17];
    assign P[5] = in1[17] ^ in2[17];
    assign G[6] = in1[16] & in2[16];
    assign P[6] = in1[16] ^ in2[16];
    assign G[7] = in1[15] & in2[15];
    assign P[7] = in1[15] ^ in2[15];
    assign G[8] = in1[14] & in2[14];
    assign P[8] = in1[14] ^ in2[14];
    assign G[9] = in1[13] & in2[13];
    assign P[9] = in1[13] ^ in2[13];
    assign G[10] = in1[12] & in2[12];
    assign P[10] = in1[12] ^ in2[12];
    assign G[11] = in1[11] & in2[11];
    assign P[11] = in1[11] ^ in2[11];
    assign G[12] = in1[10] & in2[10];
    assign P[12] = in1[10] ^ in2[10];
    assign G[13] = in1[9] & in2[9];
    assign P[13] = in1[9] ^ in2[9];
    assign G[14] = in1[8] & in2[8];
    assign P[14] = in1[8] ^ in2[8];
    assign G[15] = in1[7] & in2[7];
    assign P[15] = in1[7] ^ in2[7];
    assign G[16] = in1[6] & in2[6];
    assign P[16] = in1[6] ^ in2[6];
    assign G[17] = in1[5] & in2[5];
    assign P[17] = in1[5] ^ in2[5];
    assign G[18] = in1[4] & in2[4];
    assign P[18] = in1[4] ^ in2[4];
    assign G[19] = in1[3] & in2[3];
    assign P[19] = in1[3] ^ in2[3];
    assign G[20] = in1[2] & in2[2];
    assign P[20] = in1[2] ^ in2[2];
    assign G[21] = in1[1] & in2[1];
    assign P[21] = in1[1] ^ in2[1];
    assign G[22] = in1[0] & in2[0];
    assign P[22] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign cout = G[22] | (P[22] & C[22]);
    assign sum = P ^ C;
endmodule

module CLA_22(output [21:0] sum, output cout, input [21:0] in1, input [21:0] in2);

    wire[21:0] G;
    wire[21:0] C;
    wire[21:0] P;

    assign G[0] = in1[21] & in2[21];
    assign P[0] = in1[21] ^ in2[21];
    assign G[1] = in1[20] & in2[20];
    assign P[1] = in1[20] ^ in2[20];
    assign G[2] = in1[19] & in2[19];
    assign P[2] = in1[19] ^ in2[19];
    assign G[3] = in1[18] & in2[18];
    assign P[3] = in1[18] ^ in2[18];
    assign G[4] = in1[17] & in2[17];
    assign P[4] = in1[17] ^ in2[17];
    assign G[5] = in1[16] & in2[16];
    assign P[5] = in1[16] ^ in2[16];
    assign G[6] = in1[15] & in2[15];
    assign P[6] = in1[15] ^ in2[15];
    assign G[7] = in1[14] & in2[14];
    assign P[7] = in1[14] ^ in2[14];
    assign G[8] = in1[13] & in2[13];
    assign P[8] = in1[13] ^ in2[13];
    assign G[9] = in1[12] & in2[12];
    assign P[9] = in1[12] ^ in2[12];
    assign G[10] = in1[11] & in2[11];
    assign P[10] = in1[11] ^ in2[11];
    assign G[11] = in1[10] & in2[10];
    assign P[11] = in1[10] ^ in2[10];
    assign G[12] = in1[9] & in2[9];
    assign P[12] = in1[9] ^ in2[9];
    assign G[13] = in1[8] & in2[8];
    assign P[13] = in1[8] ^ in2[8];
    assign G[14] = in1[7] & in2[7];
    assign P[14] = in1[7] ^ in2[7];
    assign G[15] = in1[6] & in2[6];
    assign P[15] = in1[6] ^ in2[6];
    assign G[16] = in1[5] & in2[5];
    assign P[16] = in1[5] ^ in2[5];
    assign G[17] = in1[4] & in2[4];
    assign P[17] = in1[4] ^ in2[4];
    assign G[18] = in1[3] & in2[3];
    assign P[18] = in1[3] ^ in2[3];
    assign G[19] = in1[2] & in2[2];
    assign P[19] = in1[2] ^ in2[2];
    assign G[20] = in1[1] & in2[1];
    assign P[20] = in1[1] ^ in2[1];
    assign G[21] = in1[0] & in2[0];
    assign P[21] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign cout = G[21] | (P[21] & C[21]);
    assign sum = P ^ C;
endmodule

module CLA_21(output [20:0] sum, output cout, input [20:0] in1, input [20:0] in2);

    wire[20:0] G;
    wire[20:0] C;
    wire[20:0] P;

    assign G[0] = in1[20] & in2[20];
    assign P[0] = in1[20] ^ in2[20];
    assign G[1] = in1[19] & in2[19];
    assign P[1] = in1[19] ^ in2[19];
    assign G[2] = in1[18] & in2[18];
    assign P[2] = in1[18] ^ in2[18];
    assign G[3] = in1[17] & in2[17];
    assign P[3] = in1[17] ^ in2[17];
    assign G[4] = in1[16] & in2[16];
    assign P[4] = in1[16] ^ in2[16];
    assign G[5] = in1[15] & in2[15];
    assign P[5] = in1[15] ^ in2[15];
    assign G[6] = in1[14] & in2[14];
    assign P[6] = in1[14] ^ in2[14];
    assign G[7] = in1[13] & in2[13];
    assign P[7] = in1[13] ^ in2[13];
    assign G[8] = in1[12] & in2[12];
    assign P[8] = in1[12] ^ in2[12];
    assign G[9] = in1[11] & in2[11];
    assign P[9] = in1[11] ^ in2[11];
    assign G[10] = in1[10] & in2[10];
    assign P[10] = in1[10] ^ in2[10];
    assign G[11] = in1[9] & in2[9];
    assign P[11] = in1[9] ^ in2[9];
    assign G[12] = in1[8] & in2[8];
    assign P[12] = in1[8] ^ in2[8];
    assign G[13] = in1[7] & in2[7];
    assign P[13] = in1[7] ^ in2[7];
    assign G[14] = in1[6] & in2[6];
    assign P[14] = in1[6] ^ in2[6];
    assign G[15] = in1[5] & in2[5];
    assign P[15] = in1[5] ^ in2[5];
    assign G[16] = in1[4] & in2[4];
    assign P[16] = in1[4] ^ in2[4];
    assign G[17] = in1[3] & in2[3];
    assign P[17] = in1[3] ^ in2[3];
    assign G[18] = in1[2] & in2[2];
    assign P[18] = in1[2] ^ in2[2];
    assign G[19] = in1[1] & in2[1];
    assign P[19] = in1[1] ^ in2[1];
    assign G[20] = in1[0] & in2[0];
    assign P[20] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign cout = G[20] | (P[20] & C[20]);
    assign sum = P ^ C;
endmodule

module CLA_20(output [19:0] sum, output cout, input [19:0] in1, input [19:0] in2);

    wire[19:0] G;
    wire[19:0] C;
    wire[19:0] P;

    assign G[0] = in1[19] & in2[19];
    assign P[0] = in1[19] ^ in2[19];
    assign G[1] = in1[18] & in2[18];
    assign P[1] = in1[18] ^ in2[18];
    assign G[2] = in1[17] & in2[17];
    assign P[2] = in1[17] ^ in2[17];
    assign G[3] = in1[16] & in2[16];
    assign P[3] = in1[16] ^ in2[16];
    assign G[4] = in1[15] & in2[15];
    assign P[4] = in1[15] ^ in2[15];
    assign G[5] = in1[14] & in2[14];
    assign P[5] = in1[14] ^ in2[14];
    assign G[6] = in1[13] & in2[13];
    assign P[6] = in1[13] ^ in2[13];
    assign G[7] = in1[12] & in2[12];
    assign P[7] = in1[12] ^ in2[12];
    assign G[8] = in1[11] & in2[11];
    assign P[8] = in1[11] ^ in2[11];
    assign G[9] = in1[10] & in2[10];
    assign P[9] = in1[10] ^ in2[10];
    assign G[10] = in1[9] & in2[9];
    assign P[10] = in1[9] ^ in2[9];
    assign G[11] = in1[8] & in2[8];
    assign P[11] = in1[8] ^ in2[8];
    assign G[12] = in1[7] & in2[7];
    assign P[12] = in1[7] ^ in2[7];
    assign G[13] = in1[6] & in2[6];
    assign P[13] = in1[6] ^ in2[6];
    assign G[14] = in1[5] & in2[5];
    assign P[14] = in1[5] ^ in2[5];
    assign G[15] = in1[4] & in2[4];
    assign P[15] = in1[4] ^ in2[4];
    assign G[16] = in1[3] & in2[3];
    assign P[16] = in1[3] ^ in2[3];
    assign G[17] = in1[2] & in2[2];
    assign P[17] = in1[2] ^ in2[2];
    assign G[18] = in1[1] & in2[1];
    assign P[18] = in1[1] ^ in2[1];
    assign G[19] = in1[0] & in2[0];
    assign P[19] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign cout = G[19] | (P[19] & C[19]);
    assign sum = P ^ C;
endmodule

module CLA_19(output [18:0] sum, output cout, input [18:0] in1, input [18:0] in2);

    wire[18:0] G;
    wire[18:0] C;
    wire[18:0] P;

    assign G[0] = in1[18] & in2[18];
    assign P[0] = in1[18] ^ in2[18];
    assign G[1] = in1[17] & in2[17];
    assign P[1] = in1[17] ^ in2[17];
    assign G[2] = in1[16] & in2[16];
    assign P[2] = in1[16] ^ in2[16];
    assign G[3] = in1[15] & in2[15];
    assign P[3] = in1[15] ^ in2[15];
    assign G[4] = in1[14] & in2[14];
    assign P[4] = in1[14] ^ in2[14];
    assign G[5] = in1[13] & in2[13];
    assign P[5] = in1[13] ^ in2[13];
    assign G[6] = in1[12] & in2[12];
    assign P[6] = in1[12] ^ in2[12];
    assign G[7] = in1[11] & in2[11];
    assign P[7] = in1[11] ^ in2[11];
    assign G[8] = in1[10] & in2[10];
    assign P[8] = in1[10] ^ in2[10];
    assign G[9] = in1[9] & in2[9];
    assign P[9] = in1[9] ^ in2[9];
    assign G[10] = in1[8] & in2[8];
    assign P[10] = in1[8] ^ in2[8];
    assign G[11] = in1[7] & in2[7];
    assign P[11] = in1[7] ^ in2[7];
    assign G[12] = in1[6] & in2[6];
    assign P[12] = in1[6] ^ in2[6];
    assign G[13] = in1[5] & in2[5];
    assign P[13] = in1[5] ^ in2[5];
    assign G[14] = in1[4] & in2[4];
    assign P[14] = in1[4] ^ in2[4];
    assign G[15] = in1[3] & in2[3];
    assign P[15] = in1[3] ^ in2[3];
    assign G[16] = in1[2] & in2[2];
    assign P[16] = in1[2] ^ in2[2];
    assign G[17] = in1[1] & in2[1];
    assign P[17] = in1[1] ^ in2[1];
    assign G[18] = in1[0] & in2[0];
    assign P[18] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign cout = G[18] | (P[18] & C[18]);
    assign sum = P ^ C;
endmodule

module CLA_18(output [17:0] sum, output cout, input [17:0] in1, input [17:0] in2);

    wire[17:0] G;
    wire[17:0] C;
    wire[17:0] P;

    assign G[0] = in1[17] & in2[17];
    assign P[0] = in1[17] ^ in2[17];
    assign G[1] = in1[16] & in2[16];
    assign P[1] = in1[16] ^ in2[16];
    assign G[2] = in1[15] & in2[15];
    assign P[2] = in1[15] ^ in2[15];
    assign G[3] = in1[14] & in2[14];
    assign P[3] = in1[14] ^ in2[14];
    assign G[4] = in1[13] & in2[13];
    assign P[4] = in1[13] ^ in2[13];
    assign G[5] = in1[12] & in2[12];
    assign P[5] = in1[12] ^ in2[12];
    assign G[6] = in1[11] & in2[11];
    assign P[6] = in1[11] ^ in2[11];
    assign G[7] = in1[10] & in2[10];
    assign P[7] = in1[10] ^ in2[10];
    assign G[8] = in1[9] & in2[9];
    assign P[8] = in1[9] ^ in2[9];
    assign G[9] = in1[8] & in2[8];
    assign P[9] = in1[8] ^ in2[8];
    assign G[10] = in1[7] & in2[7];
    assign P[10] = in1[7] ^ in2[7];
    assign G[11] = in1[6] & in2[6];
    assign P[11] = in1[6] ^ in2[6];
    assign G[12] = in1[5] & in2[5];
    assign P[12] = in1[5] ^ in2[5];
    assign G[13] = in1[4] & in2[4];
    assign P[13] = in1[4] ^ in2[4];
    assign G[14] = in1[3] & in2[3];
    assign P[14] = in1[3] ^ in2[3];
    assign G[15] = in1[2] & in2[2];
    assign P[15] = in1[2] ^ in2[2];
    assign G[16] = in1[1] & in2[1];
    assign P[16] = in1[1] ^ in2[1];
    assign G[17] = in1[0] & in2[0];
    assign P[17] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign cout = G[17] | (P[17] & C[17]);
    assign sum = P ^ C;
endmodule

module CLA_17(output [16:0] sum, output cout, input [16:0] in1, input [16:0] in2);

    wire[16:0] G;
    wire[16:0] C;
    wire[16:0] P;

    assign G[0] = in1[16] & in2[16];
    assign P[0] = in1[16] ^ in2[16];
    assign G[1] = in1[15] & in2[15];
    assign P[1] = in1[15] ^ in2[15];
    assign G[2] = in1[14] & in2[14];
    assign P[2] = in1[14] ^ in2[14];
    assign G[3] = in1[13] & in2[13];
    assign P[3] = in1[13] ^ in2[13];
    assign G[4] = in1[12] & in2[12];
    assign P[4] = in1[12] ^ in2[12];
    assign G[5] = in1[11] & in2[11];
    assign P[5] = in1[11] ^ in2[11];
    assign G[6] = in1[10] & in2[10];
    assign P[6] = in1[10] ^ in2[10];
    assign G[7] = in1[9] & in2[9];
    assign P[7] = in1[9] ^ in2[9];
    assign G[8] = in1[8] & in2[8];
    assign P[8] = in1[8] ^ in2[8];
    assign G[9] = in1[7] & in2[7];
    assign P[9] = in1[7] ^ in2[7];
    assign G[10] = in1[6] & in2[6];
    assign P[10] = in1[6] ^ in2[6];
    assign G[11] = in1[5] & in2[5];
    assign P[11] = in1[5] ^ in2[5];
    assign G[12] = in1[4] & in2[4];
    assign P[12] = in1[4] ^ in2[4];
    assign G[13] = in1[3] & in2[3];
    assign P[13] = in1[3] ^ in2[3];
    assign G[14] = in1[2] & in2[2];
    assign P[14] = in1[2] ^ in2[2];
    assign G[15] = in1[1] & in2[1];
    assign P[15] = in1[1] ^ in2[1];
    assign G[16] = in1[0] & in2[0];
    assign P[16] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign cout = G[16] | (P[16] & C[16]);
    assign sum = P ^ C;
endmodule

module CLA_16(output [15:0] sum, output cout, input [15:0] in1, input [15:0] in2);

    wire[15:0] G;
    wire[15:0] C;
    wire[15:0] P;

    assign G[0] = in1[15] & in2[15];
    assign P[0] = in1[15] ^ in2[15];
    assign G[1] = in1[14] & in2[14];
    assign P[1] = in1[14] ^ in2[14];
    assign G[2] = in1[13] & in2[13];
    assign P[2] = in1[13] ^ in2[13];
    assign G[3] = in1[12] & in2[12];
    assign P[3] = in1[12] ^ in2[12];
    assign G[4] = in1[11] & in2[11];
    assign P[4] = in1[11] ^ in2[11];
    assign G[5] = in1[10] & in2[10];
    assign P[5] = in1[10] ^ in2[10];
    assign G[6] = in1[9] & in2[9];
    assign P[6] = in1[9] ^ in2[9];
    assign G[7] = in1[8] & in2[8];
    assign P[7] = in1[8] ^ in2[8];
    assign G[8] = in1[7] & in2[7];
    assign P[8] = in1[7] ^ in2[7];
    assign G[9] = in1[6] & in2[6];
    assign P[9] = in1[6] ^ in2[6];
    assign G[10] = in1[5] & in2[5];
    assign P[10] = in1[5] ^ in2[5];
    assign G[11] = in1[4] & in2[4];
    assign P[11] = in1[4] ^ in2[4];
    assign G[12] = in1[3] & in2[3];
    assign P[12] = in1[3] ^ in2[3];
    assign G[13] = in1[2] & in2[2];
    assign P[13] = in1[2] ^ in2[2];
    assign G[14] = in1[1] & in2[1];
    assign P[14] = in1[1] ^ in2[1];
    assign G[15] = in1[0] & in2[0];
    assign P[15] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign cout = G[15] | (P[15] & C[15]);
    assign sum = P ^ C;
endmodule

module CLA_15(output [14:0] sum, output cout, input [14:0] in1, input [14:0] in2);

    wire[14:0] G;
    wire[14:0] C;
    wire[14:0] P;

    assign G[0] = in1[14] & in2[14];
    assign P[0] = in1[14] ^ in2[14];
    assign G[1] = in1[13] & in2[13];
    assign P[1] = in1[13] ^ in2[13];
    assign G[2] = in1[12] & in2[12];
    assign P[2] = in1[12] ^ in2[12];
    assign G[3] = in1[11] & in2[11];
    assign P[3] = in1[11] ^ in2[11];
    assign G[4] = in1[10] & in2[10];
    assign P[4] = in1[10] ^ in2[10];
    assign G[5] = in1[9] & in2[9];
    assign P[5] = in1[9] ^ in2[9];
    assign G[6] = in1[8] & in2[8];
    assign P[6] = in1[8] ^ in2[8];
    assign G[7] = in1[7] & in2[7];
    assign P[7] = in1[7] ^ in2[7];
    assign G[8] = in1[6] & in2[6];
    assign P[8] = in1[6] ^ in2[6];
    assign G[9] = in1[5] & in2[5];
    assign P[9] = in1[5] ^ in2[5];
    assign G[10] = in1[4] & in2[4];
    assign P[10] = in1[4] ^ in2[4];
    assign G[11] = in1[3] & in2[3];
    assign P[11] = in1[3] ^ in2[3];
    assign G[12] = in1[2] & in2[2];
    assign P[12] = in1[2] ^ in2[2];
    assign G[13] = in1[1] & in2[1];
    assign P[13] = in1[1] ^ in2[1];
    assign G[14] = in1[0] & in2[0];
    assign P[14] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign cout = G[14] | (P[14] & C[14]);
    assign sum = P ^ C;
endmodule

module CLA_14(output [13:0] sum, output cout, input [13:0] in1, input [13:0] in2);

    wire[13:0] G;
    wire[13:0] C;
    wire[13:0] P;

    assign G[0] = in1[13] & in2[13];
    assign P[0] = in1[13] ^ in2[13];
    assign G[1] = in1[12] & in2[12];
    assign P[1] = in1[12] ^ in2[12];
    assign G[2] = in1[11] & in2[11];
    assign P[2] = in1[11] ^ in2[11];
    assign G[3] = in1[10] & in2[10];
    assign P[3] = in1[10] ^ in2[10];
    assign G[4] = in1[9] & in2[9];
    assign P[4] = in1[9] ^ in2[9];
    assign G[5] = in1[8] & in2[8];
    assign P[5] = in1[8] ^ in2[8];
    assign G[6] = in1[7] & in2[7];
    assign P[6] = in1[7] ^ in2[7];
    assign G[7] = in1[6] & in2[6];
    assign P[7] = in1[6] ^ in2[6];
    assign G[8] = in1[5] & in2[5];
    assign P[8] = in1[5] ^ in2[5];
    assign G[9] = in1[4] & in2[4];
    assign P[9] = in1[4] ^ in2[4];
    assign G[10] = in1[3] & in2[3];
    assign P[10] = in1[3] ^ in2[3];
    assign G[11] = in1[2] & in2[2];
    assign P[11] = in1[2] ^ in2[2];
    assign G[12] = in1[1] & in2[1];
    assign P[12] = in1[1] ^ in2[1];
    assign G[13] = in1[0] & in2[0];
    assign P[13] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign cout = G[13] | (P[13] & C[13]);
    assign sum = P ^ C;
endmodule

module CLA_13(output [12:0] sum, output cout, input [12:0] in1, input [12:0] in2);

    wire[12:0] G;
    wire[12:0] C;
    wire[12:0] P;

    assign G[0] = in1[12] & in2[12];
    assign P[0] = in1[12] ^ in2[12];
    assign G[1] = in1[11] & in2[11];
    assign P[1] = in1[11] ^ in2[11];
    assign G[2] = in1[10] & in2[10];
    assign P[2] = in1[10] ^ in2[10];
    assign G[3] = in1[9] & in2[9];
    assign P[3] = in1[9] ^ in2[9];
    assign G[4] = in1[8] & in2[8];
    assign P[4] = in1[8] ^ in2[8];
    assign G[5] = in1[7] & in2[7];
    assign P[5] = in1[7] ^ in2[7];
    assign G[6] = in1[6] & in2[6];
    assign P[6] = in1[6] ^ in2[6];
    assign G[7] = in1[5] & in2[5];
    assign P[7] = in1[5] ^ in2[5];
    assign G[8] = in1[4] & in2[4];
    assign P[8] = in1[4] ^ in2[4];
    assign G[9] = in1[3] & in2[3];
    assign P[9] = in1[3] ^ in2[3];
    assign G[10] = in1[2] & in2[2];
    assign P[10] = in1[2] ^ in2[2];
    assign G[11] = in1[1] & in2[1];
    assign P[11] = in1[1] ^ in2[1];
    assign G[12] = in1[0] & in2[0];
    assign P[12] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign cout = G[12] | (P[12] & C[12]);
    assign sum = P ^ C;
endmodule

module CLA_12(output [11:0] sum, output cout, input [11:0] in1, input [11:0] in2);

    wire[11:0] G;
    wire[11:0] C;
    wire[11:0] P;

    assign G[0] = in1[11] & in2[11];
    assign P[0] = in1[11] ^ in2[11];
    assign G[1] = in1[10] & in2[10];
    assign P[1] = in1[10] ^ in2[10];
    assign G[2] = in1[9] & in2[9];
    assign P[2] = in1[9] ^ in2[9];
    assign G[3] = in1[8] & in2[8];
    assign P[3] = in1[8] ^ in2[8];
    assign G[4] = in1[7] & in2[7];
    assign P[4] = in1[7] ^ in2[7];
    assign G[5] = in1[6] & in2[6];
    assign P[5] = in1[6] ^ in2[6];
    assign G[6] = in1[5] & in2[5];
    assign P[6] = in1[5] ^ in2[5];
    assign G[7] = in1[4] & in2[4];
    assign P[7] = in1[4] ^ in2[4];
    assign G[8] = in1[3] & in2[3];
    assign P[8] = in1[3] ^ in2[3];
    assign G[9] = in1[2] & in2[2];
    assign P[9] = in1[2] ^ in2[2];
    assign G[10] = in1[1] & in2[1];
    assign P[10] = in1[1] ^ in2[1];
    assign G[11] = in1[0] & in2[0];
    assign P[11] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign cout = G[11] | (P[11] & C[11]);
    assign sum = P ^ C;
endmodule

module CLA_11(output [10:0] sum, output cout, input [10:0] in1, input [10:0] in2);

    wire[10:0] G;
    wire[10:0] C;
    wire[10:0] P;

    assign G[0] = in1[10] & in2[10];
    assign P[0] = in1[10] ^ in2[10];
    assign G[1] = in1[9] & in2[9];
    assign P[1] = in1[9] ^ in2[9];
    assign G[2] = in1[8] & in2[8];
    assign P[2] = in1[8] ^ in2[8];
    assign G[3] = in1[7] & in2[7];
    assign P[3] = in1[7] ^ in2[7];
    assign G[4] = in1[6] & in2[6];
    assign P[4] = in1[6] ^ in2[6];
    assign G[5] = in1[5] & in2[5];
    assign P[5] = in1[5] ^ in2[5];
    assign G[6] = in1[4] & in2[4];
    assign P[6] = in1[4] ^ in2[4];
    assign G[7] = in1[3] & in2[3];
    assign P[7] = in1[3] ^ in2[3];
    assign G[8] = in1[2] & in2[2];
    assign P[8] = in1[2] ^ in2[2];
    assign G[9] = in1[1] & in2[1];
    assign P[9] = in1[1] ^ in2[1];
    assign G[10] = in1[0] & in2[0];
    assign P[10] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign cout = G[10] | (P[10] & C[10]);
    assign sum = P ^ C;
endmodule

module CLA_10(output [9:0] sum, output cout, input [9:0] in1, input [9:0] in2);

    wire[9:0] G;
    wire[9:0] C;
    wire[9:0] P;

    assign G[0] = in1[9] & in2[9];
    assign P[0] = in1[9] ^ in2[9];
    assign G[1] = in1[8] & in2[8];
    assign P[1] = in1[8] ^ in2[8];
    assign G[2] = in1[7] & in2[7];
    assign P[2] = in1[7] ^ in2[7];
    assign G[3] = in1[6] & in2[6];
    assign P[3] = in1[6] ^ in2[6];
    assign G[4] = in1[5] & in2[5];
    assign P[4] = in1[5] ^ in2[5];
    assign G[5] = in1[4] & in2[4];
    assign P[5] = in1[4] ^ in2[4];
    assign G[6] = in1[3] & in2[3];
    assign P[6] = in1[3] ^ in2[3];
    assign G[7] = in1[2] & in2[2];
    assign P[7] = in1[2] ^ in2[2];
    assign G[8] = in1[1] & in2[1];
    assign P[8] = in1[1] ^ in2[1];
    assign G[9] = in1[0] & in2[0];
    assign P[9] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign cout = G[9] | (P[9] & C[9]);
    assign sum = P ^ C;
endmodule

module CLA_9(output [8:0] sum, output cout, input [8:0] in1, input [8:0] in2);

    wire[8:0] G;
    wire[8:0] C;
    wire[8:0] P;

    assign G[0] = in1[8] & in2[8];
    assign P[0] = in1[8] ^ in2[8];
    assign G[1] = in1[7] & in2[7];
    assign P[1] = in1[7] ^ in2[7];
    assign G[2] = in1[6] & in2[6];
    assign P[2] = in1[6] ^ in2[6];
    assign G[3] = in1[5] & in2[5];
    assign P[3] = in1[5] ^ in2[5];
    assign G[4] = in1[4] & in2[4];
    assign P[4] = in1[4] ^ in2[4];
    assign G[5] = in1[3] & in2[3];
    assign P[5] = in1[3] ^ in2[3];
    assign G[6] = in1[2] & in2[2];
    assign P[6] = in1[2] ^ in2[2];
    assign G[7] = in1[1] & in2[1];
    assign P[7] = in1[1] ^ in2[1];
    assign G[8] = in1[0] & in2[0];
    assign P[8] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign cout = G[8] | (P[8] & C[8]);
    assign sum = P ^ C;
endmodule

module CLA_8(output [7:0] sum, output cout, input [7:0] in1, input [7:0] in2);

    wire[7:0] G;
    wire[7:0] C;
    wire[7:0] P;

    assign G[0] = in1[7] & in2[7];
    assign P[0] = in1[7] ^ in2[7];
    assign G[1] = in1[6] & in2[6];
    assign P[1] = in1[6] ^ in2[6];
    assign G[2] = in1[5] & in2[5];
    assign P[2] = in1[5] ^ in2[5];
    assign G[3] = in1[4] & in2[4];
    assign P[3] = in1[4] ^ in2[4];
    assign G[4] = in1[3] & in2[3];
    assign P[4] = in1[3] ^ in2[3];
    assign G[5] = in1[2] & in2[2];
    assign P[5] = in1[2] ^ in2[2];
    assign G[6] = in1[1] & in2[1];
    assign P[6] = in1[1] ^ in2[1];
    assign G[7] = in1[0] & in2[0];
    assign P[7] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign cout = G[7] | (P[7] & C[7]);
    assign sum = P ^ C;
endmodule

module CLA_7(output [6:0] sum, output cout, input [6:0] in1, input [6:0] in2);

    wire[6:0] G;
    wire[6:0] C;
    wire[6:0] P;

    assign G[0] = in1[6] & in2[6];
    assign P[0] = in1[6] ^ in2[6];
    assign G[1] = in1[5] & in2[5];
    assign P[1] = in1[5] ^ in2[5];
    assign G[2] = in1[4] & in2[4];
    assign P[2] = in1[4] ^ in2[4];
    assign G[3] = in1[3] & in2[3];
    assign P[3] = in1[3] ^ in2[3];
    assign G[4] = in1[2] & in2[2];
    assign P[4] = in1[2] ^ in2[2];
    assign G[5] = in1[1] & in2[1];
    assign P[5] = in1[1] ^ in2[1];
    assign G[6] = in1[0] & in2[0];
    assign P[6] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign cout = G[6] | (P[6] & C[6]);
    assign sum = P ^ C;
endmodule

module CLA_6(output [5:0] sum, output cout, input [5:0] in1, input [5:0] in2);

    wire[5:0] G;
    wire[5:0] C;
    wire[5:0] P;

    assign G[0] = in1[5] & in2[5];
    assign P[0] = in1[5] ^ in2[5];
    assign G[1] = in1[4] & in2[4];
    assign P[1] = in1[4] ^ in2[4];
    assign G[2] = in1[3] & in2[3];
    assign P[2] = in1[3] ^ in2[3];
    assign G[3] = in1[2] & in2[2];
    assign P[3] = in1[2] ^ in2[2];
    assign G[4] = in1[1] & in2[1];
    assign P[4] = in1[1] ^ in2[1];
    assign G[5] = in1[0] & in2[0];
    assign P[5] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign cout = G[5] | (P[5] & C[5]);
    assign sum = P ^ C;
endmodule

module CLA_5(output [4:0] sum, output cout, input [4:0] in1, input [4:0] in2);

    wire[4:0] G;
    wire[4:0] C;
    wire[4:0] P;

    assign G[0] = in1[4] & in2[4];
    assign P[0] = in1[4] ^ in2[4];
    assign G[1] = in1[3] & in2[3];
    assign P[1] = in1[3] ^ in2[3];
    assign G[2] = in1[2] & in2[2];
    assign P[2] = in1[2] ^ in2[2];
    assign G[3] = in1[1] & in2[1];
    assign P[3] = in1[1] ^ in2[1];
    assign G[4] = in1[0] & in2[0];
    assign P[4] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign cout = G[4] | (P[4] & C[4]);
    assign sum = P ^ C;
endmodule

module CLA_4(output [3:0] sum, output cout, input [3:0] in1, input [3:0] in2);

    wire[3:0] G;
    wire[3:0] C;
    wire[3:0] P;

    assign G[0] = in1[3] & in2[3];
    assign P[0] = in1[3] ^ in2[3];
    assign G[1] = in1[2] & in2[2];
    assign P[1] = in1[2] ^ in2[2];
    assign G[2] = in1[1] & in2[1];
    assign P[2] = in1[1] ^ in2[1];
    assign G[3] = in1[0] & in2[0];
    assign P[3] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign cout = G[3] | (P[3] & C[3]);
    assign sum = P ^ C;
endmodule

module CLA_3(output [2:0] sum, output cout, input [2:0] in1, input [2:0] in2);

    wire[2:0] G;
    wire[2:0] C;
    wire[2:0] P;

    assign G[0] = in1[2] & in2[2];
    assign P[0] = in1[2] ^ in2[2];
    assign G[1] = in1[1] & in2[1];
    assign P[1] = in1[1] ^ in2[1];
    assign G[2] = in1[0] & in2[0];
    assign P[2] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign cout = G[2] | (P[2] & C[2]);
    assign sum = P ^ C;
endmodule

module CLA_2(output [1:0] sum, output cout, input [1:0] in1, input [1:0] in2);

    wire[1:0] G;
    wire[1:0] C;
    wire[1:0] P;

    assign G[0] = in1[1] & in2[1];
    assign P[0] = in1[1] ^ in2[1];
    assign G[1] = in1[0] & in2[0];
    assign P[1] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign cout = G[1] | (P[1] & C[1]);
    assign sum = P ^ C;
endmodule



module Half_Adder(input wire in1,
                  input wire in2,
		  output wire sum,
                  output wire cout);
    xor(sum, in1, in2);
    and(cout, in1, in2);
endmodule

module Full_Adder(input wire in1,
                  input wire in2,
                  input wire cin,
		  output wire sum,
                  output wire cout);
    wire temp1;
    wire temp2;
    wire temp3;
    xor(sum, in1, in2, cin);
    and(temp1,in1,in2);
    and(temp2,in1,cin);
    and(temp3,in2,cin);
    or(cout,temp1,temp2,temp3);
endmodule
