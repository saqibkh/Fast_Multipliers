module multiplier_128bits_version14(product, A, B);

    output [255:0] product;
    input [127:0] A, B;

    /*
     * Area: 319161.534633
     * Power: 295.4140mW
     * Timing: 16.59ns
     */

    wire [127:0] pp0;
    wire [127:0] pp1;
    wire [127:0] pp2;
    wire [127:0] pp3;
    wire [127:0] pp4;
    wire [127:0] pp5;
    wire [127:0] pp6;
    wire [127:0] pp7;
    wire [127:0] pp8;
    wire [127:0] pp9;
    wire [127:0] pp10;
    wire [127:0] pp11;
    wire [127:0] pp12;
    wire [127:0] pp13;
    wire [127:0] pp14;
    wire [127:0] pp15;
    wire [127:0] pp16;
    wire [127:0] pp17;
    wire [127:0] pp18;
    wire [127:0] pp19;
    wire [127:0] pp20;
    wire [127:0] pp21;
    wire [127:0] pp22;
    wire [127:0] pp23;
    wire [127:0] pp24;
    wire [127:0] pp25;
    wire [127:0] pp26;
    wire [127:0] pp27;
    wire [127:0] pp28;
    wire [127:0] pp29;
    wire [127:0] pp30;
    wire [127:0] pp31;
    wire [127:0] pp32;
    wire [127:0] pp33;
    wire [127:0] pp34;
    wire [127:0] pp35;
    wire [127:0] pp36;
    wire [127:0] pp37;
    wire [127:0] pp38;
    wire [127:0] pp39;
    wire [127:0] pp40;
    wire [127:0] pp41;
    wire [127:0] pp42;
    wire [127:0] pp43;
    wire [127:0] pp44;
    wire [127:0] pp45;
    wire [127:0] pp46;
    wire [127:0] pp47;
    wire [127:0] pp48;
    wire [127:0] pp49;
    wire [127:0] pp50;
    wire [127:0] pp51;
    wire [127:0] pp52;
    wire [127:0] pp53;
    wire [127:0] pp54;
    wire [127:0] pp55;
    wire [127:0] pp56;
    wire [127:0] pp57;
    wire [127:0] pp58;
    wire [127:0] pp59;
    wire [127:0] pp60;
    wire [127:0] pp61;
    wire [127:0] pp62;
    wire [127:0] pp63;
    wire [127:0] pp64;
    wire [127:0] pp65;
    wire [127:0] pp66;
    wire [127:0] pp67;
    wire [127:0] pp68;
    wire [127:0] pp69;
    wire [127:0] pp70;
    wire [127:0] pp71;
    wire [127:0] pp72;
    wire [127:0] pp73;
    wire [127:0] pp74;
    wire [127:0] pp75;
    wire [127:0] pp76;
    wire [127:0] pp77;
    wire [127:0] pp78;
    wire [127:0] pp79;
    wire [127:0] pp80;
    wire [127:0] pp81;
    wire [127:0] pp82;
    wire [127:0] pp83;
    wire [127:0] pp84;
    wire [127:0] pp85;
    wire [127:0] pp86;
    wire [127:0] pp87;
    wire [127:0] pp88;
    wire [127:0] pp89;
    wire [127:0] pp90;
    wire [127:0] pp91;
    wire [127:0] pp92;
    wire [127:0] pp93;
    wire [127:0] pp94;
    wire [127:0] pp95;
    wire [127:0] pp96;
    wire [127:0] pp97;
    wire [127:0] pp98;
    wire [127:0] pp99;
    wire [127:0] pp100;
    wire [127:0] pp101;
    wire [127:0] pp102;
    wire [127:0] pp103;
    wire [127:0] pp104;
    wire [127:0] pp105;
    wire [127:0] pp106;
    wire [127:0] pp107;
    wire [127:0] pp108;
    wire [127:0] pp109;
    wire [127:0] pp110;
    wire [127:0] pp111;
    wire [127:0] pp112;
    wire [127:0] pp113;
    wire [127:0] pp114;
    wire [127:0] pp115;
    wire [127:0] pp116;
    wire [127:0] pp117;
    wire [127:0] pp118;
    wire [127:0] pp119;
    wire [127:0] pp120;
    wire [127:0] pp121;
    wire [127:0] pp122;
    wire [127:0] pp123;
    wire [127:0] pp124;
    wire [127:0] pp125;
    wire [127:0] pp126;
    wire [127:0] pp127;


    assign pp0 = A[0] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp1 = A[1] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp2 = A[2] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp3 = A[3] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp4 = A[4] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp5 = A[5] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp6 = A[6] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp7 = A[7] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp8 = A[8] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp9 = A[9] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp10 = A[10] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp11 = A[11] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp12 = A[12] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp13 = A[13] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp14 = A[14] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp15 = A[15] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp16 = A[16] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp17 = A[17] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp18 = A[18] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp19 = A[19] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp20 = A[20] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp21 = A[21] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp22 = A[22] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp23 = A[23] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp24 = A[24] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp25 = A[25] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp26 = A[26] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp27 = A[27] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp28 = A[28] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp29 = A[29] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp30 = A[30] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp31 = A[31] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp32 = A[32] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp33 = A[33] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp34 = A[34] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp35 = A[35] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp36 = A[36] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp37 = A[37] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp38 = A[38] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp39 = A[39] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp40 = A[40] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp41 = A[41] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp42 = A[42] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp43 = A[43] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp44 = A[44] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp45 = A[45] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp46 = A[46] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp47 = A[47] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp48 = A[48] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp49 = A[49] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp50 = A[50] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp51 = A[51] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp52 = A[52] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp53 = A[53] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp54 = A[54] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp55 = A[55] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp56 = A[56] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp57 = A[57] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp58 = A[58] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp59 = A[59] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp60 = A[60] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp61 = A[61] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp62 = A[62] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp63 = A[63] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp64 = A[64] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp65 = A[65] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp66 = A[66] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp67 = A[67] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp68 = A[68] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp69 = A[69] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp70 = A[70] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp71 = A[71] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp72 = A[72] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp73 = A[73] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp74 = A[74] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp75 = A[75] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp76 = A[76] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp77 = A[77] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp78 = A[78] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp79 = A[79] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp80 = A[80] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp81 = A[81] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp82 = A[82] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp83 = A[83] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp84 = A[84] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp85 = A[85] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp86 = A[86] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp87 = A[87] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp88 = A[88] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp89 = A[89] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp90 = A[90] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp91 = A[91] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp92 = A[92] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp93 = A[93] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp94 = A[94] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp95 = A[95] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp96 = A[96] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp97 = A[97] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp98 = A[98] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp99 = A[99] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp100 = A[100] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp101 = A[101] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp102 = A[102] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp103 = A[103] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp104 = A[104] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp105 = A[105] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp106 = A[106] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp107 = A[107] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp108 = A[108] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp109 = A[109] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp110 = A[110] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp111 = A[111] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp112 = A[112] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp113 = A[113] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp114 = A[114] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp115 = A[115] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp116 = A[116] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp117 = A[117] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp118 = A[118] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp119 = A[119] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp120 = A[120] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp121 = A[121] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp122 = A[122] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp123 = A[123] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp124 = A[124] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp125 = A[125] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp126 = A[126] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp127 = A[127] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


    /*Stage 1*/
    wire[0:0] s1, in1_1, in1_2;
    wire c1;
    assign in1_1 = {pp0[86]};
    assign in1_2 = {pp1[85]};
    Half_Adder HA_1(s1, c1, in1_1, in1_2);
    wire[0:0] s2, in2_1, in2_2;
    wire c2;
    assign in2_1 = {pp1[86]};
    assign in2_2 = {pp2[85]};
    Full_Adder FA_2(s2, c2, in2_1, in2_2, pp0[87]);
    wire[0:0] s3, in3_1, in3_2;
    wire c3;
    assign in3_1 = {pp3[84]};
    assign in3_2 = {pp4[83]};
    Half_Adder HA_3(s3, c3, in3_1, in3_2);
    wire[0:0] s4, in4_1, in4_2;
    wire c4;
    assign in4_1 = {pp1[87]};
    assign in4_2 = {pp2[86]};
    Full_Adder FA_4(s4, c4, in4_1, in4_2, pp0[88]);
    wire[0:0] s5, in5_1, in5_2;
    wire c5;
    assign in5_1 = {pp4[84]};
    assign in5_2 = {pp5[83]};
    Full_Adder FA_5(s5, c5, in5_1, in5_2, pp3[85]);
    wire[0:0] s6, in6_1, in6_2;
    wire c6;
    assign in6_1 = {pp6[82]};
    assign in6_2 = {pp7[81]};
    Half_Adder HA_6(s6, c6, in6_1, in6_2);
    wire[0:0] s7, in7_1, in7_2;
    wire c7;
    assign in7_1 = {pp1[88]};
    assign in7_2 = {pp2[87]};
    Full_Adder FA_7(s7, c7, in7_1, in7_2, pp0[89]);
    wire[0:0] s8, in8_1, in8_2;
    wire c8;
    assign in8_1 = {pp4[85]};
    assign in8_2 = {pp5[84]};
    Full_Adder FA_8(s8, c8, in8_1, in8_2, pp3[86]);
    wire[0:0] s9, in9_1, in9_2;
    wire c9;
    assign in9_1 = {pp7[82]};
    assign in9_2 = {pp8[81]};
    Full_Adder FA_9(s9, c9, in9_1, in9_2, pp6[83]);
    wire[0:0] s10, in10_1, in10_2;
    wire c10;
    assign in10_1 = {pp9[80]};
    assign in10_2 = {pp10[79]};
    Half_Adder HA_10(s10, c10, in10_1, in10_2);
    wire[0:0] s11, in11_1, in11_2;
    wire c11;
    assign in11_1 = {pp1[89]};
    assign in11_2 = {pp2[88]};
    Full_Adder FA_11(s11, c11, in11_1, in11_2, pp0[90]);
    wire[0:0] s12, in12_1, in12_2;
    wire c12;
    assign in12_1 = {pp4[86]};
    assign in12_2 = {pp5[85]};
    Full_Adder FA_12(s12, c12, in12_1, in12_2, pp3[87]);
    wire[0:0] s13, in13_1, in13_2;
    wire c13;
    assign in13_1 = {pp7[83]};
    assign in13_2 = {pp8[82]};
    Full_Adder FA_13(s13, c13, in13_1, in13_2, pp6[84]);
    wire[0:0] s14, in14_1, in14_2;
    wire c14;
    assign in14_1 = {pp10[80]};
    assign in14_2 = {pp11[79]};
    Full_Adder FA_14(s14, c14, in14_1, in14_2, pp9[81]);
    wire[0:0] s15, in15_1, in15_2;
    wire c15;
    assign in15_1 = {pp12[78]};
    assign in15_2 = {pp13[77]};
    Half_Adder HA_15(s15, c15, in15_1, in15_2);
    wire[0:0] s16, in16_1, in16_2;
    wire c16;
    assign in16_1 = {pp1[90]};
    assign in16_2 = {pp2[89]};
    Full_Adder FA_16(s16, c16, in16_1, in16_2, pp0[91]);
    wire[0:0] s17, in17_1, in17_2;
    wire c17;
    assign in17_1 = {pp4[87]};
    assign in17_2 = {pp5[86]};
    Full_Adder FA_17(s17, c17, in17_1, in17_2, pp3[88]);
    wire[0:0] s18, in18_1, in18_2;
    wire c18;
    assign in18_1 = {pp7[84]};
    assign in18_2 = {pp8[83]};
    Full_Adder FA_18(s18, c18, in18_1, in18_2, pp6[85]);
    wire[0:0] s19, in19_1, in19_2;
    wire c19;
    assign in19_1 = {pp10[81]};
    assign in19_2 = {pp11[80]};
    Full_Adder FA_19(s19, c19, in19_1, in19_2, pp9[82]);
    wire[0:0] s20, in20_1, in20_2;
    wire c20;
    assign in20_1 = {pp13[78]};
    assign in20_2 = {pp14[77]};
    Full_Adder FA_20(s20, c20, in20_1, in20_2, pp12[79]);
    wire[0:0] s21, in21_1, in21_2;
    wire c21;
    assign in21_1 = {pp15[76]};
    assign in21_2 = {pp16[75]};
    Half_Adder HA_21(s21, c21, in21_1, in21_2);
    wire[0:0] s22, in22_1, in22_2;
    wire c22;
    assign in22_1 = {pp1[91]};
    assign in22_2 = {pp2[90]};
    Full_Adder FA_22(s22, c22, in22_1, in22_2, pp0[92]);
    wire[0:0] s23, in23_1, in23_2;
    wire c23;
    assign in23_1 = {pp4[88]};
    assign in23_2 = {pp5[87]};
    Full_Adder FA_23(s23, c23, in23_1, in23_2, pp3[89]);
    wire[0:0] s24, in24_1, in24_2;
    wire c24;
    assign in24_1 = {pp7[85]};
    assign in24_2 = {pp8[84]};
    Full_Adder FA_24(s24, c24, in24_1, in24_2, pp6[86]);
    wire[0:0] s25, in25_1, in25_2;
    wire c25;
    assign in25_1 = {pp10[82]};
    assign in25_2 = {pp11[81]};
    Full_Adder FA_25(s25, c25, in25_1, in25_2, pp9[83]);
    wire[0:0] s26, in26_1, in26_2;
    wire c26;
    assign in26_1 = {pp13[79]};
    assign in26_2 = {pp14[78]};
    Full_Adder FA_26(s26, c26, in26_1, in26_2, pp12[80]);
    wire[0:0] s27, in27_1, in27_2;
    wire c27;
    assign in27_1 = {pp16[76]};
    assign in27_2 = {pp17[75]};
    Full_Adder FA_27(s27, c27, in27_1, in27_2, pp15[77]);
    wire[0:0] s28, in28_1, in28_2;
    wire c28;
    assign in28_1 = {pp18[74]};
    assign in28_2 = {pp19[73]};
    Half_Adder HA_28(s28, c28, in28_1, in28_2);
    wire[0:0] s29, in29_1, in29_2;
    wire c29;
    assign in29_1 = {pp1[92]};
    assign in29_2 = {pp2[91]};
    Full_Adder FA_29(s29, c29, in29_1, in29_2, pp0[93]);
    wire[0:0] s30, in30_1, in30_2;
    wire c30;
    assign in30_1 = {pp4[89]};
    assign in30_2 = {pp5[88]};
    Full_Adder FA_30(s30, c30, in30_1, in30_2, pp3[90]);
    wire[0:0] s31, in31_1, in31_2;
    wire c31;
    assign in31_1 = {pp7[86]};
    assign in31_2 = {pp8[85]};
    Full_Adder FA_31(s31, c31, in31_1, in31_2, pp6[87]);
    wire[0:0] s32, in32_1, in32_2;
    wire c32;
    assign in32_1 = {pp10[83]};
    assign in32_2 = {pp11[82]};
    Full_Adder FA_32(s32, c32, in32_1, in32_2, pp9[84]);
    wire[0:0] s33, in33_1, in33_2;
    wire c33;
    assign in33_1 = {pp13[80]};
    assign in33_2 = {pp14[79]};
    Full_Adder FA_33(s33, c33, in33_1, in33_2, pp12[81]);
    wire[0:0] s34, in34_1, in34_2;
    wire c34;
    assign in34_1 = {pp16[77]};
    assign in34_2 = {pp17[76]};
    Full_Adder FA_34(s34, c34, in34_1, in34_2, pp15[78]);
    wire[0:0] s35, in35_1, in35_2;
    wire c35;
    assign in35_1 = {pp19[74]};
    assign in35_2 = {pp20[73]};
    Full_Adder FA_35(s35, c35, in35_1, in35_2, pp18[75]);
    wire[0:0] s36, in36_1, in36_2;
    wire c36;
    assign in36_1 = {pp21[72]};
    assign in36_2 = {pp22[71]};
    Half_Adder HA_36(s36, c36, in36_1, in36_2);
    wire[0:0] s37, in37_1, in37_2;
    wire c37;
    assign in37_1 = {pp1[93]};
    assign in37_2 = {pp2[92]};
    Full_Adder FA_37(s37, c37, in37_1, in37_2, pp0[94]);
    wire[0:0] s38, in38_1, in38_2;
    wire c38;
    assign in38_1 = {pp4[90]};
    assign in38_2 = {pp5[89]};
    Full_Adder FA_38(s38, c38, in38_1, in38_2, pp3[91]);
    wire[0:0] s39, in39_1, in39_2;
    wire c39;
    assign in39_1 = {pp7[87]};
    assign in39_2 = {pp8[86]};
    Full_Adder FA_39(s39, c39, in39_1, in39_2, pp6[88]);
    wire[0:0] s40, in40_1, in40_2;
    wire c40;
    assign in40_1 = {pp10[84]};
    assign in40_2 = {pp11[83]};
    Full_Adder FA_40(s40, c40, in40_1, in40_2, pp9[85]);
    wire[0:0] s41, in41_1, in41_2;
    wire c41;
    assign in41_1 = {pp13[81]};
    assign in41_2 = {pp14[80]};
    Full_Adder FA_41(s41, c41, in41_1, in41_2, pp12[82]);
    wire[0:0] s42, in42_1, in42_2;
    wire c42;
    assign in42_1 = {pp16[78]};
    assign in42_2 = {pp17[77]};
    Full_Adder FA_42(s42, c42, in42_1, in42_2, pp15[79]);
    wire[0:0] s43, in43_1, in43_2;
    wire c43;
    assign in43_1 = {pp19[75]};
    assign in43_2 = {pp20[74]};
    Full_Adder FA_43(s43, c43, in43_1, in43_2, pp18[76]);
    wire[0:0] s44, in44_1, in44_2;
    wire c44;
    assign in44_1 = {pp22[72]};
    assign in44_2 = {pp23[71]};
    Full_Adder FA_44(s44, c44, in44_1, in44_2, pp21[73]);
    wire[0:0] s45, in45_1, in45_2;
    wire c45;
    assign in45_1 = {pp24[70]};
    assign in45_2 = {pp25[69]};
    Half_Adder HA_45(s45, c45, in45_1, in45_2);
    wire[0:0] s46, in46_1, in46_2;
    wire c46;
    assign in46_1 = {pp1[94]};
    assign in46_2 = {pp2[93]};
    Full_Adder FA_46(s46, c46, in46_1, in46_2, pp0[95]);
    wire[0:0] s47, in47_1, in47_2;
    wire c47;
    assign in47_1 = {pp4[91]};
    assign in47_2 = {pp5[90]};
    Full_Adder FA_47(s47, c47, in47_1, in47_2, pp3[92]);
    wire[0:0] s48, in48_1, in48_2;
    wire c48;
    assign in48_1 = {pp7[88]};
    assign in48_2 = {pp8[87]};
    Full_Adder FA_48(s48, c48, in48_1, in48_2, pp6[89]);
    wire[0:0] s49, in49_1, in49_2;
    wire c49;
    assign in49_1 = {pp10[85]};
    assign in49_2 = {pp11[84]};
    Full_Adder FA_49(s49, c49, in49_1, in49_2, pp9[86]);
    wire[0:0] s50, in50_1, in50_2;
    wire c50;
    assign in50_1 = {pp13[82]};
    assign in50_2 = {pp14[81]};
    Full_Adder FA_50(s50, c50, in50_1, in50_2, pp12[83]);
    wire[0:0] s51, in51_1, in51_2;
    wire c51;
    assign in51_1 = {pp16[79]};
    assign in51_2 = {pp17[78]};
    Full_Adder FA_51(s51, c51, in51_1, in51_2, pp15[80]);
    wire[0:0] s52, in52_1, in52_2;
    wire c52;
    assign in52_1 = {pp19[76]};
    assign in52_2 = {pp20[75]};
    Full_Adder FA_52(s52, c52, in52_1, in52_2, pp18[77]);
    wire[0:0] s53, in53_1, in53_2;
    wire c53;
    assign in53_1 = {pp22[73]};
    assign in53_2 = {pp23[72]};
    Full_Adder FA_53(s53, c53, in53_1, in53_2, pp21[74]);
    wire[0:0] s54, in54_1, in54_2;
    wire c54;
    assign in54_1 = {pp25[70]};
    assign in54_2 = {pp26[69]};
    Full_Adder FA_54(s54, c54, in54_1, in54_2, pp24[71]);
    wire[0:0] s55, in55_1, in55_2;
    wire c55;
    assign in55_1 = {pp27[68]};
    assign in55_2 = {pp28[67]};
    Half_Adder HA_55(s55, c55, in55_1, in55_2);
    wire[0:0] s56, in56_1, in56_2;
    wire c56;
    assign in56_1 = {pp1[95]};
    assign in56_2 = {pp2[94]};
    Full_Adder FA_56(s56, c56, in56_1, in56_2, pp0[96]);
    wire[0:0] s57, in57_1, in57_2;
    wire c57;
    assign in57_1 = {pp4[92]};
    assign in57_2 = {pp5[91]};
    Full_Adder FA_57(s57, c57, in57_1, in57_2, pp3[93]);
    wire[0:0] s58, in58_1, in58_2;
    wire c58;
    assign in58_1 = {pp7[89]};
    assign in58_2 = {pp8[88]};
    Full_Adder FA_58(s58, c58, in58_1, in58_2, pp6[90]);
    wire[0:0] s59, in59_1, in59_2;
    wire c59;
    assign in59_1 = {pp10[86]};
    assign in59_2 = {pp11[85]};
    Full_Adder FA_59(s59, c59, in59_1, in59_2, pp9[87]);
    wire[0:0] s60, in60_1, in60_2;
    wire c60;
    assign in60_1 = {pp13[83]};
    assign in60_2 = {pp14[82]};
    Full_Adder FA_60(s60, c60, in60_1, in60_2, pp12[84]);
    wire[0:0] s61, in61_1, in61_2;
    wire c61;
    assign in61_1 = {pp16[80]};
    assign in61_2 = {pp17[79]};
    Full_Adder FA_61(s61, c61, in61_1, in61_2, pp15[81]);
    wire[0:0] s62, in62_1, in62_2;
    wire c62;
    assign in62_1 = {pp19[77]};
    assign in62_2 = {pp20[76]};
    Full_Adder FA_62(s62, c62, in62_1, in62_2, pp18[78]);
    wire[0:0] s63, in63_1, in63_2;
    wire c63;
    assign in63_1 = {pp22[74]};
    assign in63_2 = {pp23[73]};
    Full_Adder FA_63(s63, c63, in63_1, in63_2, pp21[75]);
    wire[0:0] s64, in64_1, in64_2;
    wire c64;
    assign in64_1 = {pp25[71]};
    assign in64_2 = {pp26[70]};
    Full_Adder FA_64(s64, c64, in64_1, in64_2, pp24[72]);
    wire[0:0] s65, in65_1, in65_2;
    wire c65;
    assign in65_1 = {pp28[68]};
    assign in65_2 = {pp29[67]};
    Full_Adder FA_65(s65, c65, in65_1, in65_2, pp27[69]);
    wire[0:0] s66, in66_1, in66_2;
    wire c66;
    assign in66_1 = {pp30[66]};
    assign in66_2 = {pp31[65]};
    Half_Adder HA_66(s66, c66, in66_1, in66_2);
    wire[0:0] s67, in67_1, in67_2;
    wire c67;
    assign in67_1 = {pp1[96]};
    assign in67_2 = {pp2[95]};
    Full_Adder FA_67(s67, c67, in67_1, in67_2, pp0[97]);
    wire[0:0] s68, in68_1, in68_2;
    wire c68;
    assign in68_1 = {pp4[93]};
    assign in68_2 = {pp5[92]};
    Full_Adder FA_68(s68, c68, in68_1, in68_2, pp3[94]);
    wire[0:0] s69, in69_1, in69_2;
    wire c69;
    assign in69_1 = {pp7[90]};
    assign in69_2 = {pp8[89]};
    Full_Adder FA_69(s69, c69, in69_1, in69_2, pp6[91]);
    wire[0:0] s70, in70_1, in70_2;
    wire c70;
    assign in70_1 = {pp10[87]};
    assign in70_2 = {pp11[86]};
    Full_Adder FA_70(s70, c70, in70_1, in70_2, pp9[88]);
    wire[0:0] s71, in71_1, in71_2;
    wire c71;
    assign in71_1 = {pp13[84]};
    assign in71_2 = {pp14[83]};
    Full_Adder FA_71(s71, c71, in71_1, in71_2, pp12[85]);
    wire[0:0] s72, in72_1, in72_2;
    wire c72;
    assign in72_1 = {pp16[81]};
    assign in72_2 = {pp17[80]};
    Full_Adder FA_72(s72, c72, in72_1, in72_2, pp15[82]);
    wire[0:0] s73, in73_1, in73_2;
    wire c73;
    assign in73_1 = {pp19[78]};
    assign in73_2 = {pp20[77]};
    Full_Adder FA_73(s73, c73, in73_1, in73_2, pp18[79]);
    wire[0:0] s74, in74_1, in74_2;
    wire c74;
    assign in74_1 = {pp22[75]};
    assign in74_2 = {pp23[74]};
    Full_Adder FA_74(s74, c74, in74_1, in74_2, pp21[76]);
    wire[0:0] s75, in75_1, in75_2;
    wire c75;
    assign in75_1 = {pp25[72]};
    assign in75_2 = {pp26[71]};
    Full_Adder FA_75(s75, c75, in75_1, in75_2, pp24[73]);
    wire[0:0] s76, in76_1, in76_2;
    wire c76;
    assign in76_1 = {pp28[69]};
    assign in76_2 = {pp29[68]};
    Full_Adder FA_76(s76, c76, in76_1, in76_2, pp27[70]);
    wire[0:0] s77, in77_1, in77_2;
    wire c77;
    assign in77_1 = {pp31[66]};
    assign in77_2 = {pp32[65]};
    Full_Adder FA_77(s77, c77, in77_1, in77_2, pp30[67]);
    wire[0:0] s78, in78_1, in78_2;
    wire c78;
    assign in78_1 = {pp33[64]};
    assign in78_2 = {pp34[63]};
    Half_Adder HA_78(s78, c78, in78_1, in78_2);
    wire[0:0] s79, in79_1, in79_2;
    wire c79;
    assign in79_1 = {pp1[97]};
    assign in79_2 = {pp2[96]};
    Full_Adder FA_79(s79, c79, in79_1, in79_2, pp0[98]);
    wire[0:0] s80, in80_1, in80_2;
    wire c80;
    assign in80_1 = {pp4[94]};
    assign in80_2 = {pp5[93]};
    Full_Adder FA_80(s80, c80, in80_1, in80_2, pp3[95]);
    wire[0:0] s81, in81_1, in81_2;
    wire c81;
    assign in81_1 = {pp7[91]};
    assign in81_2 = {pp8[90]};
    Full_Adder FA_81(s81, c81, in81_1, in81_2, pp6[92]);
    wire[0:0] s82, in82_1, in82_2;
    wire c82;
    assign in82_1 = {pp10[88]};
    assign in82_2 = {pp11[87]};
    Full_Adder FA_82(s82, c82, in82_1, in82_2, pp9[89]);
    wire[0:0] s83, in83_1, in83_2;
    wire c83;
    assign in83_1 = {pp13[85]};
    assign in83_2 = {pp14[84]};
    Full_Adder FA_83(s83, c83, in83_1, in83_2, pp12[86]);
    wire[0:0] s84, in84_1, in84_2;
    wire c84;
    assign in84_1 = {pp16[82]};
    assign in84_2 = {pp17[81]};
    Full_Adder FA_84(s84, c84, in84_1, in84_2, pp15[83]);
    wire[0:0] s85, in85_1, in85_2;
    wire c85;
    assign in85_1 = {pp19[79]};
    assign in85_2 = {pp20[78]};
    Full_Adder FA_85(s85, c85, in85_1, in85_2, pp18[80]);
    wire[0:0] s86, in86_1, in86_2;
    wire c86;
    assign in86_1 = {pp22[76]};
    assign in86_2 = {pp23[75]};
    Full_Adder FA_86(s86, c86, in86_1, in86_2, pp21[77]);
    wire[0:0] s87, in87_1, in87_2;
    wire c87;
    assign in87_1 = {pp25[73]};
    assign in87_2 = {pp26[72]};
    Full_Adder FA_87(s87, c87, in87_1, in87_2, pp24[74]);
    wire[0:0] s88, in88_1, in88_2;
    wire c88;
    assign in88_1 = {pp28[70]};
    assign in88_2 = {pp29[69]};
    Full_Adder FA_88(s88, c88, in88_1, in88_2, pp27[71]);
    wire[0:0] s89, in89_1, in89_2;
    wire c89;
    assign in89_1 = {pp31[67]};
    assign in89_2 = {pp32[66]};
    Full_Adder FA_89(s89, c89, in89_1, in89_2, pp30[68]);
    wire[0:0] s90, in90_1, in90_2;
    wire c90;
    assign in90_1 = {pp34[64]};
    assign in90_2 = {pp35[63]};
    Full_Adder FA_90(s90, c90, in90_1, in90_2, pp33[65]);
    wire[0:0] s91, in91_1, in91_2;
    wire c91;
    assign in91_1 = {pp36[62]};
    assign in91_2 = {pp37[61]};
    Half_Adder HA_91(s91, c91, in91_1, in91_2);
    wire[0:0] s92, in92_1, in92_2;
    wire c92;
    assign in92_1 = {pp1[98]};
    assign in92_2 = {pp2[97]};
    Full_Adder FA_92(s92, c92, in92_1, in92_2, pp0[99]);
    wire[0:0] s93, in93_1, in93_2;
    wire c93;
    assign in93_1 = {pp4[95]};
    assign in93_2 = {pp5[94]};
    Full_Adder FA_93(s93, c93, in93_1, in93_2, pp3[96]);
    wire[0:0] s94, in94_1, in94_2;
    wire c94;
    assign in94_1 = {pp7[92]};
    assign in94_2 = {pp8[91]};
    Full_Adder FA_94(s94, c94, in94_1, in94_2, pp6[93]);
    wire[0:0] s95, in95_1, in95_2;
    wire c95;
    assign in95_1 = {pp10[89]};
    assign in95_2 = {pp11[88]};
    Full_Adder FA_95(s95, c95, in95_1, in95_2, pp9[90]);
    wire[0:0] s96, in96_1, in96_2;
    wire c96;
    assign in96_1 = {pp13[86]};
    assign in96_2 = {pp14[85]};
    Full_Adder FA_96(s96, c96, in96_1, in96_2, pp12[87]);
    wire[0:0] s97, in97_1, in97_2;
    wire c97;
    assign in97_1 = {pp16[83]};
    assign in97_2 = {pp17[82]};
    Full_Adder FA_97(s97, c97, in97_1, in97_2, pp15[84]);
    wire[0:0] s98, in98_1, in98_2;
    wire c98;
    assign in98_1 = {pp19[80]};
    assign in98_2 = {pp20[79]};
    Full_Adder FA_98(s98, c98, in98_1, in98_2, pp18[81]);
    wire[0:0] s99, in99_1, in99_2;
    wire c99;
    assign in99_1 = {pp22[77]};
    assign in99_2 = {pp23[76]};
    Full_Adder FA_99(s99, c99, in99_1, in99_2, pp21[78]);
    wire[0:0] s100, in100_1, in100_2;
    wire c100;
    assign in100_1 = {pp25[74]};
    assign in100_2 = {pp26[73]};
    Full_Adder FA_100(s100, c100, in100_1, in100_2, pp24[75]);
    wire[0:0] s101, in101_1, in101_2;
    wire c101;
    assign in101_1 = {pp28[71]};
    assign in101_2 = {pp29[70]};
    Full_Adder FA_101(s101, c101, in101_1, in101_2, pp27[72]);
    wire[0:0] s102, in102_1, in102_2;
    wire c102;
    assign in102_1 = {pp31[68]};
    assign in102_2 = {pp32[67]};
    Full_Adder FA_102(s102, c102, in102_1, in102_2, pp30[69]);
    wire[0:0] s103, in103_1, in103_2;
    wire c103;
    assign in103_1 = {pp34[65]};
    assign in103_2 = {pp35[64]};
    Full_Adder FA_103(s103, c103, in103_1, in103_2, pp33[66]);
    wire[0:0] s104, in104_1, in104_2;
    wire c104;
    assign in104_1 = {pp37[62]};
    assign in104_2 = {pp38[61]};
    Full_Adder FA_104(s104, c104, in104_1, in104_2, pp36[63]);
    wire[0:0] s105, in105_1, in105_2;
    wire c105;
    assign in105_1 = {pp39[60]};
    assign in105_2 = {pp40[59]};
    Half_Adder HA_105(s105, c105, in105_1, in105_2);
    wire[0:0] s106, in106_1, in106_2;
    wire c106;
    assign in106_1 = {pp1[99]};
    assign in106_2 = {pp2[98]};
    Full_Adder FA_106(s106, c106, in106_1, in106_2, pp0[100]);
    wire[0:0] s107, in107_1, in107_2;
    wire c107;
    assign in107_1 = {pp4[96]};
    assign in107_2 = {pp5[95]};
    Full_Adder FA_107(s107, c107, in107_1, in107_2, pp3[97]);
    wire[0:0] s108, in108_1, in108_2;
    wire c108;
    assign in108_1 = {pp7[93]};
    assign in108_2 = {pp8[92]};
    Full_Adder FA_108(s108, c108, in108_1, in108_2, pp6[94]);
    wire[0:0] s109, in109_1, in109_2;
    wire c109;
    assign in109_1 = {pp10[90]};
    assign in109_2 = {pp11[89]};
    Full_Adder FA_109(s109, c109, in109_1, in109_2, pp9[91]);
    wire[0:0] s110, in110_1, in110_2;
    wire c110;
    assign in110_1 = {pp13[87]};
    assign in110_2 = {pp14[86]};
    Full_Adder FA_110(s110, c110, in110_1, in110_2, pp12[88]);
    wire[0:0] s111, in111_1, in111_2;
    wire c111;
    assign in111_1 = {pp16[84]};
    assign in111_2 = {pp17[83]};
    Full_Adder FA_111(s111, c111, in111_1, in111_2, pp15[85]);
    wire[0:0] s112, in112_1, in112_2;
    wire c112;
    assign in112_1 = {pp19[81]};
    assign in112_2 = {pp20[80]};
    Full_Adder FA_112(s112, c112, in112_1, in112_2, pp18[82]);
    wire[0:0] s113, in113_1, in113_2;
    wire c113;
    assign in113_1 = {pp22[78]};
    assign in113_2 = {pp23[77]};
    Full_Adder FA_113(s113, c113, in113_1, in113_2, pp21[79]);
    wire[0:0] s114, in114_1, in114_2;
    wire c114;
    assign in114_1 = {pp25[75]};
    assign in114_2 = {pp26[74]};
    Full_Adder FA_114(s114, c114, in114_1, in114_2, pp24[76]);
    wire[0:0] s115, in115_1, in115_2;
    wire c115;
    assign in115_1 = {pp28[72]};
    assign in115_2 = {pp29[71]};
    Full_Adder FA_115(s115, c115, in115_1, in115_2, pp27[73]);
    wire[0:0] s116, in116_1, in116_2;
    wire c116;
    assign in116_1 = {pp31[69]};
    assign in116_2 = {pp32[68]};
    Full_Adder FA_116(s116, c116, in116_1, in116_2, pp30[70]);
    wire[0:0] s117, in117_1, in117_2;
    wire c117;
    assign in117_1 = {pp34[66]};
    assign in117_2 = {pp35[65]};
    Full_Adder FA_117(s117, c117, in117_1, in117_2, pp33[67]);
    wire[0:0] s118, in118_1, in118_2;
    wire c118;
    assign in118_1 = {pp37[63]};
    assign in118_2 = {pp38[62]};
    Full_Adder FA_118(s118, c118, in118_1, in118_2, pp36[64]);
    wire[0:0] s119, in119_1, in119_2;
    wire c119;
    assign in119_1 = {pp40[60]};
    assign in119_2 = {pp41[59]};
    Full_Adder FA_119(s119, c119, in119_1, in119_2, pp39[61]);
    wire[0:0] s120, in120_1, in120_2;
    wire c120;
    assign in120_1 = {pp42[58]};
    assign in120_2 = {pp43[57]};
    Half_Adder HA_120(s120, c120, in120_1, in120_2);
    wire[0:0] s121, in121_1, in121_2;
    wire c121;
    assign in121_1 = {pp1[100]};
    assign in121_2 = {pp2[99]};
    Full_Adder FA_121(s121, c121, in121_1, in121_2, pp0[101]);
    wire[0:0] s122, in122_1, in122_2;
    wire c122;
    assign in122_1 = {pp4[97]};
    assign in122_2 = {pp5[96]};
    Full_Adder FA_122(s122, c122, in122_1, in122_2, pp3[98]);
    wire[0:0] s123, in123_1, in123_2;
    wire c123;
    assign in123_1 = {pp7[94]};
    assign in123_2 = {pp8[93]};
    Full_Adder FA_123(s123, c123, in123_1, in123_2, pp6[95]);
    wire[0:0] s124, in124_1, in124_2;
    wire c124;
    assign in124_1 = {pp10[91]};
    assign in124_2 = {pp11[90]};
    Full_Adder FA_124(s124, c124, in124_1, in124_2, pp9[92]);
    wire[0:0] s125, in125_1, in125_2;
    wire c125;
    assign in125_1 = {pp13[88]};
    assign in125_2 = {pp14[87]};
    Full_Adder FA_125(s125, c125, in125_1, in125_2, pp12[89]);
    wire[0:0] s126, in126_1, in126_2;
    wire c126;
    assign in126_1 = {pp16[85]};
    assign in126_2 = {pp17[84]};
    Full_Adder FA_126(s126, c126, in126_1, in126_2, pp15[86]);
    wire[0:0] s127, in127_1, in127_2;
    wire c127;
    assign in127_1 = {pp19[82]};
    assign in127_2 = {pp20[81]};
    Full_Adder FA_127(s127, c127, in127_1, in127_2, pp18[83]);
    wire[0:0] s128, in128_1, in128_2;
    wire c128;
    assign in128_1 = {pp22[79]};
    assign in128_2 = {pp23[78]};
    Full_Adder FA_128(s128, c128, in128_1, in128_2, pp21[80]);
    wire[0:0] s129, in129_1, in129_2;
    wire c129;
    assign in129_1 = {pp25[76]};
    assign in129_2 = {pp26[75]};
    Full_Adder FA_129(s129, c129, in129_1, in129_2, pp24[77]);
    wire[0:0] s130, in130_1, in130_2;
    wire c130;
    assign in130_1 = {pp28[73]};
    assign in130_2 = {pp29[72]};
    Full_Adder FA_130(s130, c130, in130_1, in130_2, pp27[74]);
    wire[0:0] s131, in131_1, in131_2;
    wire c131;
    assign in131_1 = {pp31[70]};
    assign in131_2 = {pp32[69]};
    Full_Adder FA_131(s131, c131, in131_1, in131_2, pp30[71]);
    wire[0:0] s132, in132_1, in132_2;
    wire c132;
    assign in132_1 = {pp34[67]};
    assign in132_2 = {pp35[66]};
    Full_Adder FA_132(s132, c132, in132_1, in132_2, pp33[68]);
    wire[0:0] s133, in133_1, in133_2;
    wire c133;
    assign in133_1 = {pp37[64]};
    assign in133_2 = {pp38[63]};
    Full_Adder FA_133(s133, c133, in133_1, in133_2, pp36[65]);
    wire[0:0] s134, in134_1, in134_2;
    wire c134;
    assign in134_1 = {pp40[61]};
    assign in134_2 = {pp41[60]};
    Full_Adder FA_134(s134, c134, in134_1, in134_2, pp39[62]);
    wire[0:0] s135, in135_1, in135_2;
    wire c135;
    assign in135_1 = {pp43[58]};
    assign in135_2 = {pp44[57]};
    Full_Adder FA_135(s135, c135, in135_1, in135_2, pp42[59]);
    wire[0:0] s136, in136_1, in136_2;
    wire c136;
    assign in136_1 = {pp45[56]};
    assign in136_2 = {pp46[55]};
    Half_Adder HA_136(s136, c136, in136_1, in136_2);
    wire[0:0] s137, in137_1, in137_2;
    wire c137;
    assign in137_1 = {pp1[101]};
    assign in137_2 = {pp2[100]};
    Full_Adder FA_137(s137, c137, in137_1, in137_2, pp0[102]);
    wire[0:0] s138, in138_1, in138_2;
    wire c138;
    assign in138_1 = {pp4[98]};
    assign in138_2 = {pp5[97]};
    Full_Adder FA_138(s138, c138, in138_1, in138_2, pp3[99]);
    wire[0:0] s139, in139_1, in139_2;
    wire c139;
    assign in139_1 = {pp7[95]};
    assign in139_2 = {pp8[94]};
    Full_Adder FA_139(s139, c139, in139_1, in139_2, pp6[96]);
    wire[0:0] s140, in140_1, in140_2;
    wire c140;
    assign in140_1 = {pp10[92]};
    assign in140_2 = {pp11[91]};
    Full_Adder FA_140(s140, c140, in140_1, in140_2, pp9[93]);
    wire[0:0] s141, in141_1, in141_2;
    wire c141;
    assign in141_1 = {pp13[89]};
    assign in141_2 = {pp14[88]};
    Full_Adder FA_141(s141, c141, in141_1, in141_2, pp12[90]);
    wire[0:0] s142, in142_1, in142_2;
    wire c142;
    assign in142_1 = {pp16[86]};
    assign in142_2 = {pp17[85]};
    Full_Adder FA_142(s142, c142, in142_1, in142_2, pp15[87]);
    wire[0:0] s143, in143_1, in143_2;
    wire c143;
    assign in143_1 = {pp19[83]};
    assign in143_2 = {pp20[82]};
    Full_Adder FA_143(s143, c143, in143_1, in143_2, pp18[84]);
    wire[0:0] s144, in144_1, in144_2;
    wire c144;
    assign in144_1 = {pp22[80]};
    assign in144_2 = {pp23[79]};
    Full_Adder FA_144(s144, c144, in144_1, in144_2, pp21[81]);
    wire[0:0] s145, in145_1, in145_2;
    wire c145;
    assign in145_1 = {pp25[77]};
    assign in145_2 = {pp26[76]};
    Full_Adder FA_145(s145, c145, in145_1, in145_2, pp24[78]);
    wire[0:0] s146, in146_1, in146_2;
    wire c146;
    assign in146_1 = {pp28[74]};
    assign in146_2 = {pp29[73]};
    Full_Adder FA_146(s146, c146, in146_1, in146_2, pp27[75]);
    wire[0:0] s147, in147_1, in147_2;
    wire c147;
    assign in147_1 = {pp31[71]};
    assign in147_2 = {pp32[70]};
    Full_Adder FA_147(s147, c147, in147_1, in147_2, pp30[72]);
    wire[0:0] s148, in148_1, in148_2;
    wire c148;
    assign in148_1 = {pp34[68]};
    assign in148_2 = {pp35[67]};
    Full_Adder FA_148(s148, c148, in148_1, in148_2, pp33[69]);
    wire[0:0] s149, in149_1, in149_2;
    wire c149;
    assign in149_1 = {pp37[65]};
    assign in149_2 = {pp38[64]};
    Full_Adder FA_149(s149, c149, in149_1, in149_2, pp36[66]);
    wire[0:0] s150, in150_1, in150_2;
    wire c150;
    assign in150_1 = {pp40[62]};
    assign in150_2 = {pp41[61]};
    Full_Adder FA_150(s150, c150, in150_1, in150_2, pp39[63]);
    wire[0:0] s151, in151_1, in151_2;
    wire c151;
    assign in151_1 = {pp43[59]};
    assign in151_2 = {pp44[58]};
    Full_Adder FA_151(s151, c151, in151_1, in151_2, pp42[60]);
    wire[0:0] s152, in152_1, in152_2;
    wire c152;
    assign in152_1 = {pp46[56]};
    assign in152_2 = {pp47[55]};
    Full_Adder FA_152(s152, c152, in152_1, in152_2, pp45[57]);
    wire[0:0] s153, in153_1, in153_2;
    wire c153;
    assign in153_1 = {pp48[54]};
    assign in153_2 = {pp49[53]};
    Half_Adder HA_153(s153, c153, in153_1, in153_2);
    wire[0:0] s154, in154_1, in154_2;
    wire c154;
    assign in154_1 = {pp1[102]};
    assign in154_2 = {pp2[101]};
    Full_Adder FA_154(s154, c154, in154_1, in154_2, pp0[103]);
    wire[0:0] s155, in155_1, in155_2;
    wire c155;
    assign in155_1 = {pp4[99]};
    assign in155_2 = {pp5[98]};
    Full_Adder FA_155(s155, c155, in155_1, in155_2, pp3[100]);
    wire[0:0] s156, in156_1, in156_2;
    wire c156;
    assign in156_1 = {pp7[96]};
    assign in156_2 = {pp8[95]};
    Full_Adder FA_156(s156, c156, in156_1, in156_2, pp6[97]);
    wire[0:0] s157, in157_1, in157_2;
    wire c157;
    assign in157_1 = {pp10[93]};
    assign in157_2 = {pp11[92]};
    Full_Adder FA_157(s157, c157, in157_1, in157_2, pp9[94]);
    wire[0:0] s158, in158_1, in158_2;
    wire c158;
    assign in158_1 = {pp13[90]};
    assign in158_2 = {pp14[89]};
    Full_Adder FA_158(s158, c158, in158_1, in158_2, pp12[91]);
    wire[0:0] s159, in159_1, in159_2;
    wire c159;
    assign in159_1 = {pp16[87]};
    assign in159_2 = {pp17[86]};
    Full_Adder FA_159(s159, c159, in159_1, in159_2, pp15[88]);
    wire[0:0] s160, in160_1, in160_2;
    wire c160;
    assign in160_1 = {pp19[84]};
    assign in160_2 = {pp20[83]};
    Full_Adder FA_160(s160, c160, in160_1, in160_2, pp18[85]);
    wire[0:0] s161, in161_1, in161_2;
    wire c161;
    assign in161_1 = {pp22[81]};
    assign in161_2 = {pp23[80]};
    Full_Adder FA_161(s161, c161, in161_1, in161_2, pp21[82]);
    wire[0:0] s162, in162_1, in162_2;
    wire c162;
    assign in162_1 = {pp25[78]};
    assign in162_2 = {pp26[77]};
    Full_Adder FA_162(s162, c162, in162_1, in162_2, pp24[79]);
    wire[0:0] s163, in163_1, in163_2;
    wire c163;
    assign in163_1 = {pp28[75]};
    assign in163_2 = {pp29[74]};
    Full_Adder FA_163(s163, c163, in163_1, in163_2, pp27[76]);
    wire[0:0] s164, in164_1, in164_2;
    wire c164;
    assign in164_1 = {pp31[72]};
    assign in164_2 = {pp32[71]};
    Full_Adder FA_164(s164, c164, in164_1, in164_2, pp30[73]);
    wire[0:0] s165, in165_1, in165_2;
    wire c165;
    assign in165_1 = {pp34[69]};
    assign in165_2 = {pp35[68]};
    Full_Adder FA_165(s165, c165, in165_1, in165_2, pp33[70]);
    wire[0:0] s166, in166_1, in166_2;
    wire c166;
    assign in166_1 = {pp37[66]};
    assign in166_2 = {pp38[65]};
    Full_Adder FA_166(s166, c166, in166_1, in166_2, pp36[67]);
    wire[0:0] s167, in167_1, in167_2;
    wire c167;
    assign in167_1 = {pp40[63]};
    assign in167_2 = {pp41[62]};
    Full_Adder FA_167(s167, c167, in167_1, in167_2, pp39[64]);
    wire[0:0] s168, in168_1, in168_2;
    wire c168;
    assign in168_1 = {pp43[60]};
    assign in168_2 = {pp44[59]};
    Full_Adder FA_168(s168, c168, in168_1, in168_2, pp42[61]);
    wire[0:0] s169, in169_1, in169_2;
    wire c169;
    assign in169_1 = {pp46[57]};
    assign in169_2 = {pp47[56]};
    Full_Adder FA_169(s169, c169, in169_1, in169_2, pp45[58]);
    wire[0:0] s170, in170_1, in170_2;
    wire c170;
    assign in170_1 = {pp49[54]};
    assign in170_2 = {pp50[53]};
    Full_Adder FA_170(s170, c170, in170_1, in170_2, pp48[55]);
    wire[0:0] s171, in171_1, in171_2;
    wire c171;
    assign in171_1 = {pp51[52]};
    assign in171_2 = {pp52[51]};
    Half_Adder HA_171(s171, c171, in171_1, in171_2);
    wire[0:0] s172, in172_1, in172_2;
    wire c172;
    assign in172_1 = {pp1[103]};
    assign in172_2 = {pp2[102]};
    Full_Adder FA_172(s172, c172, in172_1, in172_2, pp0[104]);
    wire[0:0] s173, in173_1, in173_2;
    wire c173;
    assign in173_1 = {pp4[100]};
    assign in173_2 = {pp5[99]};
    Full_Adder FA_173(s173, c173, in173_1, in173_2, pp3[101]);
    wire[0:0] s174, in174_1, in174_2;
    wire c174;
    assign in174_1 = {pp7[97]};
    assign in174_2 = {pp8[96]};
    Full_Adder FA_174(s174, c174, in174_1, in174_2, pp6[98]);
    wire[0:0] s175, in175_1, in175_2;
    wire c175;
    assign in175_1 = {pp10[94]};
    assign in175_2 = {pp11[93]};
    Full_Adder FA_175(s175, c175, in175_1, in175_2, pp9[95]);
    wire[0:0] s176, in176_1, in176_2;
    wire c176;
    assign in176_1 = {pp13[91]};
    assign in176_2 = {pp14[90]};
    Full_Adder FA_176(s176, c176, in176_1, in176_2, pp12[92]);
    wire[0:0] s177, in177_1, in177_2;
    wire c177;
    assign in177_1 = {pp16[88]};
    assign in177_2 = {pp17[87]};
    Full_Adder FA_177(s177, c177, in177_1, in177_2, pp15[89]);
    wire[0:0] s178, in178_1, in178_2;
    wire c178;
    assign in178_1 = {pp19[85]};
    assign in178_2 = {pp20[84]};
    Full_Adder FA_178(s178, c178, in178_1, in178_2, pp18[86]);
    wire[0:0] s179, in179_1, in179_2;
    wire c179;
    assign in179_1 = {pp22[82]};
    assign in179_2 = {pp23[81]};
    Full_Adder FA_179(s179, c179, in179_1, in179_2, pp21[83]);
    wire[0:0] s180, in180_1, in180_2;
    wire c180;
    assign in180_1 = {pp25[79]};
    assign in180_2 = {pp26[78]};
    Full_Adder FA_180(s180, c180, in180_1, in180_2, pp24[80]);
    wire[0:0] s181, in181_1, in181_2;
    wire c181;
    assign in181_1 = {pp28[76]};
    assign in181_2 = {pp29[75]};
    Full_Adder FA_181(s181, c181, in181_1, in181_2, pp27[77]);
    wire[0:0] s182, in182_1, in182_2;
    wire c182;
    assign in182_1 = {pp31[73]};
    assign in182_2 = {pp32[72]};
    Full_Adder FA_182(s182, c182, in182_1, in182_2, pp30[74]);
    wire[0:0] s183, in183_1, in183_2;
    wire c183;
    assign in183_1 = {pp34[70]};
    assign in183_2 = {pp35[69]};
    Full_Adder FA_183(s183, c183, in183_1, in183_2, pp33[71]);
    wire[0:0] s184, in184_1, in184_2;
    wire c184;
    assign in184_1 = {pp37[67]};
    assign in184_2 = {pp38[66]};
    Full_Adder FA_184(s184, c184, in184_1, in184_2, pp36[68]);
    wire[0:0] s185, in185_1, in185_2;
    wire c185;
    assign in185_1 = {pp40[64]};
    assign in185_2 = {pp41[63]};
    Full_Adder FA_185(s185, c185, in185_1, in185_2, pp39[65]);
    wire[0:0] s186, in186_1, in186_2;
    wire c186;
    assign in186_1 = {pp43[61]};
    assign in186_2 = {pp44[60]};
    Full_Adder FA_186(s186, c186, in186_1, in186_2, pp42[62]);
    wire[0:0] s187, in187_1, in187_2;
    wire c187;
    assign in187_1 = {pp46[58]};
    assign in187_2 = {pp47[57]};
    Full_Adder FA_187(s187, c187, in187_1, in187_2, pp45[59]);
    wire[0:0] s188, in188_1, in188_2;
    wire c188;
    assign in188_1 = {pp49[55]};
    assign in188_2 = {pp50[54]};
    Full_Adder FA_188(s188, c188, in188_1, in188_2, pp48[56]);
    wire[0:0] s189, in189_1, in189_2;
    wire c189;
    assign in189_1 = {pp52[52]};
    assign in189_2 = {pp53[51]};
    Full_Adder FA_189(s189, c189, in189_1, in189_2, pp51[53]);
    wire[0:0] s190, in190_1, in190_2;
    wire c190;
    assign in190_1 = {pp54[50]};
    assign in190_2 = {pp55[49]};
    Half_Adder HA_190(s190, c190, in190_1, in190_2);
    wire[0:0] s191, in191_1, in191_2;
    wire c191;
    assign in191_1 = {pp1[104]};
    assign in191_2 = {pp2[103]};
    Full_Adder FA_191(s191, c191, in191_1, in191_2, pp0[105]);
    wire[0:0] s192, in192_1, in192_2;
    wire c192;
    assign in192_1 = {pp4[101]};
    assign in192_2 = {pp5[100]};
    Full_Adder FA_192(s192, c192, in192_1, in192_2, pp3[102]);
    wire[0:0] s193, in193_1, in193_2;
    wire c193;
    assign in193_1 = {pp7[98]};
    assign in193_2 = {pp8[97]};
    Full_Adder FA_193(s193, c193, in193_1, in193_2, pp6[99]);
    wire[0:0] s194, in194_1, in194_2;
    wire c194;
    assign in194_1 = {pp10[95]};
    assign in194_2 = {pp11[94]};
    Full_Adder FA_194(s194, c194, in194_1, in194_2, pp9[96]);
    wire[0:0] s195, in195_1, in195_2;
    wire c195;
    assign in195_1 = {pp13[92]};
    assign in195_2 = {pp14[91]};
    Full_Adder FA_195(s195, c195, in195_1, in195_2, pp12[93]);
    wire[0:0] s196, in196_1, in196_2;
    wire c196;
    assign in196_1 = {pp16[89]};
    assign in196_2 = {pp17[88]};
    Full_Adder FA_196(s196, c196, in196_1, in196_2, pp15[90]);
    wire[0:0] s197, in197_1, in197_2;
    wire c197;
    assign in197_1 = {pp19[86]};
    assign in197_2 = {pp20[85]};
    Full_Adder FA_197(s197, c197, in197_1, in197_2, pp18[87]);
    wire[0:0] s198, in198_1, in198_2;
    wire c198;
    assign in198_1 = {pp22[83]};
    assign in198_2 = {pp23[82]};
    Full_Adder FA_198(s198, c198, in198_1, in198_2, pp21[84]);
    wire[0:0] s199, in199_1, in199_2;
    wire c199;
    assign in199_1 = {pp25[80]};
    assign in199_2 = {pp26[79]};
    Full_Adder FA_199(s199, c199, in199_1, in199_2, pp24[81]);
    wire[0:0] s200, in200_1, in200_2;
    wire c200;
    assign in200_1 = {pp28[77]};
    assign in200_2 = {pp29[76]};
    Full_Adder FA_200(s200, c200, in200_1, in200_2, pp27[78]);
    wire[0:0] s201, in201_1, in201_2;
    wire c201;
    assign in201_1 = {pp31[74]};
    assign in201_2 = {pp32[73]};
    Full_Adder FA_201(s201, c201, in201_1, in201_2, pp30[75]);
    wire[0:0] s202, in202_1, in202_2;
    wire c202;
    assign in202_1 = {pp34[71]};
    assign in202_2 = {pp35[70]};
    Full_Adder FA_202(s202, c202, in202_1, in202_2, pp33[72]);
    wire[0:0] s203, in203_1, in203_2;
    wire c203;
    assign in203_1 = {pp37[68]};
    assign in203_2 = {pp38[67]};
    Full_Adder FA_203(s203, c203, in203_1, in203_2, pp36[69]);
    wire[0:0] s204, in204_1, in204_2;
    wire c204;
    assign in204_1 = {pp40[65]};
    assign in204_2 = {pp41[64]};
    Full_Adder FA_204(s204, c204, in204_1, in204_2, pp39[66]);
    wire[0:0] s205, in205_1, in205_2;
    wire c205;
    assign in205_1 = {pp43[62]};
    assign in205_2 = {pp44[61]};
    Full_Adder FA_205(s205, c205, in205_1, in205_2, pp42[63]);
    wire[0:0] s206, in206_1, in206_2;
    wire c206;
    assign in206_1 = {pp46[59]};
    assign in206_2 = {pp47[58]};
    Full_Adder FA_206(s206, c206, in206_1, in206_2, pp45[60]);
    wire[0:0] s207, in207_1, in207_2;
    wire c207;
    assign in207_1 = {pp49[56]};
    assign in207_2 = {pp50[55]};
    Full_Adder FA_207(s207, c207, in207_1, in207_2, pp48[57]);
    wire[0:0] s208, in208_1, in208_2;
    wire c208;
    assign in208_1 = {pp52[53]};
    assign in208_2 = {pp53[52]};
    Full_Adder FA_208(s208, c208, in208_1, in208_2, pp51[54]);
    wire[0:0] s209, in209_1, in209_2;
    wire c209;
    assign in209_1 = {pp55[50]};
    assign in209_2 = {pp56[49]};
    Full_Adder FA_209(s209, c209, in209_1, in209_2, pp54[51]);
    wire[0:0] s210, in210_1, in210_2;
    wire c210;
    assign in210_1 = {pp57[48]};
    assign in210_2 = {pp58[47]};
    Half_Adder HA_210(s210, c210, in210_1, in210_2);
    wire[0:0] s211, in211_1, in211_2;
    wire c211;
    assign in211_1 = {pp1[105]};
    assign in211_2 = {pp2[104]};
    Full_Adder FA_211(s211, c211, in211_1, in211_2, pp0[106]);
    wire[0:0] s212, in212_1, in212_2;
    wire c212;
    assign in212_1 = {pp4[102]};
    assign in212_2 = {pp5[101]};
    Full_Adder FA_212(s212, c212, in212_1, in212_2, pp3[103]);
    wire[0:0] s213, in213_1, in213_2;
    wire c213;
    assign in213_1 = {pp7[99]};
    assign in213_2 = {pp8[98]};
    Full_Adder FA_213(s213, c213, in213_1, in213_2, pp6[100]);
    wire[0:0] s214, in214_1, in214_2;
    wire c214;
    assign in214_1 = {pp10[96]};
    assign in214_2 = {pp11[95]};
    Full_Adder FA_214(s214, c214, in214_1, in214_2, pp9[97]);
    wire[0:0] s215, in215_1, in215_2;
    wire c215;
    assign in215_1 = {pp13[93]};
    assign in215_2 = {pp14[92]};
    Full_Adder FA_215(s215, c215, in215_1, in215_2, pp12[94]);
    wire[0:0] s216, in216_1, in216_2;
    wire c216;
    assign in216_1 = {pp16[90]};
    assign in216_2 = {pp17[89]};
    Full_Adder FA_216(s216, c216, in216_1, in216_2, pp15[91]);
    wire[0:0] s217, in217_1, in217_2;
    wire c217;
    assign in217_1 = {pp19[87]};
    assign in217_2 = {pp20[86]};
    Full_Adder FA_217(s217, c217, in217_1, in217_2, pp18[88]);
    wire[0:0] s218, in218_1, in218_2;
    wire c218;
    assign in218_1 = {pp22[84]};
    assign in218_2 = {pp23[83]};
    Full_Adder FA_218(s218, c218, in218_1, in218_2, pp21[85]);
    wire[0:0] s219, in219_1, in219_2;
    wire c219;
    assign in219_1 = {pp25[81]};
    assign in219_2 = {pp26[80]};
    Full_Adder FA_219(s219, c219, in219_1, in219_2, pp24[82]);
    wire[0:0] s220, in220_1, in220_2;
    wire c220;
    assign in220_1 = {pp28[78]};
    assign in220_2 = {pp29[77]};
    Full_Adder FA_220(s220, c220, in220_1, in220_2, pp27[79]);
    wire[0:0] s221, in221_1, in221_2;
    wire c221;
    assign in221_1 = {pp31[75]};
    assign in221_2 = {pp32[74]};
    Full_Adder FA_221(s221, c221, in221_1, in221_2, pp30[76]);
    wire[0:0] s222, in222_1, in222_2;
    wire c222;
    assign in222_1 = {pp34[72]};
    assign in222_2 = {pp35[71]};
    Full_Adder FA_222(s222, c222, in222_1, in222_2, pp33[73]);
    wire[0:0] s223, in223_1, in223_2;
    wire c223;
    assign in223_1 = {pp37[69]};
    assign in223_2 = {pp38[68]};
    Full_Adder FA_223(s223, c223, in223_1, in223_2, pp36[70]);
    wire[0:0] s224, in224_1, in224_2;
    wire c224;
    assign in224_1 = {pp40[66]};
    assign in224_2 = {pp41[65]};
    Full_Adder FA_224(s224, c224, in224_1, in224_2, pp39[67]);
    wire[0:0] s225, in225_1, in225_2;
    wire c225;
    assign in225_1 = {pp43[63]};
    assign in225_2 = {pp44[62]};
    Full_Adder FA_225(s225, c225, in225_1, in225_2, pp42[64]);
    wire[0:0] s226, in226_1, in226_2;
    wire c226;
    assign in226_1 = {pp46[60]};
    assign in226_2 = {pp47[59]};
    Full_Adder FA_226(s226, c226, in226_1, in226_2, pp45[61]);
    wire[0:0] s227, in227_1, in227_2;
    wire c227;
    assign in227_1 = {pp49[57]};
    assign in227_2 = {pp50[56]};
    Full_Adder FA_227(s227, c227, in227_1, in227_2, pp48[58]);
    wire[0:0] s228, in228_1, in228_2;
    wire c228;
    assign in228_1 = {pp52[54]};
    assign in228_2 = {pp53[53]};
    Full_Adder FA_228(s228, c228, in228_1, in228_2, pp51[55]);
    wire[0:0] s229, in229_1, in229_2;
    wire c229;
    assign in229_1 = {pp55[51]};
    assign in229_2 = {pp56[50]};
    Full_Adder FA_229(s229, c229, in229_1, in229_2, pp54[52]);
    wire[0:0] s230, in230_1, in230_2;
    wire c230;
    assign in230_1 = {pp58[48]};
    assign in230_2 = {pp59[47]};
    Full_Adder FA_230(s230, c230, in230_1, in230_2, pp57[49]);
    wire[0:0] s231, in231_1, in231_2;
    wire c231;
    assign in231_1 = {pp60[46]};
    assign in231_2 = {pp61[45]};
    Half_Adder HA_231(s231, c231, in231_1, in231_2);
    wire[0:0] s232, in232_1, in232_2;
    wire c232;
    assign in232_1 = {pp1[106]};
    assign in232_2 = {pp2[105]};
    Full_Adder FA_232(s232, c232, in232_1, in232_2, pp0[107]);
    wire[0:0] s233, in233_1, in233_2;
    wire c233;
    assign in233_1 = {pp4[103]};
    assign in233_2 = {pp5[102]};
    Full_Adder FA_233(s233, c233, in233_1, in233_2, pp3[104]);
    wire[0:0] s234, in234_1, in234_2;
    wire c234;
    assign in234_1 = {pp7[100]};
    assign in234_2 = {pp8[99]};
    Full_Adder FA_234(s234, c234, in234_1, in234_2, pp6[101]);
    wire[0:0] s235, in235_1, in235_2;
    wire c235;
    assign in235_1 = {pp10[97]};
    assign in235_2 = {pp11[96]};
    Full_Adder FA_235(s235, c235, in235_1, in235_2, pp9[98]);
    wire[0:0] s236, in236_1, in236_2;
    wire c236;
    assign in236_1 = {pp13[94]};
    assign in236_2 = {pp14[93]};
    Full_Adder FA_236(s236, c236, in236_1, in236_2, pp12[95]);
    wire[0:0] s237, in237_1, in237_2;
    wire c237;
    assign in237_1 = {pp16[91]};
    assign in237_2 = {pp17[90]};
    Full_Adder FA_237(s237, c237, in237_1, in237_2, pp15[92]);
    wire[0:0] s238, in238_1, in238_2;
    wire c238;
    assign in238_1 = {pp19[88]};
    assign in238_2 = {pp20[87]};
    Full_Adder FA_238(s238, c238, in238_1, in238_2, pp18[89]);
    wire[0:0] s239, in239_1, in239_2;
    wire c239;
    assign in239_1 = {pp22[85]};
    assign in239_2 = {pp23[84]};
    Full_Adder FA_239(s239, c239, in239_1, in239_2, pp21[86]);
    wire[0:0] s240, in240_1, in240_2;
    wire c240;
    assign in240_1 = {pp25[82]};
    assign in240_2 = {pp26[81]};
    Full_Adder FA_240(s240, c240, in240_1, in240_2, pp24[83]);
    wire[0:0] s241, in241_1, in241_2;
    wire c241;
    assign in241_1 = {pp28[79]};
    assign in241_2 = {pp29[78]};
    Full_Adder FA_241(s241, c241, in241_1, in241_2, pp27[80]);
    wire[0:0] s242, in242_1, in242_2;
    wire c242;
    assign in242_1 = {pp31[76]};
    assign in242_2 = {pp32[75]};
    Full_Adder FA_242(s242, c242, in242_1, in242_2, pp30[77]);
    wire[0:0] s243, in243_1, in243_2;
    wire c243;
    assign in243_1 = {pp34[73]};
    assign in243_2 = {pp35[72]};
    Full_Adder FA_243(s243, c243, in243_1, in243_2, pp33[74]);
    wire[0:0] s244, in244_1, in244_2;
    wire c244;
    assign in244_1 = {pp37[70]};
    assign in244_2 = {pp38[69]};
    Full_Adder FA_244(s244, c244, in244_1, in244_2, pp36[71]);
    wire[0:0] s245, in245_1, in245_2;
    wire c245;
    assign in245_1 = {pp40[67]};
    assign in245_2 = {pp41[66]};
    Full_Adder FA_245(s245, c245, in245_1, in245_2, pp39[68]);
    wire[0:0] s246, in246_1, in246_2;
    wire c246;
    assign in246_1 = {pp43[64]};
    assign in246_2 = {pp44[63]};
    Full_Adder FA_246(s246, c246, in246_1, in246_2, pp42[65]);
    wire[0:0] s247, in247_1, in247_2;
    wire c247;
    assign in247_1 = {pp46[61]};
    assign in247_2 = {pp47[60]};
    Full_Adder FA_247(s247, c247, in247_1, in247_2, pp45[62]);
    wire[0:0] s248, in248_1, in248_2;
    wire c248;
    assign in248_1 = {pp49[58]};
    assign in248_2 = {pp50[57]};
    Full_Adder FA_248(s248, c248, in248_1, in248_2, pp48[59]);
    wire[0:0] s249, in249_1, in249_2;
    wire c249;
    assign in249_1 = {pp52[55]};
    assign in249_2 = {pp53[54]};
    Full_Adder FA_249(s249, c249, in249_1, in249_2, pp51[56]);
    wire[0:0] s250, in250_1, in250_2;
    wire c250;
    assign in250_1 = {pp55[52]};
    assign in250_2 = {pp56[51]};
    Full_Adder FA_250(s250, c250, in250_1, in250_2, pp54[53]);
    wire[0:0] s251, in251_1, in251_2;
    wire c251;
    assign in251_1 = {pp58[49]};
    assign in251_2 = {pp59[48]};
    Full_Adder FA_251(s251, c251, in251_1, in251_2, pp57[50]);
    wire[0:0] s252, in252_1, in252_2;
    wire c252;
    assign in252_1 = {pp61[46]};
    assign in252_2 = {pp62[45]};
    Full_Adder FA_252(s252, c252, in252_1, in252_2, pp60[47]);
    wire[0:0] s253, in253_1, in253_2;
    wire c253;
    assign in253_1 = {pp63[44]};
    assign in253_2 = {pp64[43]};
    Half_Adder HA_253(s253, c253, in253_1, in253_2);
    wire[0:0] s254, in254_1, in254_2;
    wire c254;
    assign in254_1 = {pp1[107]};
    assign in254_2 = {pp2[106]};
    Full_Adder FA_254(s254, c254, in254_1, in254_2, pp0[108]);
    wire[0:0] s255, in255_1, in255_2;
    wire c255;
    assign in255_1 = {pp4[104]};
    assign in255_2 = {pp5[103]};
    Full_Adder FA_255(s255, c255, in255_1, in255_2, pp3[105]);
    wire[0:0] s256, in256_1, in256_2;
    wire c256;
    assign in256_1 = {pp7[101]};
    assign in256_2 = {pp8[100]};
    Full_Adder FA_256(s256, c256, in256_1, in256_2, pp6[102]);
    wire[0:0] s257, in257_1, in257_2;
    wire c257;
    assign in257_1 = {pp10[98]};
    assign in257_2 = {pp11[97]};
    Full_Adder FA_257(s257, c257, in257_1, in257_2, pp9[99]);
    wire[0:0] s258, in258_1, in258_2;
    wire c258;
    assign in258_1 = {pp13[95]};
    assign in258_2 = {pp14[94]};
    Full_Adder FA_258(s258, c258, in258_1, in258_2, pp12[96]);
    wire[0:0] s259, in259_1, in259_2;
    wire c259;
    assign in259_1 = {pp16[92]};
    assign in259_2 = {pp17[91]};
    Full_Adder FA_259(s259, c259, in259_1, in259_2, pp15[93]);
    wire[0:0] s260, in260_1, in260_2;
    wire c260;
    assign in260_1 = {pp19[89]};
    assign in260_2 = {pp20[88]};
    Full_Adder FA_260(s260, c260, in260_1, in260_2, pp18[90]);
    wire[0:0] s261, in261_1, in261_2;
    wire c261;
    assign in261_1 = {pp22[86]};
    assign in261_2 = {pp23[85]};
    Full_Adder FA_261(s261, c261, in261_1, in261_2, pp21[87]);
    wire[0:0] s262, in262_1, in262_2;
    wire c262;
    assign in262_1 = {pp25[83]};
    assign in262_2 = {pp26[82]};
    Full_Adder FA_262(s262, c262, in262_1, in262_2, pp24[84]);
    wire[0:0] s263, in263_1, in263_2;
    wire c263;
    assign in263_1 = {pp28[80]};
    assign in263_2 = {pp29[79]};
    Full_Adder FA_263(s263, c263, in263_1, in263_2, pp27[81]);
    wire[0:0] s264, in264_1, in264_2;
    wire c264;
    assign in264_1 = {pp31[77]};
    assign in264_2 = {pp32[76]};
    Full_Adder FA_264(s264, c264, in264_1, in264_2, pp30[78]);
    wire[0:0] s265, in265_1, in265_2;
    wire c265;
    assign in265_1 = {pp34[74]};
    assign in265_2 = {pp35[73]};
    Full_Adder FA_265(s265, c265, in265_1, in265_2, pp33[75]);
    wire[0:0] s266, in266_1, in266_2;
    wire c266;
    assign in266_1 = {pp37[71]};
    assign in266_2 = {pp38[70]};
    Full_Adder FA_266(s266, c266, in266_1, in266_2, pp36[72]);
    wire[0:0] s267, in267_1, in267_2;
    wire c267;
    assign in267_1 = {pp40[68]};
    assign in267_2 = {pp41[67]};
    Full_Adder FA_267(s267, c267, in267_1, in267_2, pp39[69]);
    wire[0:0] s268, in268_1, in268_2;
    wire c268;
    assign in268_1 = {pp43[65]};
    assign in268_2 = {pp44[64]};
    Full_Adder FA_268(s268, c268, in268_1, in268_2, pp42[66]);
    wire[0:0] s269, in269_1, in269_2;
    wire c269;
    assign in269_1 = {pp46[62]};
    assign in269_2 = {pp47[61]};
    Full_Adder FA_269(s269, c269, in269_1, in269_2, pp45[63]);
    wire[0:0] s270, in270_1, in270_2;
    wire c270;
    assign in270_1 = {pp49[59]};
    assign in270_2 = {pp50[58]};
    Full_Adder FA_270(s270, c270, in270_1, in270_2, pp48[60]);
    wire[0:0] s271, in271_1, in271_2;
    wire c271;
    assign in271_1 = {pp52[56]};
    assign in271_2 = {pp53[55]};
    Full_Adder FA_271(s271, c271, in271_1, in271_2, pp51[57]);
    wire[0:0] s272, in272_1, in272_2;
    wire c272;
    assign in272_1 = {pp55[53]};
    assign in272_2 = {pp56[52]};
    Full_Adder FA_272(s272, c272, in272_1, in272_2, pp54[54]);
    wire[0:0] s273, in273_1, in273_2;
    wire c273;
    assign in273_1 = {pp58[50]};
    assign in273_2 = {pp59[49]};
    Full_Adder FA_273(s273, c273, in273_1, in273_2, pp57[51]);
    wire[0:0] s274, in274_1, in274_2;
    wire c274;
    assign in274_1 = {pp61[47]};
    assign in274_2 = {pp62[46]};
    Full_Adder FA_274(s274, c274, in274_1, in274_2, pp60[48]);
    wire[0:0] s275, in275_1, in275_2;
    wire c275;
    assign in275_1 = {pp64[44]};
    assign in275_2 = {pp65[43]};
    Full_Adder FA_275(s275, c275, in275_1, in275_2, pp63[45]);
    wire[0:0] s276, in276_1, in276_2;
    wire c276;
    assign in276_1 = {pp66[42]};
    assign in276_2 = {pp67[41]};
    Half_Adder HA_276(s276, c276, in276_1, in276_2);
    wire[0:0] s277, in277_1, in277_2;
    wire c277;
    assign in277_1 = {pp1[108]};
    assign in277_2 = {pp2[107]};
    Full_Adder FA_277(s277, c277, in277_1, in277_2, pp0[109]);
    wire[0:0] s278, in278_1, in278_2;
    wire c278;
    assign in278_1 = {pp4[105]};
    assign in278_2 = {pp5[104]};
    Full_Adder FA_278(s278, c278, in278_1, in278_2, pp3[106]);
    wire[0:0] s279, in279_1, in279_2;
    wire c279;
    assign in279_1 = {pp7[102]};
    assign in279_2 = {pp8[101]};
    Full_Adder FA_279(s279, c279, in279_1, in279_2, pp6[103]);
    wire[0:0] s280, in280_1, in280_2;
    wire c280;
    assign in280_1 = {pp10[99]};
    assign in280_2 = {pp11[98]};
    Full_Adder FA_280(s280, c280, in280_1, in280_2, pp9[100]);
    wire[0:0] s281, in281_1, in281_2;
    wire c281;
    assign in281_1 = {pp13[96]};
    assign in281_2 = {pp14[95]};
    Full_Adder FA_281(s281, c281, in281_1, in281_2, pp12[97]);
    wire[0:0] s282, in282_1, in282_2;
    wire c282;
    assign in282_1 = {pp16[93]};
    assign in282_2 = {pp17[92]};
    Full_Adder FA_282(s282, c282, in282_1, in282_2, pp15[94]);
    wire[0:0] s283, in283_1, in283_2;
    wire c283;
    assign in283_1 = {pp19[90]};
    assign in283_2 = {pp20[89]};
    Full_Adder FA_283(s283, c283, in283_1, in283_2, pp18[91]);
    wire[0:0] s284, in284_1, in284_2;
    wire c284;
    assign in284_1 = {pp22[87]};
    assign in284_2 = {pp23[86]};
    Full_Adder FA_284(s284, c284, in284_1, in284_2, pp21[88]);
    wire[0:0] s285, in285_1, in285_2;
    wire c285;
    assign in285_1 = {pp25[84]};
    assign in285_2 = {pp26[83]};
    Full_Adder FA_285(s285, c285, in285_1, in285_2, pp24[85]);
    wire[0:0] s286, in286_1, in286_2;
    wire c286;
    assign in286_1 = {pp28[81]};
    assign in286_2 = {pp29[80]};
    Full_Adder FA_286(s286, c286, in286_1, in286_2, pp27[82]);
    wire[0:0] s287, in287_1, in287_2;
    wire c287;
    assign in287_1 = {pp31[78]};
    assign in287_2 = {pp32[77]};
    Full_Adder FA_287(s287, c287, in287_1, in287_2, pp30[79]);
    wire[0:0] s288, in288_1, in288_2;
    wire c288;
    assign in288_1 = {pp34[75]};
    assign in288_2 = {pp35[74]};
    Full_Adder FA_288(s288, c288, in288_1, in288_2, pp33[76]);
    wire[0:0] s289, in289_1, in289_2;
    wire c289;
    assign in289_1 = {pp37[72]};
    assign in289_2 = {pp38[71]};
    Full_Adder FA_289(s289, c289, in289_1, in289_2, pp36[73]);
    wire[0:0] s290, in290_1, in290_2;
    wire c290;
    assign in290_1 = {pp40[69]};
    assign in290_2 = {pp41[68]};
    Full_Adder FA_290(s290, c290, in290_1, in290_2, pp39[70]);
    wire[0:0] s291, in291_1, in291_2;
    wire c291;
    assign in291_1 = {pp43[66]};
    assign in291_2 = {pp44[65]};
    Full_Adder FA_291(s291, c291, in291_1, in291_2, pp42[67]);
    wire[0:0] s292, in292_1, in292_2;
    wire c292;
    assign in292_1 = {pp46[63]};
    assign in292_2 = {pp47[62]};
    Full_Adder FA_292(s292, c292, in292_1, in292_2, pp45[64]);
    wire[0:0] s293, in293_1, in293_2;
    wire c293;
    assign in293_1 = {pp49[60]};
    assign in293_2 = {pp50[59]};
    Full_Adder FA_293(s293, c293, in293_1, in293_2, pp48[61]);
    wire[0:0] s294, in294_1, in294_2;
    wire c294;
    assign in294_1 = {pp52[57]};
    assign in294_2 = {pp53[56]};
    Full_Adder FA_294(s294, c294, in294_1, in294_2, pp51[58]);
    wire[0:0] s295, in295_1, in295_2;
    wire c295;
    assign in295_1 = {pp55[54]};
    assign in295_2 = {pp56[53]};
    Full_Adder FA_295(s295, c295, in295_1, in295_2, pp54[55]);
    wire[0:0] s296, in296_1, in296_2;
    wire c296;
    assign in296_1 = {pp58[51]};
    assign in296_2 = {pp59[50]};
    Full_Adder FA_296(s296, c296, in296_1, in296_2, pp57[52]);
    wire[0:0] s297, in297_1, in297_2;
    wire c297;
    assign in297_1 = {pp61[48]};
    assign in297_2 = {pp62[47]};
    Full_Adder FA_297(s297, c297, in297_1, in297_2, pp60[49]);
    wire[0:0] s298, in298_1, in298_2;
    wire c298;
    assign in298_1 = {pp64[45]};
    assign in298_2 = {pp65[44]};
    Full_Adder FA_298(s298, c298, in298_1, in298_2, pp63[46]);
    wire[0:0] s299, in299_1, in299_2;
    wire c299;
    assign in299_1 = {pp67[42]};
    assign in299_2 = {pp68[41]};
    Full_Adder FA_299(s299, c299, in299_1, in299_2, pp66[43]);
    wire[0:0] s300, in300_1, in300_2;
    wire c300;
    assign in300_1 = {pp69[40]};
    assign in300_2 = {pp70[39]};
    Half_Adder HA_300(s300, c300, in300_1, in300_2);
    wire[0:0] s301, in301_1, in301_2;
    wire c301;
    assign in301_1 = {pp1[109]};
    assign in301_2 = {pp2[108]};
    Full_Adder FA_301(s301, c301, in301_1, in301_2, pp0[110]);
    wire[0:0] s302, in302_1, in302_2;
    wire c302;
    assign in302_1 = {pp4[106]};
    assign in302_2 = {pp5[105]};
    Full_Adder FA_302(s302, c302, in302_1, in302_2, pp3[107]);
    wire[0:0] s303, in303_1, in303_2;
    wire c303;
    assign in303_1 = {pp7[103]};
    assign in303_2 = {pp8[102]};
    Full_Adder FA_303(s303, c303, in303_1, in303_2, pp6[104]);
    wire[0:0] s304, in304_1, in304_2;
    wire c304;
    assign in304_1 = {pp10[100]};
    assign in304_2 = {pp11[99]};
    Full_Adder FA_304(s304, c304, in304_1, in304_2, pp9[101]);
    wire[0:0] s305, in305_1, in305_2;
    wire c305;
    assign in305_1 = {pp13[97]};
    assign in305_2 = {pp14[96]};
    Full_Adder FA_305(s305, c305, in305_1, in305_2, pp12[98]);
    wire[0:0] s306, in306_1, in306_2;
    wire c306;
    assign in306_1 = {pp16[94]};
    assign in306_2 = {pp17[93]};
    Full_Adder FA_306(s306, c306, in306_1, in306_2, pp15[95]);
    wire[0:0] s307, in307_1, in307_2;
    wire c307;
    assign in307_1 = {pp19[91]};
    assign in307_2 = {pp20[90]};
    Full_Adder FA_307(s307, c307, in307_1, in307_2, pp18[92]);
    wire[0:0] s308, in308_1, in308_2;
    wire c308;
    assign in308_1 = {pp22[88]};
    assign in308_2 = {pp23[87]};
    Full_Adder FA_308(s308, c308, in308_1, in308_2, pp21[89]);
    wire[0:0] s309, in309_1, in309_2;
    wire c309;
    assign in309_1 = {pp25[85]};
    assign in309_2 = {pp26[84]};
    Full_Adder FA_309(s309, c309, in309_1, in309_2, pp24[86]);
    wire[0:0] s310, in310_1, in310_2;
    wire c310;
    assign in310_1 = {pp28[82]};
    assign in310_2 = {pp29[81]};
    Full_Adder FA_310(s310, c310, in310_1, in310_2, pp27[83]);
    wire[0:0] s311, in311_1, in311_2;
    wire c311;
    assign in311_1 = {pp31[79]};
    assign in311_2 = {pp32[78]};
    Full_Adder FA_311(s311, c311, in311_1, in311_2, pp30[80]);
    wire[0:0] s312, in312_1, in312_2;
    wire c312;
    assign in312_1 = {pp34[76]};
    assign in312_2 = {pp35[75]};
    Full_Adder FA_312(s312, c312, in312_1, in312_2, pp33[77]);
    wire[0:0] s313, in313_1, in313_2;
    wire c313;
    assign in313_1 = {pp37[73]};
    assign in313_2 = {pp38[72]};
    Full_Adder FA_313(s313, c313, in313_1, in313_2, pp36[74]);
    wire[0:0] s314, in314_1, in314_2;
    wire c314;
    assign in314_1 = {pp40[70]};
    assign in314_2 = {pp41[69]};
    Full_Adder FA_314(s314, c314, in314_1, in314_2, pp39[71]);
    wire[0:0] s315, in315_1, in315_2;
    wire c315;
    assign in315_1 = {pp43[67]};
    assign in315_2 = {pp44[66]};
    Full_Adder FA_315(s315, c315, in315_1, in315_2, pp42[68]);
    wire[0:0] s316, in316_1, in316_2;
    wire c316;
    assign in316_1 = {pp46[64]};
    assign in316_2 = {pp47[63]};
    Full_Adder FA_316(s316, c316, in316_1, in316_2, pp45[65]);
    wire[0:0] s317, in317_1, in317_2;
    wire c317;
    assign in317_1 = {pp49[61]};
    assign in317_2 = {pp50[60]};
    Full_Adder FA_317(s317, c317, in317_1, in317_2, pp48[62]);
    wire[0:0] s318, in318_1, in318_2;
    wire c318;
    assign in318_1 = {pp52[58]};
    assign in318_2 = {pp53[57]};
    Full_Adder FA_318(s318, c318, in318_1, in318_2, pp51[59]);
    wire[0:0] s319, in319_1, in319_2;
    wire c319;
    assign in319_1 = {pp55[55]};
    assign in319_2 = {pp56[54]};
    Full_Adder FA_319(s319, c319, in319_1, in319_2, pp54[56]);
    wire[0:0] s320, in320_1, in320_2;
    wire c320;
    assign in320_1 = {pp58[52]};
    assign in320_2 = {pp59[51]};
    Full_Adder FA_320(s320, c320, in320_1, in320_2, pp57[53]);
    wire[0:0] s321, in321_1, in321_2;
    wire c321;
    assign in321_1 = {pp61[49]};
    assign in321_2 = {pp62[48]};
    Full_Adder FA_321(s321, c321, in321_1, in321_2, pp60[50]);
    wire[0:0] s322, in322_1, in322_2;
    wire c322;
    assign in322_1 = {pp64[46]};
    assign in322_2 = {pp65[45]};
    Full_Adder FA_322(s322, c322, in322_1, in322_2, pp63[47]);
    wire[0:0] s323, in323_1, in323_2;
    wire c323;
    assign in323_1 = {pp67[43]};
    assign in323_2 = {pp68[42]};
    Full_Adder FA_323(s323, c323, in323_1, in323_2, pp66[44]);
    wire[0:0] s324, in324_1, in324_2;
    wire c324;
    assign in324_1 = {pp70[40]};
    assign in324_2 = {pp71[39]};
    Full_Adder FA_324(s324, c324, in324_1, in324_2, pp69[41]);
    wire[0:0] s325, in325_1, in325_2;
    wire c325;
    assign in325_1 = {pp72[38]};
    assign in325_2 = {pp73[37]};
    Half_Adder HA_325(s325, c325, in325_1, in325_2);
    wire[0:0] s326, in326_1, in326_2;
    wire c326;
    assign in326_1 = {pp1[110]};
    assign in326_2 = {pp2[109]};
    Full_Adder FA_326(s326, c326, in326_1, in326_2, pp0[111]);
    wire[0:0] s327, in327_1, in327_2;
    wire c327;
    assign in327_1 = {pp4[107]};
    assign in327_2 = {pp5[106]};
    Full_Adder FA_327(s327, c327, in327_1, in327_2, pp3[108]);
    wire[0:0] s328, in328_1, in328_2;
    wire c328;
    assign in328_1 = {pp7[104]};
    assign in328_2 = {pp8[103]};
    Full_Adder FA_328(s328, c328, in328_1, in328_2, pp6[105]);
    wire[0:0] s329, in329_1, in329_2;
    wire c329;
    assign in329_1 = {pp10[101]};
    assign in329_2 = {pp11[100]};
    Full_Adder FA_329(s329, c329, in329_1, in329_2, pp9[102]);
    wire[0:0] s330, in330_1, in330_2;
    wire c330;
    assign in330_1 = {pp13[98]};
    assign in330_2 = {pp14[97]};
    Full_Adder FA_330(s330, c330, in330_1, in330_2, pp12[99]);
    wire[0:0] s331, in331_1, in331_2;
    wire c331;
    assign in331_1 = {pp16[95]};
    assign in331_2 = {pp17[94]};
    Full_Adder FA_331(s331, c331, in331_1, in331_2, pp15[96]);
    wire[0:0] s332, in332_1, in332_2;
    wire c332;
    assign in332_1 = {pp19[92]};
    assign in332_2 = {pp20[91]};
    Full_Adder FA_332(s332, c332, in332_1, in332_2, pp18[93]);
    wire[0:0] s333, in333_1, in333_2;
    wire c333;
    assign in333_1 = {pp22[89]};
    assign in333_2 = {pp23[88]};
    Full_Adder FA_333(s333, c333, in333_1, in333_2, pp21[90]);
    wire[0:0] s334, in334_1, in334_2;
    wire c334;
    assign in334_1 = {pp25[86]};
    assign in334_2 = {pp26[85]};
    Full_Adder FA_334(s334, c334, in334_1, in334_2, pp24[87]);
    wire[0:0] s335, in335_1, in335_2;
    wire c335;
    assign in335_1 = {pp28[83]};
    assign in335_2 = {pp29[82]};
    Full_Adder FA_335(s335, c335, in335_1, in335_2, pp27[84]);
    wire[0:0] s336, in336_1, in336_2;
    wire c336;
    assign in336_1 = {pp31[80]};
    assign in336_2 = {pp32[79]};
    Full_Adder FA_336(s336, c336, in336_1, in336_2, pp30[81]);
    wire[0:0] s337, in337_1, in337_2;
    wire c337;
    assign in337_1 = {pp34[77]};
    assign in337_2 = {pp35[76]};
    Full_Adder FA_337(s337, c337, in337_1, in337_2, pp33[78]);
    wire[0:0] s338, in338_1, in338_2;
    wire c338;
    assign in338_1 = {pp37[74]};
    assign in338_2 = {pp38[73]};
    Full_Adder FA_338(s338, c338, in338_1, in338_2, pp36[75]);
    wire[0:0] s339, in339_1, in339_2;
    wire c339;
    assign in339_1 = {pp40[71]};
    assign in339_2 = {pp41[70]};
    Full_Adder FA_339(s339, c339, in339_1, in339_2, pp39[72]);
    wire[0:0] s340, in340_1, in340_2;
    wire c340;
    assign in340_1 = {pp43[68]};
    assign in340_2 = {pp44[67]};
    Full_Adder FA_340(s340, c340, in340_1, in340_2, pp42[69]);
    wire[0:0] s341, in341_1, in341_2;
    wire c341;
    assign in341_1 = {pp46[65]};
    assign in341_2 = {pp47[64]};
    Full_Adder FA_341(s341, c341, in341_1, in341_2, pp45[66]);
    wire[0:0] s342, in342_1, in342_2;
    wire c342;
    assign in342_1 = {pp49[62]};
    assign in342_2 = {pp50[61]};
    Full_Adder FA_342(s342, c342, in342_1, in342_2, pp48[63]);
    wire[0:0] s343, in343_1, in343_2;
    wire c343;
    assign in343_1 = {pp52[59]};
    assign in343_2 = {pp53[58]};
    Full_Adder FA_343(s343, c343, in343_1, in343_2, pp51[60]);
    wire[0:0] s344, in344_1, in344_2;
    wire c344;
    assign in344_1 = {pp55[56]};
    assign in344_2 = {pp56[55]};
    Full_Adder FA_344(s344, c344, in344_1, in344_2, pp54[57]);
    wire[0:0] s345, in345_1, in345_2;
    wire c345;
    assign in345_1 = {pp58[53]};
    assign in345_2 = {pp59[52]};
    Full_Adder FA_345(s345, c345, in345_1, in345_2, pp57[54]);
    wire[0:0] s346, in346_1, in346_2;
    wire c346;
    assign in346_1 = {pp61[50]};
    assign in346_2 = {pp62[49]};
    Full_Adder FA_346(s346, c346, in346_1, in346_2, pp60[51]);
    wire[0:0] s347, in347_1, in347_2;
    wire c347;
    assign in347_1 = {pp64[47]};
    assign in347_2 = {pp65[46]};
    Full_Adder FA_347(s347, c347, in347_1, in347_2, pp63[48]);
    wire[0:0] s348, in348_1, in348_2;
    wire c348;
    assign in348_1 = {pp67[44]};
    assign in348_2 = {pp68[43]};
    Full_Adder FA_348(s348, c348, in348_1, in348_2, pp66[45]);
    wire[0:0] s349, in349_1, in349_2;
    wire c349;
    assign in349_1 = {pp70[41]};
    assign in349_2 = {pp71[40]};
    Full_Adder FA_349(s349, c349, in349_1, in349_2, pp69[42]);
    wire[0:0] s350, in350_1, in350_2;
    wire c350;
    assign in350_1 = {pp73[38]};
    assign in350_2 = {pp74[37]};
    Full_Adder FA_350(s350, c350, in350_1, in350_2, pp72[39]);
    wire[0:0] s351, in351_1, in351_2;
    wire c351;
    assign in351_1 = {pp75[36]};
    assign in351_2 = {pp76[35]};
    Half_Adder HA_351(s351, c351, in351_1, in351_2);
    wire[0:0] s352, in352_1, in352_2;
    wire c352;
    assign in352_1 = {pp1[111]};
    assign in352_2 = {pp2[110]};
    Full_Adder FA_352(s352, c352, in352_1, in352_2, pp0[112]);
    wire[0:0] s353, in353_1, in353_2;
    wire c353;
    assign in353_1 = {pp4[108]};
    assign in353_2 = {pp5[107]};
    Full_Adder FA_353(s353, c353, in353_1, in353_2, pp3[109]);
    wire[0:0] s354, in354_1, in354_2;
    wire c354;
    assign in354_1 = {pp7[105]};
    assign in354_2 = {pp8[104]};
    Full_Adder FA_354(s354, c354, in354_1, in354_2, pp6[106]);
    wire[0:0] s355, in355_1, in355_2;
    wire c355;
    assign in355_1 = {pp10[102]};
    assign in355_2 = {pp11[101]};
    Full_Adder FA_355(s355, c355, in355_1, in355_2, pp9[103]);
    wire[0:0] s356, in356_1, in356_2;
    wire c356;
    assign in356_1 = {pp13[99]};
    assign in356_2 = {pp14[98]};
    Full_Adder FA_356(s356, c356, in356_1, in356_2, pp12[100]);
    wire[0:0] s357, in357_1, in357_2;
    wire c357;
    assign in357_1 = {pp16[96]};
    assign in357_2 = {pp17[95]};
    Full_Adder FA_357(s357, c357, in357_1, in357_2, pp15[97]);
    wire[0:0] s358, in358_1, in358_2;
    wire c358;
    assign in358_1 = {pp19[93]};
    assign in358_2 = {pp20[92]};
    Full_Adder FA_358(s358, c358, in358_1, in358_2, pp18[94]);
    wire[0:0] s359, in359_1, in359_2;
    wire c359;
    assign in359_1 = {pp22[90]};
    assign in359_2 = {pp23[89]};
    Full_Adder FA_359(s359, c359, in359_1, in359_2, pp21[91]);
    wire[0:0] s360, in360_1, in360_2;
    wire c360;
    assign in360_1 = {pp25[87]};
    assign in360_2 = {pp26[86]};
    Full_Adder FA_360(s360, c360, in360_1, in360_2, pp24[88]);
    wire[0:0] s361, in361_1, in361_2;
    wire c361;
    assign in361_1 = {pp28[84]};
    assign in361_2 = {pp29[83]};
    Full_Adder FA_361(s361, c361, in361_1, in361_2, pp27[85]);
    wire[0:0] s362, in362_1, in362_2;
    wire c362;
    assign in362_1 = {pp31[81]};
    assign in362_2 = {pp32[80]};
    Full_Adder FA_362(s362, c362, in362_1, in362_2, pp30[82]);
    wire[0:0] s363, in363_1, in363_2;
    wire c363;
    assign in363_1 = {pp34[78]};
    assign in363_2 = {pp35[77]};
    Full_Adder FA_363(s363, c363, in363_1, in363_2, pp33[79]);
    wire[0:0] s364, in364_1, in364_2;
    wire c364;
    assign in364_1 = {pp37[75]};
    assign in364_2 = {pp38[74]};
    Full_Adder FA_364(s364, c364, in364_1, in364_2, pp36[76]);
    wire[0:0] s365, in365_1, in365_2;
    wire c365;
    assign in365_1 = {pp40[72]};
    assign in365_2 = {pp41[71]};
    Full_Adder FA_365(s365, c365, in365_1, in365_2, pp39[73]);
    wire[0:0] s366, in366_1, in366_2;
    wire c366;
    assign in366_1 = {pp43[69]};
    assign in366_2 = {pp44[68]};
    Full_Adder FA_366(s366, c366, in366_1, in366_2, pp42[70]);
    wire[0:0] s367, in367_1, in367_2;
    wire c367;
    assign in367_1 = {pp46[66]};
    assign in367_2 = {pp47[65]};
    Full_Adder FA_367(s367, c367, in367_1, in367_2, pp45[67]);
    wire[0:0] s368, in368_1, in368_2;
    wire c368;
    assign in368_1 = {pp49[63]};
    assign in368_2 = {pp50[62]};
    Full_Adder FA_368(s368, c368, in368_1, in368_2, pp48[64]);
    wire[0:0] s369, in369_1, in369_2;
    wire c369;
    assign in369_1 = {pp52[60]};
    assign in369_2 = {pp53[59]};
    Full_Adder FA_369(s369, c369, in369_1, in369_2, pp51[61]);
    wire[0:0] s370, in370_1, in370_2;
    wire c370;
    assign in370_1 = {pp55[57]};
    assign in370_2 = {pp56[56]};
    Full_Adder FA_370(s370, c370, in370_1, in370_2, pp54[58]);
    wire[0:0] s371, in371_1, in371_2;
    wire c371;
    assign in371_1 = {pp58[54]};
    assign in371_2 = {pp59[53]};
    Full_Adder FA_371(s371, c371, in371_1, in371_2, pp57[55]);
    wire[0:0] s372, in372_1, in372_2;
    wire c372;
    assign in372_1 = {pp61[51]};
    assign in372_2 = {pp62[50]};
    Full_Adder FA_372(s372, c372, in372_1, in372_2, pp60[52]);
    wire[0:0] s373, in373_1, in373_2;
    wire c373;
    assign in373_1 = {pp64[48]};
    assign in373_2 = {pp65[47]};
    Full_Adder FA_373(s373, c373, in373_1, in373_2, pp63[49]);
    wire[0:0] s374, in374_1, in374_2;
    wire c374;
    assign in374_1 = {pp67[45]};
    assign in374_2 = {pp68[44]};
    Full_Adder FA_374(s374, c374, in374_1, in374_2, pp66[46]);
    wire[0:0] s375, in375_1, in375_2;
    wire c375;
    assign in375_1 = {pp70[42]};
    assign in375_2 = {pp71[41]};
    Full_Adder FA_375(s375, c375, in375_1, in375_2, pp69[43]);
    wire[0:0] s376, in376_1, in376_2;
    wire c376;
    assign in376_1 = {pp73[39]};
    assign in376_2 = {pp74[38]};
    Full_Adder FA_376(s376, c376, in376_1, in376_2, pp72[40]);
    wire[0:0] s377, in377_1, in377_2;
    wire c377;
    assign in377_1 = {pp76[36]};
    assign in377_2 = {pp77[35]};
    Full_Adder FA_377(s377, c377, in377_1, in377_2, pp75[37]);
    wire[0:0] s378, in378_1, in378_2;
    wire c378;
    assign in378_1 = {pp78[34]};
    assign in378_2 = {pp79[33]};
    Half_Adder HA_378(s378, c378, in378_1, in378_2);
    wire[0:0] s379, in379_1, in379_2;
    wire c379;
    assign in379_1 = {pp1[112]};
    assign in379_2 = {pp2[111]};
    Full_Adder FA_379(s379, c379, in379_1, in379_2, pp0[113]);
    wire[0:0] s380, in380_1, in380_2;
    wire c380;
    assign in380_1 = {pp4[109]};
    assign in380_2 = {pp5[108]};
    Full_Adder FA_380(s380, c380, in380_1, in380_2, pp3[110]);
    wire[0:0] s381, in381_1, in381_2;
    wire c381;
    assign in381_1 = {pp7[106]};
    assign in381_2 = {pp8[105]};
    Full_Adder FA_381(s381, c381, in381_1, in381_2, pp6[107]);
    wire[0:0] s382, in382_1, in382_2;
    wire c382;
    assign in382_1 = {pp10[103]};
    assign in382_2 = {pp11[102]};
    Full_Adder FA_382(s382, c382, in382_1, in382_2, pp9[104]);
    wire[0:0] s383, in383_1, in383_2;
    wire c383;
    assign in383_1 = {pp13[100]};
    assign in383_2 = {pp14[99]};
    Full_Adder FA_383(s383, c383, in383_1, in383_2, pp12[101]);
    wire[0:0] s384, in384_1, in384_2;
    wire c384;
    assign in384_1 = {pp16[97]};
    assign in384_2 = {pp17[96]};
    Full_Adder FA_384(s384, c384, in384_1, in384_2, pp15[98]);
    wire[0:0] s385, in385_1, in385_2;
    wire c385;
    assign in385_1 = {pp19[94]};
    assign in385_2 = {pp20[93]};
    Full_Adder FA_385(s385, c385, in385_1, in385_2, pp18[95]);
    wire[0:0] s386, in386_1, in386_2;
    wire c386;
    assign in386_1 = {pp22[91]};
    assign in386_2 = {pp23[90]};
    Full_Adder FA_386(s386, c386, in386_1, in386_2, pp21[92]);
    wire[0:0] s387, in387_1, in387_2;
    wire c387;
    assign in387_1 = {pp25[88]};
    assign in387_2 = {pp26[87]};
    Full_Adder FA_387(s387, c387, in387_1, in387_2, pp24[89]);
    wire[0:0] s388, in388_1, in388_2;
    wire c388;
    assign in388_1 = {pp28[85]};
    assign in388_2 = {pp29[84]};
    Full_Adder FA_388(s388, c388, in388_1, in388_2, pp27[86]);
    wire[0:0] s389, in389_1, in389_2;
    wire c389;
    assign in389_1 = {pp31[82]};
    assign in389_2 = {pp32[81]};
    Full_Adder FA_389(s389, c389, in389_1, in389_2, pp30[83]);
    wire[0:0] s390, in390_1, in390_2;
    wire c390;
    assign in390_1 = {pp34[79]};
    assign in390_2 = {pp35[78]};
    Full_Adder FA_390(s390, c390, in390_1, in390_2, pp33[80]);
    wire[0:0] s391, in391_1, in391_2;
    wire c391;
    assign in391_1 = {pp37[76]};
    assign in391_2 = {pp38[75]};
    Full_Adder FA_391(s391, c391, in391_1, in391_2, pp36[77]);
    wire[0:0] s392, in392_1, in392_2;
    wire c392;
    assign in392_1 = {pp40[73]};
    assign in392_2 = {pp41[72]};
    Full_Adder FA_392(s392, c392, in392_1, in392_2, pp39[74]);
    wire[0:0] s393, in393_1, in393_2;
    wire c393;
    assign in393_1 = {pp43[70]};
    assign in393_2 = {pp44[69]};
    Full_Adder FA_393(s393, c393, in393_1, in393_2, pp42[71]);
    wire[0:0] s394, in394_1, in394_2;
    wire c394;
    assign in394_1 = {pp46[67]};
    assign in394_2 = {pp47[66]};
    Full_Adder FA_394(s394, c394, in394_1, in394_2, pp45[68]);
    wire[0:0] s395, in395_1, in395_2;
    wire c395;
    assign in395_1 = {pp49[64]};
    assign in395_2 = {pp50[63]};
    Full_Adder FA_395(s395, c395, in395_1, in395_2, pp48[65]);
    wire[0:0] s396, in396_1, in396_2;
    wire c396;
    assign in396_1 = {pp52[61]};
    assign in396_2 = {pp53[60]};
    Full_Adder FA_396(s396, c396, in396_1, in396_2, pp51[62]);
    wire[0:0] s397, in397_1, in397_2;
    wire c397;
    assign in397_1 = {pp55[58]};
    assign in397_2 = {pp56[57]};
    Full_Adder FA_397(s397, c397, in397_1, in397_2, pp54[59]);
    wire[0:0] s398, in398_1, in398_2;
    wire c398;
    assign in398_1 = {pp58[55]};
    assign in398_2 = {pp59[54]};
    Full_Adder FA_398(s398, c398, in398_1, in398_2, pp57[56]);
    wire[0:0] s399, in399_1, in399_2;
    wire c399;
    assign in399_1 = {pp61[52]};
    assign in399_2 = {pp62[51]};
    Full_Adder FA_399(s399, c399, in399_1, in399_2, pp60[53]);
    wire[0:0] s400, in400_1, in400_2;
    wire c400;
    assign in400_1 = {pp64[49]};
    assign in400_2 = {pp65[48]};
    Full_Adder FA_400(s400, c400, in400_1, in400_2, pp63[50]);
    wire[0:0] s401, in401_1, in401_2;
    wire c401;
    assign in401_1 = {pp67[46]};
    assign in401_2 = {pp68[45]};
    Full_Adder FA_401(s401, c401, in401_1, in401_2, pp66[47]);
    wire[0:0] s402, in402_1, in402_2;
    wire c402;
    assign in402_1 = {pp70[43]};
    assign in402_2 = {pp71[42]};
    Full_Adder FA_402(s402, c402, in402_1, in402_2, pp69[44]);
    wire[0:0] s403, in403_1, in403_2;
    wire c403;
    assign in403_1 = {pp73[40]};
    assign in403_2 = {pp74[39]};
    Full_Adder FA_403(s403, c403, in403_1, in403_2, pp72[41]);
    wire[0:0] s404, in404_1, in404_2;
    wire c404;
    assign in404_1 = {pp76[37]};
    assign in404_2 = {pp77[36]};
    Full_Adder FA_404(s404, c404, in404_1, in404_2, pp75[38]);
    wire[0:0] s405, in405_1, in405_2;
    wire c405;
    assign in405_1 = {pp79[34]};
    assign in405_2 = {pp80[33]};
    Full_Adder FA_405(s405, c405, in405_1, in405_2, pp78[35]);
    wire[0:0] s406, in406_1, in406_2;
    wire c406;
    assign in406_1 = {pp81[32]};
    assign in406_2 = {pp82[31]};
    Half_Adder HA_406(s406, c406, in406_1, in406_2);
    wire[0:0] s407, in407_1, in407_2;
    wire c407;
    assign in407_1 = {pp1[113]};
    assign in407_2 = {pp2[112]};
    Full_Adder FA_407(s407, c407, in407_1, in407_2, pp0[114]);
    wire[0:0] s408, in408_1, in408_2;
    wire c408;
    assign in408_1 = {pp4[110]};
    assign in408_2 = {pp5[109]};
    Full_Adder FA_408(s408, c408, in408_1, in408_2, pp3[111]);
    wire[0:0] s409, in409_1, in409_2;
    wire c409;
    assign in409_1 = {pp7[107]};
    assign in409_2 = {pp8[106]};
    Full_Adder FA_409(s409, c409, in409_1, in409_2, pp6[108]);
    wire[0:0] s410, in410_1, in410_2;
    wire c410;
    assign in410_1 = {pp10[104]};
    assign in410_2 = {pp11[103]};
    Full_Adder FA_410(s410, c410, in410_1, in410_2, pp9[105]);
    wire[0:0] s411, in411_1, in411_2;
    wire c411;
    assign in411_1 = {pp13[101]};
    assign in411_2 = {pp14[100]};
    Full_Adder FA_411(s411, c411, in411_1, in411_2, pp12[102]);
    wire[0:0] s412, in412_1, in412_2;
    wire c412;
    assign in412_1 = {pp16[98]};
    assign in412_2 = {pp17[97]};
    Full_Adder FA_412(s412, c412, in412_1, in412_2, pp15[99]);
    wire[0:0] s413, in413_1, in413_2;
    wire c413;
    assign in413_1 = {pp19[95]};
    assign in413_2 = {pp20[94]};
    Full_Adder FA_413(s413, c413, in413_1, in413_2, pp18[96]);
    wire[0:0] s414, in414_1, in414_2;
    wire c414;
    assign in414_1 = {pp22[92]};
    assign in414_2 = {pp23[91]};
    Full_Adder FA_414(s414, c414, in414_1, in414_2, pp21[93]);
    wire[0:0] s415, in415_1, in415_2;
    wire c415;
    assign in415_1 = {pp25[89]};
    assign in415_2 = {pp26[88]};
    Full_Adder FA_415(s415, c415, in415_1, in415_2, pp24[90]);
    wire[0:0] s416, in416_1, in416_2;
    wire c416;
    assign in416_1 = {pp28[86]};
    assign in416_2 = {pp29[85]};
    Full_Adder FA_416(s416, c416, in416_1, in416_2, pp27[87]);
    wire[0:0] s417, in417_1, in417_2;
    wire c417;
    assign in417_1 = {pp31[83]};
    assign in417_2 = {pp32[82]};
    Full_Adder FA_417(s417, c417, in417_1, in417_2, pp30[84]);
    wire[0:0] s418, in418_1, in418_2;
    wire c418;
    assign in418_1 = {pp34[80]};
    assign in418_2 = {pp35[79]};
    Full_Adder FA_418(s418, c418, in418_1, in418_2, pp33[81]);
    wire[0:0] s419, in419_1, in419_2;
    wire c419;
    assign in419_1 = {pp37[77]};
    assign in419_2 = {pp38[76]};
    Full_Adder FA_419(s419, c419, in419_1, in419_2, pp36[78]);
    wire[0:0] s420, in420_1, in420_2;
    wire c420;
    assign in420_1 = {pp40[74]};
    assign in420_2 = {pp41[73]};
    Full_Adder FA_420(s420, c420, in420_1, in420_2, pp39[75]);
    wire[0:0] s421, in421_1, in421_2;
    wire c421;
    assign in421_1 = {pp43[71]};
    assign in421_2 = {pp44[70]};
    Full_Adder FA_421(s421, c421, in421_1, in421_2, pp42[72]);
    wire[0:0] s422, in422_1, in422_2;
    wire c422;
    assign in422_1 = {pp46[68]};
    assign in422_2 = {pp47[67]};
    Full_Adder FA_422(s422, c422, in422_1, in422_2, pp45[69]);
    wire[0:0] s423, in423_1, in423_2;
    wire c423;
    assign in423_1 = {pp49[65]};
    assign in423_2 = {pp50[64]};
    Full_Adder FA_423(s423, c423, in423_1, in423_2, pp48[66]);
    wire[0:0] s424, in424_1, in424_2;
    wire c424;
    assign in424_1 = {pp52[62]};
    assign in424_2 = {pp53[61]};
    Full_Adder FA_424(s424, c424, in424_1, in424_2, pp51[63]);
    wire[0:0] s425, in425_1, in425_2;
    wire c425;
    assign in425_1 = {pp55[59]};
    assign in425_2 = {pp56[58]};
    Full_Adder FA_425(s425, c425, in425_1, in425_2, pp54[60]);
    wire[0:0] s426, in426_1, in426_2;
    wire c426;
    assign in426_1 = {pp58[56]};
    assign in426_2 = {pp59[55]};
    Full_Adder FA_426(s426, c426, in426_1, in426_2, pp57[57]);
    wire[0:0] s427, in427_1, in427_2;
    wire c427;
    assign in427_1 = {pp61[53]};
    assign in427_2 = {pp62[52]};
    Full_Adder FA_427(s427, c427, in427_1, in427_2, pp60[54]);
    wire[0:0] s428, in428_1, in428_2;
    wire c428;
    assign in428_1 = {pp64[50]};
    assign in428_2 = {pp65[49]};
    Full_Adder FA_428(s428, c428, in428_1, in428_2, pp63[51]);
    wire[0:0] s429, in429_1, in429_2;
    wire c429;
    assign in429_1 = {pp67[47]};
    assign in429_2 = {pp68[46]};
    Full_Adder FA_429(s429, c429, in429_1, in429_2, pp66[48]);
    wire[0:0] s430, in430_1, in430_2;
    wire c430;
    assign in430_1 = {pp70[44]};
    assign in430_2 = {pp71[43]};
    Full_Adder FA_430(s430, c430, in430_1, in430_2, pp69[45]);
    wire[0:0] s431, in431_1, in431_2;
    wire c431;
    assign in431_1 = {pp73[41]};
    assign in431_2 = {pp74[40]};
    Full_Adder FA_431(s431, c431, in431_1, in431_2, pp72[42]);
    wire[0:0] s432, in432_1, in432_2;
    wire c432;
    assign in432_1 = {pp76[38]};
    assign in432_2 = {pp77[37]};
    Full_Adder FA_432(s432, c432, in432_1, in432_2, pp75[39]);
    wire[0:0] s433, in433_1, in433_2;
    wire c433;
    assign in433_1 = {pp79[35]};
    assign in433_2 = {pp80[34]};
    Full_Adder FA_433(s433, c433, in433_1, in433_2, pp78[36]);
    wire[0:0] s434, in434_1, in434_2;
    wire c434;
    assign in434_1 = {pp82[32]};
    assign in434_2 = {pp83[31]};
    Full_Adder FA_434(s434, c434, in434_1, in434_2, pp81[33]);
    wire[0:0] s435, in435_1, in435_2;
    wire c435;
    assign in435_1 = {pp84[30]};
    assign in435_2 = {pp85[29]};
    Half_Adder HA_435(s435, c435, in435_1, in435_2);
    wire[0:0] s436, in436_1, in436_2;
    wire c436;
    assign in436_1 = {pp1[114]};
    assign in436_2 = {pp2[113]};
    Full_Adder FA_436(s436, c436, in436_1, in436_2, pp0[115]);
    wire[0:0] s437, in437_1, in437_2;
    wire c437;
    assign in437_1 = {pp4[111]};
    assign in437_2 = {pp5[110]};
    Full_Adder FA_437(s437, c437, in437_1, in437_2, pp3[112]);
    wire[0:0] s438, in438_1, in438_2;
    wire c438;
    assign in438_1 = {pp7[108]};
    assign in438_2 = {pp8[107]};
    Full_Adder FA_438(s438, c438, in438_1, in438_2, pp6[109]);
    wire[0:0] s439, in439_1, in439_2;
    wire c439;
    assign in439_1 = {pp10[105]};
    assign in439_2 = {pp11[104]};
    Full_Adder FA_439(s439, c439, in439_1, in439_2, pp9[106]);
    wire[0:0] s440, in440_1, in440_2;
    wire c440;
    assign in440_1 = {pp13[102]};
    assign in440_2 = {pp14[101]};
    Full_Adder FA_440(s440, c440, in440_1, in440_2, pp12[103]);
    wire[0:0] s441, in441_1, in441_2;
    wire c441;
    assign in441_1 = {pp16[99]};
    assign in441_2 = {pp17[98]};
    Full_Adder FA_441(s441, c441, in441_1, in441_2, pp15[100]);
    wire[0:0] s442, in442_1, in442_2;
    wire c442;
    assign in442_1 = {pp19[96]};
    assign in442_2 = {pp20[95]};
    Full_Adder FA_442(s442, c442, in442_1, in442_2, pp18[97]);
    wire[0:0] s443, in443_1, in443_2;
    wire c443;
    assign in443_1 = {pp22[93]};
    assign in443_2 = {pp23[92]};
    Full_Adder FA_443(s443, c443, in443_1, in443_2, pp21[94]);
    wire[0:0] s444, in444_1, in444_2;
    wire c444;
    assign in444_1 = {pp25[90]};
    assign in444_2 = {pp26[89]};
    Full_Adder FA_444(s444, c444, in444_1, in444_2, pp24[91]);
    wire[0:0] s445, in445_1, in445_2;
    wire c445;
    assign in445_1 = {pp28[87]};
    assign in445_2 = {pp29[86]};
    Full_Adder FA_445(s445, c445, in445_1, in445_2, pp27[88]);
    wire[0:0] s446, in446_1, in446_2;
    wire c446;
    assign in446_1 = {pp31[84]};
    assign in446_2 = {pp32[83]};
    Full_Adder FA_446(s446, c446, in446_1, in446_2, pp30[85]);
    wire[0:0] s447, in447_1, in447_2;
    wire c447;
    assign in447_1 = {pp34[81]};
    assign in447_2 = {pp35[80]};
    Full_Adder FA_447(s447, c447, in447_1, in447_2, pp33[82]);
    wire[0:0] s448, in448_1, in448_2;
    wire c448;
    assign in448_1 = {pp37[78]};
    assign in448_2 = {pp38[77]};
    Full_Adder FA_448(s448, c448, in448_1, in448_2, pp36[79]);
    wire[0:0] s449, in449_1, in449_2;
    wire c449;
    assign in449_1 = {pp40[75]};
    assign in449_2 = {pp41[74]};
    Full_Adder FA_449(s449, c449, in449_1, in449_2, pp39[76]);
    wire[0:0] s450, in450_1, in450_2;
    wire c450;
    assign in450_1 = {pp43[72]};
    assign in450_2 = {pp44[71]};
    Full_Adder FA_450(s450, c450, in450_1, in450_2, pp42[73]);
    wire[0:0] s451, in451_1, in451_2;
    wire c451;
    assign in451_1 = {pp46[69]};
    assign in451_2 = {pp47[68]};
    Full_Adder FA_451(s451, c451, in451_1, in451_2, pp45[70]);
    wire[0:0] s452, in452_1, in452_2;
    wire c452;
    assign in452_1 = {pp49[66]};
    assign in452_2 = {pp50[65]};
    Full_Adder FA_452(s452, c452, in452_1, in452_2, pp48[67]);
    wire[0:0] s453, in453_1, in453_2;
    wire c453;
    assign in453_1 = {pp52[63]};
    assign in453_2 = {pp53[62]};
    Full_Adder FA_453(s453, c453, in453_1, in453_2, pp51[64]);
    wire[0:0] s454, in454_1, in454_2;
    wire c454;
    assign in454_1 = {pp55[60]};
    assign in454_2 = {pp56[59]};
    Full_Adder FA_454(s454, c454, in454_1, in454_2, pp54[61]);
    wire[0:0] s455, in455_1, in455_2;
    wire c455;
    assign in455_1 = {pp58[57]};
    assign in455_2 = {pp59[56]};
    Full_Adder FA_455(s455, c455, in455_1, in455_2, pp57[58]);
    wire[0:0] s456, in456_1, in456_2;
    wire c456;
    assign in456_1 = {pp61[54]};
    assign in456_2 = {pp62[53]};
    Full_Adder FA_456(s456, c456, in456_1, in456_2, pp60[55]);
    wire[0:0] s457, in457_1, in457_2;
    wire c457;
    assign in457_1 = {pp64[51]};
    assign in457_2 = {pp65[50]};
    Full_Adder FA_457(s457, c457, in457_1, in457_2, pp63[52]);
    wire[0:0] s458, in458_1, in458_2;
    wire c458;
    assign in458_1 = {pp67[48]};
    assign in458_2 = {pp68[47]};
    Full_Adder FA_458(s458, c458, in458_1, in458_2, pp66[49]);
    wire[0:0] s459, in459_1, in459_2;
    wire c459;
    assign in459_1 = {pp70[45]};
    assign in459_2 = {pp71[44]};
    Full_Adder FA_459(s459, c459, in459_1, in459_2, pp69[46]);
    wire[0:0] s460, in460_1, in460_2;
    wire c460;
    assign in460_1 = {pp73[42]};
    assign in460_2 = {pp74[41]};
    Full_Adder FA_460(s460, c460, in460_1, in460_2, pp72[43]);
    wire[0:0] s461, in461_1, in461_2;
    wire c461;
    assign in461_1 = {pp76[39]};
    assign in461_2 = {pp77[38]};
    Full_Adder FA_461(s461, c461, in461_1, in461_2, pp75[40]);
    wire[0:0] s462, in462_1, in462_2;
    wire c462;
    assign in462_1 = {pp79[36]};
    assign in462_2 = {pp80[35]};
    Full_Adder FA_462(s462, c462, in462_1, in462_2, pp78[37]);
    wire[0:0] s463, in463_1, in463_2;
    wire c463;
    assign in463_1 = {pp82[33]};
    assign in463_2 = {pp83[32]};
    Full_Adder FA_463(s463, c463, in463_1, in463_2, pp81[34]);
    wire[0:0] s464, in464_1, in464_2;
    wire c464;
    assign in464_1 = {pp85[30]};
    assign in464_2 = {pp86[29]};
    Full_Adder FA_464(s464, c464, in464_1, in464_2, pp84[31]);
    wire[0:0] s465, in465_1, in465_2;
    wire c465;
    assign in465_1 = {pp87[28]};
    assign in465_2 = {pp88[27]};
    Half_Adder HA_465(s465, c465, in465_1, in465_2);
    wire[0:0] s466, in466_1, in466_2;
    wire c466;
    assign in466_1 = {pp1[115]};
    assign in466_2 = {pp2[114]};
    Full_Adder FA_466(s466, c466, in466_1, in466_2, pp0[116]);
    wire[0:0] s467, in467_1, in467_2;
    wire c467;
    assign in467_1 = {pp4[112]};
    assign in467_2 = {pp5[111]};
    Full_Adder FA_467(s467, c467, in467_1, in467_2, pp3[113]);
    wire[0:0] s468, in468_1, in468_2;
    wire c468;
    assign in468_1 = {pp7[109]};
    assign in468_2 = {pp8[108]};
    Full_Adder FA_468(s468, c468, in468_1, in468_2, pp6[110]);
    wire[0:0] s469, in469_1, in469_2;
    wire c469;
    assign in469_1 = {pp10[106]};
    assign in469_2 = {pp11[105]};
    Full_Adder FA_469(s469, c469, in469_1, in469_2, pp9[107]);
    wire[0:0] s470, in470_1, in470_2;
    wire c470;
    assign in470_1 = {pp13[103]};
    assign in470_2 = {pp14[102]};
    Full_Adder FA_470(s470, c470, in470_1, in470_2, pp12[104]);
    wire[0:0] s471, in471_1, in471_2;
    wire c471;
    assign in471_1 = {pp16[100]};
    assign in471_2 = {pp17[99]};
    Full_Adder FA_471(s471, c471, in471_1, in471_2, pp15[101]);
    wire[0:0] s472, in472_1, in472_2;
    wire c472;
    assign in472_1 = {pp19[97]};
    assign in472_2 = {pp20[96]};
    Full_Adder FA_472(s472, c472, in472_1, in472_2, pp18[98]);
    wire[0:0] s473, in473_1, in473_2;
    wire c473;
    assign in473_1 = {pp22[94]};
    assign in473_2 = {pp23[93]};
    Full_Adder FA_473(s473, c473, in473_1, in473_2, pp21[95]);
    wire[0:0] s474, in474_1, in474_2;
    wire c474;
    assign in474_1 = {pp25[91]};
    assign in474_2 = {pp26[90]};
    Full_Adder FA_474(s474, c474, in474_1, in474_2, pp24[92]);
    wire[0:0] s475, in475_1, in475_2;
    wire c475;
    assign in475_1 = {pp28[88]};
    assign in475_2 = {pp29[87]};
    Full_Adder FA_475(s475, c475, in475_1, in475_2, pp27[89]);
    wire[0:0] s476, in476_1, in476_2;
    wire c476;
    assign in476_1 = {pp31[85]};
    assign in476_2 = {pp32[84]};
    Full_Adder FA_476(s476, c476, in476_1, in476_2, pp30[86]);
    wire[0:0] s477, in477_1, in477_2;
    wire c477;
    assign in477_1 = {pp34[82]};
    assign in477_2 = {pp35[81]};
    Full_Adder FA_477(s477, c477, in477_1, in477_2, pp33[83]);
    wire[0:0] s478, in478_1, in478_2;
    wire c478;
    assign in478_1 = {pp37[79]};
    assign in478_2 = {pp38[78]};
    Full_Adder FA_478(s478, c478, in478_1, in478_2, pp36[80]);
    wire[0:0] s479, in479_1, in479_2;
    wire c479;
    assign in479_1 = {pp40[76]};
    assign in479_2 = {pp41[75]};
    Full_Adder FA_479(s479, c479, in479_1, in479_2, pp39[77]);
    wire[0:0] s480, in480_1, in480_2;
    wire c480;
    assign in480_1 = {pp43[73]};
    assign in480_2 = {pp44[72]};
    Full_Adder FA_480(s480, c480, in480_1, in480_2, pp42[74]);
    wire[0:0] s481, in481_1, in481_2;
    wire c481;
    assign in481_1 = {pp46[70]};
    assign in481_2 = {pp47[69]};
    Full_Adder FA_481(s481, c481, in481_1, in481_2, pp45[71]);
    wire[0:0] s482, in482_1, in482_2;
    wire c482;
    assign in482_1 = {pp49[67]};
    assign in482_2 = {pp50[66]};
    Full_Adder FA_482(s482, c482, in482_1, in482_2, pp48[68]);
    wire[0:0] s483, in483_1, in483_2;
    wire c483;
    assign in483_1 = {pp52[64]};
    assign in483_2 = {pp53[63]};
    Full_Adder FA_483(s483, c483, in483_1, in483_2, pp51[65]);
    wire[0:0] s484, in484_1, in484_2;
    wire c484;
    assign in484_1 = {pp55[61]};
    assign in484_2 = {pp56[60]};
    Full_Adder FA_484(s484, c484, in484_1, in484_2, pp54[62]);
    wire[0:0] s485, in485_1, in485_2;
    wire c485;
    assign in485_1 = {pp58[58]};
    assign in485_2 = {pp59[57]};
    Full_Adder FA_485(s485, c485, in485_1, in485_2, pp57[59]);
    wire[0:0] s486, in486_1, in486_2;
    wire c486;
    assign in486_1 = {pp61[55]};
    assign in486_2 = {pp62[54]};
    Full_Adder FA_486(s486, c486, in486_1, in486_2, pp60[56]);
    wire[0:0] s487, in487_1, in487_2;
    wire c487;
    assign in487_1 = {pp64[52]};
    assign in487_2 = {pp65[51]};
    Full_Adder FA_487(s487, c487, in487_1, in487_2, pp63[53]);
    wire[0:0] s488, in488_1, in488_2;
    wire c488;
    assign in488_1 = {pp67[49]};
    assign in488_2 = {pp68[48]};
    Full_Adder FA_488(s488, c488, in488_1, in488_2, pp66[50]);
    wire[0:0] s489, in489_1, in489_2;
    wire c489;
    assign in489_1 = {pp70[46]};
    assign in489_2 = {pp71[45]};
    Full_Adder FA_489(s489, c489, in489_1, in489_2, pp69[47]);
    wire[0:0] s490, in490_1, in490_2;
    wire c490;
    assign in490_1 = {pp73[43]};
    assign in490_2 = {pp74[42]};
    Full_Adder FA_490(s490, c490, in490_1, in490_2, pp72[44]);
    wire[0:0] s491, in491_1, in491_2;
    wire c491;
    assign in491_1 = {pp76[40]};
    assign in491_2 = {pp77[39]};
    Full_Adder FA_491(s491, c491, in491_1, in491_2, pp75[41]);
    wire[0:0] s492, in492_1, in492_2;
    wire c492;
    assign in492_1 = {pp79[37]};
    assign in492_2 = {pp80[36]};
    Full_Adder FA_492(s492, c492, in492_1, in492_2, pp78[38]);
    wire[0:0] s493, in493_1, in493_2;
    wire c493;
    assign in493_1 = {pp82[34]};
    assign in493_2 = {pp83[33]};
    Full_Adder FA_493(s493, c493, in493_1, in493_2, pp81[35]);
    wire[0:0] s494, in494_1, in494_2;
    wire c494;
    assign in494_1 = {pp85[31]};
    assign in494_2 = {pp86[30]};
    Full_Adder FA_494(s494, c494, in494_1, in494_2, pp84[32]);
    wire[0:0] s495, in495_1, in495_2;
    wire c495;
    assign in495_1 = {pp88[28]};
    assign in495_2 = {pp89[27]};
    Full_Adder FA_495(s495, c495, in495_1, in495_2, pp87[29]);
    wire[0:0] s496, in496_1, in496_2;
    wire c496;
    assign in496_1 = {pp90[26]};
    assign in496_2 = {pp91[25]};
    Half_Adder HA_496(s496, c496, in496_1, in496_2);
    wire[0:0] s497, in497_1, in497_2;
    wire c497;
    assign in497_1 = {pp1[116]};
    assign in497_2 = {pp2[115]};
    Full_Adder FA_497(s497, c497, in497_1, in497_2, pp0[117]);
    wire[0:0] s498, in498_1, in498_2;
    wire c498;
    assign in498_1 = {pp4[113]};
    assign in498_2 = {pp5[112]};
    Full_Adder FA_498(s498, c498, in498_1, in498_2, pp3[114]);
    wire[0:0] s499, in499_1, in499_2;
    wire c499;
    assign in499_1 = {pp7[110]};
    assign in499_2 = {pp8[109]};
    Full_Adder FA_499(s499, c499, in499_1, in499_2, pp6[111]);
    wire[0:0] s500, in500_1, in500_2;
    wire c500;
    assign in500_1 = {pp10[107]};
    assign in500_2 = {pp11[106]};
    Full_Adder FA_500(s500, c500, in500_1, in500_2, pp9[108]);
    wire[0:0] s501, in501_1, in501_2;
    wire c501;
    assign in501_1 = {pp13[104]};
    assign in501_2 = {pp14[103]};
    Full_Adder FA_501(s501, c501, in501_1, in501_2, pp12[105]);
    wire[0:0] s502, in502_1, in502_2;
    wire c502;
    assign in502_1 = {pp16[101]};
    assign in502_2 = {pp17[100]};
    Full_Adder FA_502(s502, c502, in502_1, in502_2, pp15[102]);
    wire[0:0] s503, in503_1, in503_2;
    wire c503;
    assign in503_1 = {pp19[98]};
    assign in503_2 = {pp20[97]};
    Full_Adder FA_503(s503, c503, in503_1, in503_2, pp18[99]);
    wire[0:0] s504, in504_1, in504_2;
    wire c504;
    assign in504_1 = {pp22[95]};
    assign in504_2 = {pp23[94]};
    Full_Adder FA_504(s504, c504, in504_1, in504_2, pp21[96]);
    wire[0:0] s505, in505_1, in505_2;
    wire c505;
    assign in505_1 = {pp25[92]};
    assign in505_2 = {pp26[91]};
    Full_Adder FA_505(s505, c505, in505_1, in505_2, pp24[93]);
    wire[0:0] s506, in506_1, in506_2;
    wire c506;
    assign in506_1 = {pp28[89]};
    assign in506_2 = {pp29[88]};
    Full_Adder FA_506(s506, c506, in506_1, in506_2, pp27[90]);
    wire[0:0] s507, in507_1, in507_2;
    wire c507;
    assign in507_1 = {pp31[86]};
    assign in507_2 = {pp32[85]};
    Full_Adder FA_507(s507, c507, in507_1, in507_2, pp30[87]);
    wire[0:0] s508, in508_1, in508_2;
    wire c508;
    assign in508_1 = {pp34[83]};
    assign in508_2 = {pp35[82]};
    Full_Adder FA_508(s508, c508, in508_1, in508_2, pp33[84]);
    wire[0:0] s509, in509_1, in509_2;
    wire c509;
    assign in509_1 = {pp37[80]};
    assign in509_2 = {pp38[79]};
    Full_Adder FA_509(s509, c509, in509_1, in509_2, pp36[81]);
    wire[0:0] s510, in510_1, in510_2;
    wire c510;
    assign in510_1 = {pp40[77]};
    assign in510_2 = {pp41[76]};
    Full_Adder FA_510(s510, c510, in510_1, in510_2, pp39[78]);
    wire[0:0] s511, in511_1, in511_2;
    wire c511;
    assign in511_1 = {pp43[74]};
    assign in511_2 = {pp44[73]};
    Full_Adder FA_511(s511, c511, in511_1, in511_2, pp42[75]);
    wire[0:0] s512, in512_1, in512_2;
    wire c512;
    assign in512_1 = {pp46[71]};
    assign in512_2 = {pp47[70]};
    Full_Adder FA_512(s512, c512, in512_1, in512_2, pp45[72]);
    wire[0:0] s513, in513_1, in513_2;
    wire c513;
    assign in513_1 = {pp49[68]};
    assign in513_2 = {pp50[67]};
    Full_Adder FA_513(s513, c513, in513_1, in513_2, pp48[69]);
    wire[0:0] s514, in514_1, in514_2;
    wire c514;
    assign in514_1 = {pp52[65]};
    assign in514_2 = {pp53[64]};
    Full_Adder FA_514(s514, c514, in514_1, in514_2, pp51[66]);
    wire[0:0] s515, in515_1, in515_2;
    wire c515;
    assign in515_1 = {pp55[62]};
    assign in515_2 = {pp56[61]};
    Full_Adder FA_515(s515, c515, in515_1, in515_2, pp54[63]);
    wire[0:0] s516, in516_1, in516_2;
    wire c516;
    assign in516_1 = {pp58[59]};
    assign in516_2 = {pp59[58]};
    Full_Adder FA_516(s516, c516, in516_1, in516_2, pp57[60]);
    wire[0:0] s517, in517_1, in517_2;
    wire c517;
    assign in517_1 = {pp61[56]};
    assign in517_2 = {pp62[55]};
    Full_Adder FA_517(s517, c517, in517_1, in517_2, pp60[57]);
    wire[0:0] s518, in518_1, in518_2;
    wire c518;
    assign in518_1 = {pp64[53]};
    assign in518_2 = {pp65[52]};
    Full_Adder FA_518(s518, c518, in518_1, in518_2, pp63[54]);
    wire[0:0] s519, in519_1, in519_2;
    wire c519;
    assign in519_1 = {pp67[50]};
    assign in519_2 = {pp68[49]};
    Full_Adder FA_519(s519, c519, in519_1, in519_2, pp66[51]);
    wire[0:0] s520, in520_1, in520_2;
    wire c520;
    assign in520_1 = {pp70[47]};
    assign in520_2 = {pp71[46]};
    Full_Adder FA_520(s520, c520, in520_1, in520_2, pp69[48]);
    wire[0:0] s521, in521_1, in521_2;
    wire c521;
    assign in521_1 = {pp73[44]};
    assign in521_2 = {pp74[43]};
    Full_Adder FA_521(s521, c521, in521_1, in521_2, pp72[45]);
    wire[0:0] s522, in522_1, in522_2;
    wire c522;
    assign in522_1 = {pp76[41]};
    assign in522_2 = {pp77[40]};
    Full_Adder FA_522(s522, c522, in522_1, in522_2, pp75[42]);
    wire[0:0] s523, in523_1, in523_2;
    wire c523;
    assign in523_1 = {pp79[38]};
    assign in523_2 = {pp80[37]};
    Full_Adder FA_523(s523, c523, in523_1, in523_2, pp78[39]);
    wire[0:0] s524, in524_1, in524_2;
    wire c524;
    assign in524_1 = {pp82[35]};
    assign in524_2 = {pp83[34]};
    Full_Adder FA_524(s524, c524, in524_1, in524_2, pp81[36]);
    wire[0:0] s525, in525_1, in525_2;
    wire c525;
    assign in525_1 = {pp85[32]};
    assign in525_2 = {pp86[31]};
    Full_Adder FA_525(s525, c525, in525_1, in525_2, pp84[33]);
    wire[0:0] s526, in526_1, in526_2;
    wire c526;
    assign in526_1 = {pp88[29]};
    assign in526_2 = {pp89[28]};
    Full_Adder FA_526(s526, c526, in526_1, in526_2, pp87[30]);
    wire[0:0] s527, in527_1, in527_2;
    wire c527;
    assign in527_1 = {pp91[26]};
    assign in527_2 = {pp92[25]};
    Full_Adder FA_527(s527, c527, in527_1, in527_2, pp90[27]);
    wire[0:0] s528, in528_1, in528_2;
    wire c528;
    assign in528_1 = {pp93[24]};
    assign in528_2 = {pp94[23]};
    Half_Adder HA_528(s528, c528, in528_1, in528_2);
    wire[0:0] s529, in529_1, in529_2;
    wire c529;
    assign in529_1 = {pp1[117]};
    assign in529_2 = {pp2[116]};
    Full_Adder FA_529(s529, c529, in529_1, in529_2, pp0[118]);
    wire[0:0] s530, in530_1, in530_2;
    wire c530;
    assign in530_1 = {pp4[114]};
    assign in530_2 = {pp5[113]};
    Full_Adder FA_530(s530, c530, in530_1, in530_2, pp3[115]);
    wire[0:0] s531, in531_1, in531_2;
    wire c531;
    assign in531_1 = {pp7[111]};
    assign in531_2 = {pp8[110]};
    Full_Adder FA_531(s531, c531, in531_1, in531_2, pp6[112]);
    wire[0:0] s532, in532_1, in532_2;
    wire c532;
    assign in532_1 = {pp10[108]};
    assign in532_2 = {pp11[107]};
    Full_Adder FA_532(s532, c532, in532_1, in532_2, pp9[109]);
    wire[0:0] s533, in533_1, in533_2;
    wire c533;
    assign in533_1 = {pp13[105]};
    assign in533_2 = {pp14[104]};
    Full_Adder FA_533(s533, c533, in533_1, in533_2, pp12[106]);
    wire[0:0] s534, in534_1, in534_2;
    wire c534;
    assign in534_1 = {pp16[102]};
    assign in534_2 = {pp17[101]};
    Full_Adder FA_534(s534, c534, in534_1, in534_2, pp15[103]);
    wire[0:0] s535, in535_1, in535_2;
    wire c535;
    assign in535_1 = {pp19[99]};
    assign in535_2 = {pp20[98]};
    Full_Adder FA_535(s535, c535, in535_1, in535_2, pp18[100]);
    wire[0:0] s536, in536_1, in536_2;
    wire c536;
    assign in536_1 = {pp22[96]};
    assign in536_2 = {pp23[95]};
    Full_Adder FA_536(s536, c536, in536_1, in536_2, pp21[97]);
    wire[0:0] s537, in537_1, in537_2;
    wire c537;
    assign in537_1 = {pp25[93]};
    assign in537_2 = {pp26[92]};
    Full_Adder FA_537(s537, c537, in537_1, in537_2, pp24[94]);
    wire[0:0] s538, in538_1, in538_2;
    wire c538;
    assign in538_1 = {pp28[90]};
    assign in538_2 = {pp29[89]};
    Full_Adder FA_538(s538, c538, in538_1, in538_2, pp27[91]);
    wire[0:0] s539, in539_1, in539_2;
    wire c539;
    assign in539_1 = {pp31[87]};
    assign in539_2 = {pp32[86]};
    Full_Adder FA_539(s539, c539, in539_1, in539_2, pp30[88]);
    wire[0:0] s540, in540_1, in540_2;
    wire c540;
    assign in540_1 = {pp34[84]};
    assign in540_2 = {pp35[83]};
    Full_Adder FA_540(s540, c540, in540_1, in540_2, pp33[85]);
    wire[0:0] s541, in541_1, in541_2;
    wire c541;
    assign in541_1 = {pp37[81]};
    assign in541_2 = {pp38[80]};
    Full_Adder FA_541(s541, c541, in541_1, in541_2, pp36[82]);
    wire[0:0] s542, in542_1, in542_2;
    wire c542;
    assign in542_1 = {pp40[78]};
    assign in542_2 = {pp41[77]};
    Full_Adder FA_542(s542, c542, in542_1, in542_2, pp39[79]);
    wire[0:0] s543, in543_1, in543_2;
    wire c543;
    assign in543_1 = {pp43[75]};
    assign in543_2 = {pp44[74]};
    Full_Adder FA_543(s543, c543, in543_1, in543_2, pp42[76]);
    wire[0:0] s544, in544_1, in544_2;
    wire c544;
    assign in544_1 = {pp46[72]};
    assign in544_2 = {pp47[71]};
    Full_Adder FA_544(s544, c544, in544_1, in544_2, pp45[73]);
    wire[0:0] s545, in545_1, in545_2;
    wire c545;
    assign in545_1 = {pp49[69]};
    assign in545_2 = {pp50[68]};
    Full_Adder FA_545(s545, c545, in545_1, in545_2, pp48[70]);
    wire[0:0] s546, in546_1, in546_2;
    wire c546;
    assign in546_1 = {pp52[66]};
    assign in546_2 = {pp53[65]};
    Full_Adder FA_546(s546, c546, in546_1, in546_2, pp51[67]);
    wire[0:0] s547, in547_1, in547_2;
    wire c547;
    assign in547_1 = {pp55[63]};
    assign in547_2 = {pp56[62]};
    Full_Adder FA_547(s547, c547, in547_1, in547_2, pp54[64]);
    wire[0:0] s548, in548_1, in548_2;
    wire c548;
    assign in548_1 = {pp58[60]};
    assign in548_2 = {pp59[59]};
    Full_Adder FA_548(s548, c548, in548_1, in548_2, pp57[61]);
    wire[0:0] s549, in549_1, in549_2;
    wire c549;
    assign in549_1 = {pp61[57]};
    assign in549_2 = {pp62[56]};
    Full_Adder FA_549(s549, c549, in549_1, in549_2, pp60[58]);
    wire[0:0] s550, in550_1, in550_2;
    wire c550;
    assign in550_1 = {pp64[54]};
    assign in550_2 = {pp65[53]};
    Full_Adder FA_550(s550, c550, in550_1, in550_2, pp63[55]);
    wire[0:0] s551, in551_1, in551_2;
    wire c551;
    assign in551_1 = {pp67[51]};
    assign in551_2 = {pp68[50]};
    Full_Adder FA_551(s551, c551, in551_1, in551_2, pp66[52]);
    wire[0:0] s552, in552_1, in552_2;
    wire c552;
    assign in552_1 = {pp70[48]};
    assign in552_2 = {pp71[47]};
    Full_Adder FA_552(s552, c552, in552_1, in552_2, pp69[49]);
    wire[0:0] s553, in553_1, in553_2;
    wire c553;
    assign in553_1 = {pp73[45]};
    assign in553_2 = {pp74[44]};
    Full_Adder FA_553(s553, c553, in553_1, in553_2, pp72[46]);
    wire[0:0] s554, in554_1, in554_2;
    wire c554;
    assign in554_1 = {pp76[42]};
    assign in554_2 = {pp77[41]};
    Full_Adder FA_554(s554, c554, in554_1, in554_2, pp75[43]);
    wire[0:0] s555, in555_1, in555_2;
    wire c555;
    assign in555_1 = {pp79[39]};
    assign in555_2 = {pp80[38]};
    Full_Adder FA_555(s555, c555, in555_1, in555_2, pp78[40]);
    wire[0:0] s556, in556_1, in556_2;
    wire c556;
    assign in556_1 = {pp82[36]};
    assign in556_2 = {pp83[35]};
    Full_Adder FA_556(s556, c556, in556_1, in556_2, pp81[37]);
    wire[0:0] s557, in557_1, in557_2;
    wire c557;
    assign in557_1 = {pp85[33]};
    assign in557_2 = {pp86[32]};
    Full_Adder FA_557(s557, c557, in557_1, in557_2, pp84[34]);
    wire[0:0] s558, in558_1, in558_2;
    wire c558;
    assign in558_1 = {pp88[30]};
    assign in558_2 = {pp89[29]};
    Full_Adder FA_558(s558, c558, in558_1, in558_2, pp87[31]);
    wire[0:0] s559, in559_1, in559_2;
    wire c559;
    assign in559_1 = {pp91[27]};
    assign in559_2 = {pp92[26]};
    Full_Adder FA_559(s559, c559, in559_1, in559_2, pp90[28]);
    wire[0:0] s560, in560_1, in560_2;
    wire c560;
    assign in560_1 = {pp94[24]};
    assign in560_2 = {pp95[23]};
    Full_Adder FA_560(s560, c560, in560_1, in560_2, pp93[25]);
    wire[0:0] s561, in561_1, in561_2;
    wire c561;
    assign in561_1 = {pp96[22]};
    assign in561_2 = {pp97[21]};
    Half_Adder HA_561(s561, c561, in561_1, in561_2);
    wire[0:0] s562, in562_1, in562_2;
    wire c562;
    assign in562_1 = {pp1[118]};
    assign in562_2 = {pp2[117]};
    Full_Adder FA_562(s562, c562, in562_1, in562_2, pp0[119]);
    wire[0:0] s563, in563_1, in563_2;
    wire c563;
    assign in563_1 = {pp4[115]};
    assign in563_2 = {pp5[114]};
    Full_Adder FA_563(s563, c563, in563_1, in563_2, pp3[116]);
    wire[0:0] s564, in564_1, in564_2;
    wire c564;
    assign in564_1 = {pp7[112]};
    assign in564_2 = {pp8[111]};
    Full_Adder FA_564(s564, c564, in564_1, in564_2, pp6[113]);
    wire[0:0] s565, in565_1, in565_2;
    wire c565;
    assign in565_1 = {pp10[109]};
    assign in565_2 = {pp11[108]};
    Full_Adder FA_565(s565, c565, in565_1, in565_2, pp9[110]);
    wire[0:0] s566, in566_1, in566_2;
    wire c566;
    assign in566_1 = {pp13[106]};
    assign in566_2 = {pp14[105]};
    Full_Adder FA_566(s566, c566, in566_1, in566_2, pp12[107]);
    wire[0:0] s567, in567_1, in567_2;
    wire c567;
    assign in567_1 = {pp16[103]};
    assign in567_2 = {pp17[102]};
    Full_Adder FA_567(s567, c567, in567_1, in567_2, pp15[104]);
    wire[0:0] s568, in568_1, in568_2;
    wire c568;
    assign in568_1 = {pp19[100]};
    assign in568_2 = {pp20[99]};
    Full_Adder FA_568(s568, c568, in568_1, in568_2, pp18[101]);
    wire[0:0] s569, in569_1, in569_2;
    wire c569;
    assign in569_1 = {pp22[97]};
    assign in569_2 = {pp23[96]};
    Full_Adder FA_569(s569, c569, in569_1, in569_2, pp21[98]);
    wire[0:0] s570, in570_1, in570_2;
    wire c570;
    assign in570_1 = {pp25[94]};
    assign in570_2 = {pp26[93]};
    Full_Adder FA_570(s570, c570, in570_1, in570_2, pp24[95]);
    wire[0:0] s571, in571_1, in571_2;
    wire c571;
    assign in571_1 = {pp28[91]};
    assign in571_2 = {pp29[90]};
    Full_Adder FA_571(s571, c571, in571_1, in571_2, pp27[92]);
    wire[0:0] s572, in572_1, in572_2;
    wire c572;
    assign in572_1 = {pp31[88]};
    assign in572_2 = {pp32[87]};
    Full_Adder FA_572(s572, c572, in572_1, in572_2, pp30[89]);
    wire[0:0] s573, in573_1, in573_2;
    wire c573;
    assign in573_1 = {pp34[85]};
    assign in573_2 = {pp35[84]};
    Full_Adder FA_573(s573, c573, in573_1, in573_2, pp33[86]);
    wire[0:0] s574, in574_1, in574_2;
    wire c574;
    assign in574_1 = {pp37[82]};
    assign in574_2 = {pp38[81]};
    Full_Adder FA_574(s574, c574, in574_1, in574_2, pp36[83]);
    wire[0:0] s575, in575_1, in575_2;
    wire c575;
    assign in575_1 = {pp40[79]};
    assign in575_2 = {pp41[78]};
    Full_Adder FA_575(s575, c575, in575_1, in575_2, pp39[80]);
    wire[0:0] s576, in576_1, in576_2;
    wire c576;
    assign in576_1 = {pp43[76]};
    assign in576_2 = {pp44[75]};
    Full_Adder FA_576(s576, c576, in576_1, in576_2, pp42[77]);
    wire[0:0] s577, in577_1, in577_2;
    wire c577;
    assign in577_1 = {pp46[73]};
    assign in577_2 = {pp47[72]};
    Full_Adder FA_577(s577, c577, in577_1, in577_2, pp45[74]);
    wire[0:0] s578, in578_1, in578_2;
    wire c578;
    assign in578_1 = {pp49[70]};
    assign in578_2 = {pp50[69]};
    Full_Adder FA_578(s578, c578, in578_1, in578_2, pp48[71]);
    wire[0:0] s579, in579_1, in579_2;
    wire c579;
    assign in579_1 = {pp52[67]};
    assign in579_2 = {pp53[66]};
    Full_Adder FA_579(s579, c579, in579_1, in579_2, pp51[68]);
    wire[0:0] s580, in580_1, in580_2;
    wire c580;
    assign in580_1 = {pp55[64]};
    assign in580_2 = {pp56[63]};
    Full_Adder FA_580(s580, c580, in580_1, in580_2, pp54[65]);
    wire[0:0] s581, in581_1, in581_2;
    wire c581;
    assign in581_1 = {pp58[61]};
    assign in581_2 = {pp59[60]};
    Full_Adder FA_581(s581, c581, in581_1, in581_2, pp57[62]);
    wire[0:0] s582, in582_1, in582_2;
    wire c582;
    assign in582_1 = {pp61[58]};
    assign in582_2 = {pp62[57]};
    Full_Adder FA_582(s582, c582, in582_1, in582_2, pp60[59]);
    wire[0:0] s583, in583_1, in583_2;
    wire c583;
    assign in583_1 = {pp64[55]};
    assign in583_2 = {pp65[54]};
    Full_Adder FA_583(s583, c583, in583_1, in583_2, pp63[56]);
    wire[0:0] s584, in584_1, in584_2;
    wire c584;
    assign in584_1 = {pp67[52]};
    assign in584_2 = {pp68[51]};
    Full_Adder FA_584(s584, c584, in584_1, in584_2, pp66[53]);
    wire[0:0] s585, in585_1, in585_2;
    wire c585;
    assign in585_1 = {pp70[49]};
    assign in585_2 = {pp71[48]};
    Full_Adder FA_585(s585, c585, in585_1, in585_2, pp69[50]);
    wire[0:0] s586, in586_1, in586_2;
    wire c586;
    assign in586_1 = {pp73[46]};
    assign in586_2 = {pp74[45]};
    Full_Adder FA_586(s586, c586, in586_1, in586_2, pp72[47]);
    wire[0:0] s587, in587_1, in587_2;
    wire c587;
    assign in587_1 = {pp76[43]};
    assign in587_2 = {pp77[42]};
    Full_Adder FA_587(s587, c587, in587_1, in587_2, pp75[44]);
    wire[0:0] s588, in588_1, in588_2;
    wire c588;
    assign in588_1 = {pp79[40]};
    assign in588_2 = {pp80[39]};
    Full_Adder FA_588(s588, c588, in588_1, in588_2, pp78[41]);
    wire[0:0] s589, in589_1, in589_2;
    wire c589;
    assign in589_1 = {pp82[37]};
    assign in589_2 = {pp83[36]};
    Full_Adder FA_589(s589, c589, in589_1, in589_2, pp81[38]);
    wire[0:0] s590, in590_1, in590_2;
    wire c590;
    assign in590_1 = {pp85[34]};
    assign in590_2 = {pp86[33]};
    Full_Adder FA_590(s590, c590, in590_1, in590_2, pp84[35]);
    wire[0:0] s591, in591_1, in591_2;
    wire c591;
    assign in591_1 = {pp88[31]};
    assign in591_2 = {pp89[30]};
    Full_Adder FA_591(s591, c591, in591_1, in591_2, pp87[32]);
    wire[0:0] s592, in592_1, in592_2;
    wire c592;
    assign in592_1 = {pp91[28]};
    assign in592_2 = {pp92[27]};
    Full_Adder FA_592(s592, c592, in592_1, in592_2, pp90[29]);
    wire[0:0] s593, in593_1, in593_2;
    wire c593;
    assign in593_1 = {pp94[25]};
    assign in593_2 = {pp95[24]};
    Full_Adder FA_593(s593, c593, in593_1, in593_2, pp93[26]);
    wire[0:0] s594, in594_1, in594_2;
    wire c594;
    assign in594_1 = {pp97[22]};
    assign in594_2 = {pp98[21]};
    Full_Adder FA_594(s594, c594, in594_1, in594_2, pp96[23]);
    wire[0:0] s595, in595_1, in595_2;
    wire c595;
    assign in595_1 = {pp99[20]};
    assign in595_2 = {pp100[19]};
    Half_Adder HA_595(s595, c595, in595_1, in595_2);
    wire[0:0] s596, in596_1, in596_2;
    wire c596;
    assign in596_1 = {pp1[119]};
    assign in596_2 = {pp2[118]};
    Full_Adder FA_596(s596, c596, in596_1, in596_2, pp0[120]);
    wire[0:0] s597, in597_1, in597_2;
    wire c597;
    assign in597_1 = {pp4[116]};
    assign in597_2 = {pp5[115]};
    Full_Adder FA_597(s597, c597, in597_1, in597_2, pp3[117]);
    wire[0:0] s598, in598_1, in598_2;
    wire c598;
    assign in598_1 = {pp7[113]};
    assign in598_2 = {pp8[112]};
    Full_Adder FA_598(s598, c598, in598_1, in598_2, pp6[114]);
    wire[0:0] s599, in599_1, in599_2;
    wire c599;
    assign in599_1 = {pp10[110]};
    assign in599_2 = {pp11[109]};
    Full_Adder FA_599(s599, c599, in599_1, in599_2, pp9[111]);
    wire[0:0] s600, in600_1, in600_2;
    wire c600;
    assign in600_1 = {pp13[107]};
    assign in600_2 = {pp14[106]};
    Full_Adder FA_600(s600, c600, in600_1, in600_2, pp12[108]);
    wire[0:0] s601, in601_1, in601_2;
    wire c601;
    assign in601_1 = {pp16[104]};
    assign in601_2 = {pp17[103]};
    Full_Adder FA_601(s601, c601, in601_1, in601_2, pp15[105]);
    wire[0:0] s602, in602_1, in602_2;
    wire c602;
    assign in602_1 = {pp19[101]};
    assign in602_2 = {pp20[100]};
    Full_Adder FA_602(s602, c602, in602_1, in602_2, pp18[102]);
    wire[0:0] s603, in603_1, in603_2;
    wire c603;
    assign in603_1 = {pp22[98]};
    assign in603_2 = {pp23[97]};
    Full_Adder FA_603(s603, c603, in603_1, in603_2, pp21[99]);
    wire[0:0] s604, in604_1, in604_2;
    wire c604;
    assign in604_1 = {pp25[95]};
    assign in604_2 = {pp26[94]};
    Full_Adder FA_604(s604, c604, in604_1, in604_2, pp24[96]);
    wire[0:0] s605, in605_1, in605_2;
    wire c605;
    assign in605_1 = {pp28[92]};
    assign in605_2 = {pp29[91]};
    Full_Adder FA_605(s605, c605, in605_1, in605_2, pp27[93]);
    wire[0:0] s606, in606_1, in606_2;
    wire c606;
    assign in606_1 = {pp31[89]};
    assign in606_2 = {pp32[88]};
    Full_Adder FA_606(s606, c606, in606_1, in606_2, pp30[90]);
    wire[0:0] s607, in607_1, in607_2;
    wire c607;
    assign in607_1 = {pp34[86]};
    assign in607_2 = {pp35[85]};
    Full_Adder FA_607(s607, c607, in607_1, in607_2, pp33[87]);
    wire[0:0] s608, in608_1, in608_2;
    wire c608;
    assign in608_1 = {pp37[83]};
    assign in608_2 = {pp38[82]};
    Full_Adder FA_608(s608, c608, in608_1, in608_2, pp36[84]);
    wire[0:0] s609, in609_1, in609_2;
    wire c609;
    assign in609_1 = {pp40[80]};
    assign in609_2 = {pp41[79]};
    Full_Adder FA_609(s609, c609, in609_1, in609_2, pp39[81]);
    wire[0:0] s610, in610_1, in610_2;
    wire c610;
    assign in610_1 = {pp43[77]};
    assign in610_2 = {pp44[76]};
    Full_Adder FA_610(s610, c610, in610_1, in610_2, pp42[78]);
    wire[0:0] s611, in611_1, in611_2;
    wire c611;
    assign in611_1 = {pp46[74]};
    assign in611_2 = {pp47[73]};
    Full_Adder FA_611(s611, c611, in611_1, in611_2, pp45[75]);
    wire[0:0] s612, in612_1, in612_2;
    wire c612;
    assign in612_1 = {pp49[71]};
    assign in612_2 = {pp50[70]};
    Full_Adder FA_612(s612, c612, in612_1, in612_2, pp48[72]);
    wire[0:0] s613, in613_1, in613_2;
    wire c613;
    assign in613_1 = {pp52[68]};
    assign in613_2 = {pp53[67]};
    Full_Adder FA_613(s613, c613, in613_1, in613_2, pp51[69]);
    wire[0:0] s614, in614_1, in614_2;
    wire c614;
    assign in614_1 = {pp55[65]};
    assign in614_2 = {pp56[64]};
    Full_Adder FA_614(s614, c614, in614_1, in614_2, pp54[66]);
    wire[0:0] s615, in615_1, in615_2;
    wire c615;
    assign in615_1 = {pp58[62]};
    assign in615_2 = {pp59[61]};
    Full_Adder FA_615(s615, c615, in615_1, in615_2, pp57[63]);
    wire[0:0] s616, in616_1, in616_2;
    wire c616;
    assign in616_1 = {pp61[59]};
    assign in616_2 = {pp62[58]};
    Full_Adder FA_616(s616, c616, in616_1, in616_2, pp60[60]);
    wire[0:0] s617, in617_1, in617_2;
    wire c617;
    assign in617_1 = {pp64[56]};
    assign in617_2 = {pp65[55]};
    Full_Adder FA_617(s617, c617, in617_1, in617_2, pp63[57]);
    wire[0:0] s618, in618_1, in618_2;
    wire c618;
    assign in618_1 = {pp67[53]};
    assign in618_2 = {pp68[52]};
    Full_Adder FA_618(s618, c618, in618_1, in618_2, pp66[54]);
    wire[0:0] s619, in619_1, in619_2;
    wire c619;
    assign in619_1 = {pp70[50]};
    assign in619_2 = {pp71[49]};
    Full_Adder FA_619(s619, c619, in619_1, in619_2, pp69[51]);
    wire[0:0] s620, in620_1, in620_2;
    wire c620;
    assign in620_1 = {pp73[47]};
    assign in620_2 = {pp74[46]};
    Full_Adder FA_620(s620, c620, in620_1, in620_2, pp72[48]);
    wire[0:0] s621, in621_1, in621_2;
    wire c621;
    assign in621_1 = {pp76[44]};
    assign in621_2 = {pp77[43]};
    Full_Adder FA_621(s621, c621, in621_1, in621_2, pp75[45]);
    wire[0:0] s622, in622_1, in622_2;
    wire c622;
    assign in622_1 = {pp79[41]};
    assign in622_2 = {pp80[40]};
    Full_Adder FA_622(s622, c622, in622_1, in622_2, pp78[42]);
    wire[0:0] s623, in623_1, in623_2;
    wire c623;
    assign in623_1 = {pp82[38]};
    assign in623_2 = {pp83[37]};
    Full_Adder FA_623(s623, c623, in623_1, in623_2, pp81[39]);
    wire[0:0] s624, in624_1, in624_2;
    wire c624;
    assign in624_1 = {pp85[35]};
    assign in624_2 = {pp86[34]};
    Full_Adder FA_624(s624, c624, in624_1, in624_2, pp84[36]);
    wire[0:0] s625, in625_1, in625_2;
    wire c625;
    assign in625_1 = {pp88[32]};
    assign in625_2 = {pp89[31]};
    Full_Adder FA_625(s625, c625, in625_1, in625_2, pp87[33]);
    wire[0:0] s626, in626_1, in626_2;
    wire c626;
    assign in626_1 = {pp91[29]};
    assign in626_2 = {pp92[28]};
    Full_Adder FA_626(s626, c626, in626_1, in626_2, pp90[30]);
    wire[0:0] s627, in627_1, in627_2;
    wire c627;
    assign in627_1 = {pp94[26]};
    assign in627_2 = {pp95[25]};
    Full_Adder FA_627(s627, c627, in627_1, in627_2, pp93[27]);
    wire[0:0] s628, in628_1, in628_2;
    wire c628;
    assign in628_1 = {pp97[23]};
    assign in628_2 = {pp98[22]};
    Full_Adder FA_628(s628, c628, in628_1, in628_2, pp96[24]);
    wire[0:0] s629, in629_1, in629_2;
    wire c629;
    assign in629_1 = {pp100[20]};
    assign in629_2 = {pp101[19]};
    Full_Adder FA_629(s629, c629, in629_1, in629_2, pp99[21]);
    wire[0:0] s630, in630_1, in630_2;
    wire c630;
    assign in630_1 = {pp102[18]};
    assign in630_2 = {pp103[17]};
    Half_Adder HA_630(s630, c630, in630_1, in630_2);
    wire[0:0] s631, in631_1, in631_2;
    wire c631;
    assign in631_1 = {pp1[120]};
    assign in631_2 = {pp2[119]};
    Full_Adder FA_631(s631, c631, in631_1, in631_2, pp0[121]);
    wire[0:0] s632, in632_1, in632_2;
    wire c632;
    assign in632_1 = {pp4[117]};
    assign in632_2 = {pp5[116]};
    Full_Adder FA_632(s632, c632, in632_1, in632_2, pp3[118]);
    wire[0:0] s633, in633_1, in633_2;
    wire c633;
    assign in633_1 = {pp7[114]};
    assign in633_2 = {pp8[113]};
    Full_Adder FA_633(s633, c633, in633_1, in633_2, pp6[115]);
    wire[0:0] s634, in634_1, in634_2;
    wire c634;
    assign in634_1 = {pp10[111]};
    assign in634_2 = {pp11[110]};
    Full_Adder FA_634(s634, c634, in634_1, in634_2, pp9[112]);
    wire[0:0] s635, in635_1, in635_2;
    wire c635;
    assign in635_1 = {pp13[108]};
    assign in635_2 = {pp14[107]};
    Full_Adder FA_635(s635, c635, in635_1, in635_2, pp12[109]);
    wire[0:0] s636, in636_1, in636_2;
    wire c636;
    assign in636_1 = {pp16[105]};
    assign in636_2 = {pp17[104]};
    Full_Adder FA_636(s636, c636, in636_1, in636_2, pp15[106]);
    wire[0:0] s637, in637_1, in637_2;
    wire c637;
    assign in637_1 = {pp19[102]};
    assign in637_2 = {pp20[101]};
    Full_Adder FA_637(s637, c637, in637_1, in637_2, pp18[103]);
    wire[0:0] s638, in638_1, in638_2;
    wire c638;
    assign in638_1 = {pp22[99]};
    assign in638_2 = {pp23[98]};
    Full_Adder FA_638(s638, c638, in638_1, in638_2, pp21[100]);
    wire[0:0] s639, in639_1, in639_2;
    wire c639;
    assign in639_1 = {pp25[96]};
    assign in639_2 = {pp26[95]};
    Full_Adder FA_639(s639, c639, in639_1, in639_2, pp24[97]);
    wire[0:0] s640, in640_1, in640_2;
    wire c640;
    assign in640_1 = {pp28[93]};
    assign in640_2 = {pp29[92]};
    Full_Adder FA_640(s640, c640, in640_1, in640_2, pp27[94]);
    wire[0:0] s641, in641_1, in641_2;
    wire c641;
    assign in641_1 = {pp31[90]};
    assign in641_2 = {pp32[89]};
    Full_Adder FA_641(s641, c641, in641_1, in641_2, pp30[91]);
    wire[0:0] s642, in642_1, in642_2;
    wire c642;
    assign in642_1 = {pp34[87]};
    assign in642_2 = {pp35[86]};
    Full_Adder FA_642(s642, c642, in642_1, in642_2, pp33[88]);
    wire[0:0] s643, in643_1, in643_2;
    wire c643;
    assign in643_1 = {pp37[84]};
    assign in643_2 = {pp38[83]};
    Full_Adder FA_643(s643, c643, in643_1, in643_2, pp36[85]);
    wire[0:0] s644, in644_1, in644_2;
    wire c644;
    assign in644_1 = {pp40[81]};
    assign in644_2 = {pp41[80]};
    Full_Adder FA_644(s644, c644, in644_1, in644_2, pp39[82]);
    wire[0:0] s645, in645_1, in645_2;
    wire c645;
    assign in645_1 = {pp43[78]};
    assign in645_2 = {pp44[77]};
    Full_Adder FA_645(s645, c645, in645_1, in645_2, pp42[79]);
    wire[0:0] s646, in646_1, in646_2;
    wire c646;
    assign in646_1 = {pp46[75]};
    assign in646_2 = {pp47[74]};
    Full_Adder FA_646(s646, c646, in646_1, in646_2, pp45[76]);
    wire[0:0] s647, in647_1, in647_2;
    wire c647;
    assign in647_1 = {pp49[72]};
    assign in647_2 = {pp50[71]};
    Full_Adder FA_647(s647, c647, in647_1, in647_2, pp48[73]);
    wire[0:0] s648, in648_1, in648_2;
    wire c648;
    assign in648_1 = {pp52[69]};
    assign in648_2 = {pp53[68]};
    Full_Adder FA_648(s648, c648, in648_1, in648_2, pp51[70]);
    wire[0:0] s649, in649_1, in649_2;
    wire c649;
    assign in649_1 = {pp55[66]};
    assign in649_2 = {pp56[65]};
    Full_Adder FA_649(s649, c649, in649_1, in649_2, pp54[67]);
    wire[0:0] s650, in650_1, in650_2;
    wire c650;
    assign in650_1 = {pp58[63]};
    assign in650_2 = {pp59[62]};
    Full_Adder FA_650(s650, c650, in650_1, in650_2, pp57[64]);
    wire[0:0] s651, in651_1, in651_2;
    wire c651;
    assign in651_1 = {pp61[60]};
    assign in651_2 = {pp62[59]};
    Full_Adder FA_651(s651, c651, in651_1, in651_2, pp60[61]);
    wire[0:0] s652, in652_1, in652_2;
    wire c652;
    assign in652_1 = {pp64[57]};
    assign in652_2 = {pp65[56]};
    Full_Adder FA_652(s652, c652, in652_1, in652_2, pp63[58]);
    wire[0:0] s653, in653_1, in653_2;
    wire c653;
    assign in653_1 = {pp67[54]};
    assign in653_2 = {pp68[53]};
    Full_Adder FA_653(s653, c653, in653_1, in653_2, pp66[55]);
    wire[0:0] s654, in654_1, in654_2;
    wire c654;
    assign in654_1 = {pp70[51]};
    assign in654_2 = {pp71[50]};
    Full_Adder FA_654(s654, c654, in654_1, in654_2, pp69[52]);
    wire[0:0] s655, in655_1, in655_2;
    wire c655;
    assign in655_1 = {pp73[48]};
    assign in655_2 = {pp74[47]};
    Full_Adder FA_655(s655, c655, in655_1, in655_2, pp72[49]);
    wire[0:0] s656, in656_1, in656_2;
    wire c656;
    assign in656_1 = {pp76[45]};
    assign in656_2 = {pp77[44]};
    Full_Adder FA_656(s656, c656, in656_1, in656_2, pp75[46]);
    wire[0:0] s657, in657_1, in657_2;
    wire c657;
    assign in657_1 = {pp79[42]};
    assign in657_2 = {pp80[41]};
    Full_Adder FA_657(s657, c657, in657_1, in657_2, pp78[43]);
    wire[0:0] s658, in658_1, in658_2;
    wire c658;
    assign in658_1 = {pp82[39]};
    assign in658_2 = {pp83[38]};
    Full_Adder FA_658(s658, c658, in658_1, in658_2, pp81[40]);
    wire[0:0] s659, in659_1, in659_2;
    wire c659;
    assign in659_1 = {pp85[36]};
    assign in659_2 = {pp86[35]};
    Full_Adder FA_659(s659, c659, in659_1, in659_2, pp84[37]);
    wire[0:0] s660, in660_1, in660_2;
    wire c660;
    assign in660_1 = {pp88[33]};
    assign in660_2 = {pp89[32]};
    Full_Adder FA_660(s660, c660, in660_1, in660_2, pp87[34]);
    wire[0:0] s661, in661_1, in661_2;
    wire c661;
    assign in661_1 = {pp91[30]};
    assign in661_2 = {pp92[29]};
    Full_Adder FA_661(s661, c661, in661_1, in661_2, pp90[31]);
    wire[0:0] s662, in662_1, in662_2;
    wire c662;
    assign in662_1 = {pp94[27]};
    assign in662_2 = {pp95[26]};
    Full_Adder FA_662(s662, c662, in662_1, in662_2, pp93[28]);
    wire[0:0] s663, in663_1, in663_2;
    wire c663;
    assign in663_1 = {pp97[24]};
    assign in663_2 = {pp98[23]};
    Full_Adder FA_663(s663, c663, in663_1, in663_2, pp96[25]);
    wire[0:0] s664, in664_1, in664_2;
    wire c664;
    assign in664_1 = {pp100[21]};
    assign in664_2 = {pp101[20]};
    Full_Adder FA_664(s664, c664, in664_1, in664_2, pp99[22]);
    wire[0:0] s665, in665_1, in665_2;
    wire c665;
    assign in665_1 = {pp103[18]};
    assign in665_2 = {pp104[17]};
    Full_Adder FA_665(s665, c665, in665_1, in665_2, pp102[19]);
    wire[0:0] s666, in666_1, in666_2;
    wire c666;
    assign in666_1 = {pp105[16]};
    assign in666_2 = {pp106[15]};
    Half_Adder HA_666(s666, c666, in666_1, in666_2);
    wire[0:0] s667, in667_1, in667_2;
    wire c667;
    assign in667_1 = {pp1[121]};
    assign in667_2 = {pp2[120]};
    Full_Adder FA_667(s667, c667, in667_1, in667_2, pp0[122]);
    wire[0:0] s668, in668_1, in668_2;
    wire c668;
    assign in668_1 = {pp4[118]};
    assign in668_2 = {pp5[117]};
    Full_Adder FA_668(s668, c668, in668_1, in668_2, pp3[119]);
    wire[0:0] s669, in669_1, in669_2;
    wire c669;
    assign in669_1 = {pp7[115]};
    assign in669_2 = {pp8[114]};
    Full_Adder FA_669(s669, c669, in669_1, in669_2, pp6[116]);
    wire[0:0] s670, in670_1, in670_2;
    wire c670;
    assign in670_1 = {pp10[112]};
    assign in670_2 = {pp11[111]};
    Full_Adder FA_670(s670, c670, in670_1, in670_2, pp9[113]);
    wire[0:0] s671, in671_1, in671_2;
    wire c671;
    assign in671_1 = {pp13[109]};
    assign in671_2 = {pp14[108]};
    Full_Adder FA_671(s671, c671, in671_1, in671_2, pp12[110]);
    wire[0:0] s672, in672_1, in672_2;
    wire c672;
    assign in672_1 = {pp16[106]};
    assign in672_2 = {pp17[105]};
    Full_Adder FA_672(s672, c672, in672_1, in672_2, pp15[107]);
    wire[0:0] s673, in673_1, in673_2;
    wire c673;
    assign in673_1 = {pp19[103]};
    assign in673_2 = {pp20[102]};
    Full_Adder FA_673(s673, c673, in673_1, in673_2, pp18[104]);
    wire[0:0] s674, in674_1, in674_2;
    wire c674;
    assign in674_1 = {pp22[100]};
    assign in674_2 = {pp23[99]};
    Full_Adder FA_674(s674, c674, in674_1, in674_2, pp21[101]);
    wire[0:0] s675, in675_1, in675_2;
    wire c675;
    assign in675_1 = {pp25[97]};
    assign in675_2 = {pp26[96]};
    Full_Adder FA_675(s675, c675, in675_1, in675_2, pp24[98]);
    wire[0:0] s676, in676_1, in676_2;
    wire c676;
    assign in676_1 = {pp28[94]};
    assign in676_2 = {pp29[93]};
    Full_Adder FA_676(s676, c676, in676_1, in676_2, pp27[95]);
    wire[0:0] s677, in677_1, in677_2;
    wire c677;
    assign in677_1 = {pp31[91]};
    assign in677_2 = {pp32[90]};
    Full_Adder FA_677(s677, c677, in677_1, in677_2, pp30[92]);
    wire[0:0] s678, in678_1, in678_2;
    wire c678;
    assign in678_1 = {pp34[88]};
    assign in678_2 = {pp35[87]};
    Full_Adder FA_678(s678, c678, in678_1, in678_2, pp33[89]);
    wire[0:0] s679, in679_1, in679_2;
    wire c679;
    assign in679_1 = {pp37[85]};
    assign in679_2 = {pp38[84]};
    Full_Adder FA_679(s679, c679, in679_1, in679_2, pp36[86]);
    wire[0:0] s680, in680_1, in680_2;
    wire c680;
    assign in680_1 = {pp40[82]};
    assign in680_2 = {pp41[81]};
    Full_Adder FA_680(s680, c680, in680_1, in680_2, pp39[83]);
    wire[0:0] s681, in681_1, in681_2;
    wire c681;
    assign in681_1 = {pp43[79]};
    assign in681_2 = {pp44[78]};
    Full_Adder FA_681(s681, c681, in681_1, in681_2, pp42[80]);
    wire[0:0] s682, in682_1, in682_2;
    wire c682;
    assign in682_1 = {pp46[76]};
    assign in682_2 = {pp47[75]};
    Full_Adder FA_682(s682, c682, in682_1, in682_2, pp45[77]);
    wire[0:0] s683, in683_1, in683_2;
    wire c683;
    assign in683_1 = {pp49[73]};
    assign in683_2 = {pp50[72]};
    Full_Adder FA_683(s683, c683, in683_1, in683_2, pp48[74]);
    wire[0:0] s684, in684_1, in684_2;
    wire c684;
    assign in684_1 = {pp52[70]};
    assign in684_2 = {pp53[69]};
    Full_Adder FA_684(s684, c684, in684_1, in684_2, pp51[71]);
    wire[0:0] s685, in685_1, in685_2;
    wire c685;
    assign in685_1 = {pp55[67]};
    assign in685_2 = {pp56[66]};
    Full_Adder FA_685(s685, c685, in685_1, in685_2, pp54[68]);
    wire[0:0] s686, in686_1, in686_2;
    wire c686;
    assign in686_1 = {pp58[64]};
    assign in686_2 = {pp59[63]};
    Full_Adder FA_686(s686, c686, in686_1, in686_2, pp57[65]);
    wire[0:0] s687, in687_1, in687_2;
    wire c687;
    assign in687_1 = {pp61[61]};
    assign in687_2 = {pp62[60]};
    Full_Adder FA_687(s687, c687, in687_1, in687_2, pp60[62]);
    wire[0:0] s688, in688_1, in688_2;
    wire c688;
    assign in688_1 = {pp64[58]};
    assign in688_2 = {pp65[57]};
    Full_Adder FA_688(s688, c688, in688_1, in688_2, pp63[59]);
    wire[0:0] s689, in689_1, in689_2;
    wire c689;
    assign in689_1 = {pp67[55]};
    assign in689_2 = {pp68[54]};
    Full_Adder FA_689(s689, c689, in689_1, in689_2, pp66[56]);
    wire[0:0] s690, in690_1, in690_2;
    wire c690;
    assign in690_1 = {pp70[52]};
    assign in690_2 = {pp71[51]};
    Full_Adder FA_690(s690, c690, in690_1, in690_2, pp69[53]);
    wire[0:0] s691, in691_1, in691_2;
    wire c691;
    assign in691_1 = {pp73[49]};
    assign in691_2 = {pp74[48]};
    Full_Adder FA_691(s691, c691, in691_1, in691_2, pp72[50]);
    wire[0:0] s692, in692_1, in692_2;
    wire c692;
    assign in692_1 = {pp76[46]};
    assign in692_2 = {pp77[45]};
    Full_Adder FA_692(s692, c692, in692_1, in692_2, pp75[47]);
    wire[0:0] s693, in693_1, in693_2;
    wire c693;
    assign in693_1 = {pp79[43]};
    assign in693_2 = {pp80[42]};
    Full_Adder FA_693(s693, c693, in693_1, in693_2, pp78[44]);
    wire[0:0] s694, in694_1, in694_2;
    wire c694;
    assign in694_1 = {pp82[40]};
    assign in694_2 = {pp83[39]};
    Full_Adder FA_694(s694, c694, in694_1, in694_2, pp81[41]);
    wire[0:0] s695, in695_1, in695_2;
    wire c695;
    assign in695_1 = {pp85[37]};
    assign in695_2 = {pp86[36]};
    Full_Adder FA_695(s695, c695, in695_1, in695_2, pp84[38]);
    wire[0:0] s696, in696_1, in696_2;
    wire c696;
    assign in696_1 = {pp88[34]};
    assign in696_2 = {pp89[33]};
    Full_Adder FA_696(s696, c696, in696_1, in696_2, pp87[35]);
    wire[0:0] s697, in697_1, in697_2;
    wire c697;
    assign in697_1 = {pp91[31]};
    assign in697_2 = {pp92[30]};
    Full_Adder FA_697(s697, c697, in697_1, in697_2, pp90[32]);
    wire[0:0] s698, in698_1, in698_2;
    wire c698;
    assign in698_1 = {pp94[28]};
    assign in698_2 = {pp95[27]};
    Full_Adder FA_698(s698, c698, in698_1, in698_2, pp93[29]);
    wire[0:0] s699, in699_1, in699_2;
    wire c699;
    assign in699_1 = {pp97[25]};
    assign in699_2 = {pp98[24]};
    Full_Adder FA_699(s699, c699, in699_1, in699_2, pp96[26]);
    wire[0:0] s700, in700_1, in700_2;
    wire c700;
    assign in700_1 = {pp100[22]};
    assign in700_2 = {pp101[21]};
    Full_Adder FA_700(s700, c700, in700_1, in700_2, pp99[23]);
    wire[0:0] s701, in701_1, in701_2;
    wire c701;
    assign in701_1 = {pp103[19]};
    assign in701_2 = {pp104[18]};
    Full_Adder FA_701(s701, c701, in701_1, in701_2, pp102[20]);
    wire[0:0] s702, in702_1, in702_2;
    wire c702;
    assign in702_1 = {pp106[16]};
    assign in702_2 = {pp107[15]};
    Full_Adder FA_702(s702, c702, in702_1, in702_2, pp105[17]);
    wire[0:0] s703, in703_1, in703_2;
    wire c703;
    assign in703_1 = {pp108[14]};
    assign in703_2 = {pp109[13]};
    Half_Adder HA_703(s703, c703, in703_1, in703_2);
    wire[0:0] s704, in704_1, in704_2;
    wire c704;
    assign in704_1 = {pp1[122]};
    assign in704_2 = {pp2[121]};
    Full_Adder FA_704(s704, c704, in704_1, in704_2, pp0[123]);
    wire[0:0] s705, in705_1, in705_2;
    wire c705;
    assign in705_1 = {pp4[119]};
    assign in705_2 = {pp5[118]};
    Full_Adder FA_705(s705, c705, in705_1, in705_2, pp3[120]);
    wire[0:0] s706, in706_1, in706_2;
    wire c706;
    assign in706_1 = {pp7[116]};
    assign in706_2 = {pp8[115]};
    Full_Adder FA_706(s706, c706, in706_1, in706_2, pp6[117]);
    wire[0:0] s707, in707_1, in707_2;
    wire c707;
    assign in707_1 = {pp10[113]};
    assign in707_2 = {pp11[112]};
    Full_Adder FA_707(s707, c707, in707_1, in707_2, pp9[114]);
    wire[0:0] s708, in708_1, in708_2;
    wire c708;
    assign in708_1 = {pp13[110]};
    assign in708_2 = {pp14[109]};
    Full_Adder FA_708(s708, c708, in708_1, in708_2, pp12[111]);
    wire[0:0] s709, in709_1, in709_2;
    wire c709;
    assign in709_1 = {pp16[107]};
    assign in709_2 = {pp17[106]};
    Full_Adder FA_709(s709, c709, in709_1, in709_2, pp15[108]);
    wire[0:0] s710, in710_1, in710_2;
    wire c710;
    assign in710_1 = {pp19[104]};
    assign in710_2 = {pp20[103]};
    Full_Adder FA_710(s710, c710, in710_1, in710_2, pp18[105]);
    wire[0:0] s711, in711_1, in711_2;
    wire c711;
    assign in711_1 = {pp22[101]};
    assign in711_2 = {pp23[100]};
    Full_Adder FA_711(s711, c711, in711_1, in711_2, pp21[102]);
    wire[0:0] s712, in712_1, in712_2;
    wire c712;
    assign in712_1 = {pp25[98]};
    assign in712_2 = {pp26[97]};
    Full_Adder FA_712(s712, c712, in712_1, in712_2, pp24[99]);
    wire[0:0] s713, in713_1, in713_2;
    wire c713;
    assign in713_1 = {pp28[95]};
    assign in713_2 = {pp29[94]};
    Full_Adder FA_713(s713, c713, in713_1, in713_2, pp27[96]);
    wire[0:0] s714, in714_1, in714_2;
    wire c714;
    assign in714_1 = {pp31[92]};
    assign in714_2 = {pp32[91]};
    Full_Adder FA_714(s714, c714, in714_1, in714_2, pp30[93]);
    wire[0:0] s715, in715_1, in715_2;
    wire c715;
    assign in715_1 = {pp34[89]};
    assign in715_2 = {pp35[88]};
    Full_Adder FA_715(s715, c715, in715_1, in715_2, pp33[90]);
    wire[0:0] s716, in716_1, in716_2;
    wire c716;
    assign in716_1 = {pp37[86]};
    assign in716_2 = {pp38[85]};
    Full_Adder FA_716(s716, c716, in716_1, in716_2, pp36[87]);
    wire[0:0] s717, in717_1, in717_2;
    wire c717;
    assign in717_1 = {pp40[83]};
    assign in717_2 = {pp41[82]};
    Full_Adder FA_717(s717, c717, in717_1, in717_2, pp39[84]);
    wire[0:0] s718, in718_1, in718_2;
    wire c718;
    assign in718_1 = {pp43[80]};
    assign in718_2 = {pp44[79]};
    Full_Adder FA_718(s718, c718, in718_1, in718_2, pp42[81]);
    wire[0:0] s719, in719_1, in719_2;
    wire c719;
    assign in719_1 = {pp46[77]};
    assign in719_2 = {pp47[76]};
    Full_Adder FA_719(s719, c719, in719_1, in719_2, pp45[78]);
    wire[0:0] s720, in720_1, in720_2;
    wire c720;
    assign in720_1 = {pp49[74]};
    assign in720_2 = {pp50[73]};
    Full_Adder FA_720(s720, c720, in720_1, in720_2, pp48[75]);
    wire[0:0] s721, in721_1, in721_2;
    wire c721;
    assign in721_1 = {pp52[71]};
    assign in721_2 = {pp53[70]};
    Full_Adder FA_721(s721, c721, in721_1, in721_2, pp51[72]);
    wire[0:0] s722, in722_1, in722_2;
    wire c722;
    assign in722_1 = {pp55[68]};
    assign in722_2 = {pp56[67]};
    Full_Adder FA_722(s722, c722, in722_1, in722_2, pp54[69]);
    wire[0:0] s723, in723_1, in723_2;
    wire c723;
    assign in723_1 = {pp58[65]};
    assign in723_2 = {pp59[64]};
    Full_Adder FA_723(s723, c723, in723_1, in723_2, pp57[66]);
    wire[0:0] s724, in724_1, in724_2;
    wire c724;
    assign in724_1 = {pp61[62]};
    assign in724_2 = {pp62[61]};
    Full_Adder FA_724(s724, c724, in724_1, in724_2, pp60[63]);
    wire[0:0] s725, in725_1, in725_2;
    wire c725;
    assign in725_1 = {pp64[59]};
    assign in725_2 = {pp65[58]};
    Full_Adder FA_725(s725, c725, in725_1, in725_2, pp63[60]);
    wire[0:0] s726, in726_1, in726_2;
    wire c726;
    assign in726_1 = {pp67[56]};
    assign in726_2 = {pp68[55]};
    Full_Adder FA_726(s726, c726, in726_1, in726_2, pp66[57]);
    wire[0:0] s727, in727_1, in727_2;
    wire c727;
    assign in727_1 = {pp70[53]};
    assign in727_2 = {pp71[52]};
    Full_Adder FA_727(s727, c727, in727_1, in727_2, pp69[54]);
    wire[0:0] s728, in728_1, in728_2;
    wire c728;
    assign in728_1 = {pp73[50]};
    assign in728_2 = {pp74[49]};
    Full_Adder FA_728(s728, c728, in728_1, in728_2, pp72[51]);
    wire[0:0] s729, in729_1, in729_2;
    wire c729;
    assign in729_1 = {pp76[47]};
    assign in729_2 = {pp77[46]};
    Full_Adder FA_729(s729, c729, in729_1, in729_2, pp75[48]);
    wire[0:0] s730, in730_1, in730_2;
    wire c730;
    assign in730_1 = {pp79[44]};
    assign in730_2 = {pp80[43]};
    Full_Adder FA_730(s730, c730, in730_1, in730_2, pp78[45]);
    wire[0:0] s731, in731_1, in731_2;
    wire c731;
    assign in731_1 = {pp82[41]};
    assign in731_2 = {pp83[40]};
    Full_Adder FA_731(s731, c731, in731_1, in731_2, pp81[42]);
    wire[0:0] s732, in732_1, in732_2;
    wire c732;
    assign in732_1 = {pp85[38]};
    assign in732_2 = {pp86[37]};
    Full_Adder FA_732(s732, c732, in732_1, in732_2, pp84[39]);
    wire[0:0] s733, in733_1, in733_2;
    wire c733;
    assign in733_1 = {pp88[35]};
    assign in733_2 = {pp89[34]};
    Full_Adder FA_733(s733, c733, in733_1, in733_2, pp87[36]);
    wire[0:0] s734, in734_1, in734_2;
    wire c734;
    assign in734_1 = {pp91[32]};
    assign in734_2 = {pp92[31]};
    Full_Adder FA_734(s734, c734, in734_1, in734_2, pp90[33]);
    wire[0:0] s735, in735_1, in735_2;
    wire c735;
    assign in735_1 = {pp94[29]};
    assign in735_2 = {pp95[28]};
    Full_Adder FA_735(s735, c735, in735_1, in735_2, pp93[30]);
    wire[0:0] s736, in736_1, in736_2;
    wire c736;
    assign in736_1 = {pp97[26]};
    assign in736_2 = {pp98[25]};
    Full_Adder FA_736(s736, c736, in736_1, in736_2, pp96[27]);
    wire[0:0] s737, in737_1, in737_2;
    wire c737;
    assign in737_1 = {pp100[23]};
    assign in737_2 = {pp101[22]};
    Full_Adder FA_737(s737, c737, in737_1, in737_2, pp99[24]);
    wire[0:0] s738, in738_1, in738_2;
    wire c738;
    assign in738_1 = {pp103[20]};
    assign in738_2 = {pp104[19]};
    Full_Adder FA_738(s738, c738, in738_1, in738_2, pp102[21]);
    wire[0:0] s739, in739_1, in739_2;
    wire c739;
    assign in739_1 = {pp106[17]};
    assign in739_2 = {pp107[16]};
    Full_Adder FA_739(s739, c739, in739_1, in739_2, pp105[18]);
    wire[0:0] s740, in740_1, in740_2;
    wire c740;
    assign in740_1 = {pp109[14]};
    assign in740_2 = {pp110[13]};
    Full_Adder FA_740(s740, c740, in740_1, in740_2, pp108[15]);
    wire[0:0] s741, in741_1, in741_2;
    wire c741;
    assign in741_1 = {pp111[12]};
    assign in741_2 = {pp112[11]};
    Half_Adder HA_741(s741, c741, in741_1, in741_2);
    wire[0:0] s742, in742_1, in742_2;
    wire c742;
    assign in742_1 = {pp1[123]};
    assign in742_2 = {pp2[122]};
    Full_Adder FA_742(s742, c742, in742_1, in742_2, pp0[124]);
    wire[0:0] s743, in743_1, in743_2;
    wire c743;
    assign in743_1 = {pp4[120]};
    assign in743_2 = {pp5[119]};
    Full_Adder FA_743(s743, c743, in743_1, in743_2, pp3[121]);
    wire[0:0] s744, in744_1, in744_2;
    wire c744;
    assign in744_1 = {pp7[117]};
    assign in744_2 = {pp8[116]};
    Full_Adder FA_744(s744, c744, in744_1, in744_2, pp6[118]);
    wire[0:0] s745, in745_1, in745_2;
    wire c745;
    assign in745_1 = {pp10[114]};
    assign in745_2 = {pp11[113]};
    Full_Adder FA_745(s745, c745, in745_1, in745_2, pp9[115]);
    wire[0:0] s746, in746_1, in746_2;
    wire c746;
    assign in746_1 = {pp13[111]};
    assign in746_2 = {pp14[110]};
    Full_Adder FA_746(s746, c746, in746_1, in746_2, pp12[112]);
    wire[0:0] s747, in747_1, in747_2;
    wire c747;
    assign in747_1 = {pp16[108]};
    assign in747_2 = {pp17[107]};
    Full_Adder FA_747(s747, c747, in747_1, in747_2, pp15[109]);
    wire[0:0] s748, in748_1, in748_2;
    wire c748;
    assign in748_1 = {pp19[105]};
    assign in748_2 = {pp20[104]};
    Full_Adder FA_748(s748, c748, in748_1, in748_2, pp18[106]);
    wire[0:0] s749, in749_1, in749_2;
    wire c749;
    assign in749_1 = {pp22[102]};
    assign in749_2 = {pp23[101]};
    Full_Adder FA_749(s749, c749, in749_1, in749_2, pp21[103]);
    wire[0:0] s750, in750_1, in750_2;
    wire c750;
    assign in750_1 = {pp25[99]};
    assign in750_2 = {pp26[98]};
    Full_Adder FA_750(s750, c750, in750_1, in750_2, pp24[100]);
    wire[0:0] s751, in751_1, in751_2;
    wire c751;
    assign in751_1 = {pp28[96]};
    assign in751_2 = {pp29[95]};
    Full_Adder FA_751(s751, c751, in751_1, in751_2, pp27[97]);
    wire[0:0] s752, in752_1, in752_2;
    wire c752;
    assign in752_1 = {pp31[93]};
    assign in752_2 = {pp32[92]};
    Full_Adder FA_752(s752, c752, in752_1, in752_2, pp30[94]);
    wire[0:0] s753, in753_1, in753_2;
    wire c753;
    assign in753_1 = {pp34[90]};
    assign in753_2 = {pp35[89]};
    Full_Adder FA_753(s753, c753, in753_1, in753_2, pp33[91]);
    wire[0:0] s754, in754_1, in754_2;
    wire c754;
    assign in754_1 = {pp37[87]};
    assign in754_2 = {pp38[86]};
    Full_Adder FA_754(s754, c754, in754_1, in754_2, pp36[88]);
    wire[0:0] s755, in755_1, in755_2;
    wire c755;
    assign in755_1 = {pp40[84]};
    assign in755_2 = {pp41[83]};
    Full_Adder FA_755(s755, c755, in755_1, in755_2, pp39[85]);
    wire[0:0] s756, in756_1, in756_2;
    wire c756;
    assign in756_1 = {pp43[81]};
    assign in756_2 = {pp44[80]};
    Full_Adder FA_756(s756, c756, in756_1, in756_2, pp42[82]);
    wire[0:0] s757, in757_1, in757_2;
    wire c757;
    assign in757_1 = {pp46[78]};
    assign in757_2 = {pp47[77]};
    Full_Adder FA_757(s757, c757, in757_1, in757_2, pp45[79]);
    wire[0:0] s758, in758_1, in758_2;
    wire c758;
    assign in758_1 = {pp49[75]};
    assign in758_2 = {pp50[74]};
    Full_Adder FA_758(s758, c758, in758_1, in758_2, pp48[76]);
    wire[0:0] s759, in759_1, in759_2;
    wire c759;
    assign in759_1 = {pp52[72]};
    assign in759_2 = {pp53[71]};
    Full_Adder FA_759(s759, c759, in759_1, in759_2, pp51[73]);
    wire[0:0] s760, in760_1, in760_2;
    wire c760;
    assign in760_1 = {pp55[69]};
    assign in760_2 = {pp56[68]};
    Full_Adder FA_760(s760, c760, in760_1, in760_2, pp54[70]);
    wire[0:0] s761, in761_1, in761_2;
    wire c761;
    assign in761_1 = {pp58[66]};
    assign in761_2 = {pp59[65]};
    Full_Adder FA_761(s761, c761, in761_1, in761_2, pp57[67]);
    wire[0:0] s762, in762_1, in762_2;
    wire c762;
    assign in762_1 = {pp61[63]};
    assign in762_2 = {pp62[62]};
    Full_Adder FA_762(s762, c762, in762_1, in762_2, pp60[64]);
    wire[0:0] s763, in763_1, in763_2;
    wire c763;
    assign in763_1 = {pp64[60]};
    assign in763_2 = {pp65[59]};
    Full_Adder FA_763(s763, c763, in763_1, in763_2, pp63[61]);
    wire[0:0] s764, in764_1, in764_2;
    wire c764;
    assign in764_1 = {pp67[57]};
    assign in764_2 = {pp68[56]};
    Full_Adder FA_764(s764, c764, in764_1, in764_2, pp66[58]);
    wire[0:0] s765, in765_1, in765_2;
    wire c765;
    assign in765_1 = {pp70[54]};
    assign in765_2 = {pp71[53]};
    Full_Adder FA_765(s765, c765, in765_1, in765_2, pp69[55]);
    wire[0:0] s766, in766_1, in766_2;
    wire c766;
    assign in766_1 = {pp73[51]};
    assign in766_2 = {pp74[50]};
    Full_Adder FA_766(s766, c766, in766_1, in766_2, pp72[52]);
    wire[0:0] s767, in767_1, in767_2;
    wire c767;
    assign in767_1 = {pp76[48]};
    assign in767_2 = {pp77[47]};
    Full_Adder FA_767(s767, c767, in767_1, in767_2, pp75[49]);
    wire[0:0] s768, in768_1, in768_2;
    wire c768;
    assign in768_1 = {pp79[45]};
    assign in768_2 = {pp80[44]};
    Full_Adder FA_768(s768, c768, in768_1, in768_2, pp78[46]);
    wire[0:0] s769, in769_1, in769_2;
    wire c769;
    assign in769_1 = {pp82[42]};
    assign in769_2 = {pp83[41]};
    Full_Adder FA_769(s769, c769, in769_1, in769_2, pp81[43]);
    wire[0:0] s770, in770_1, in770_2;
    wire c770;
    assign in770_1 = {pp85[39]};
    assign in770_2 = {pp86[38]};
    Full_Adder FA_770(s770, c770, in770_1, in770_2, pp84[40]);
    wire[0:0] s771, in771_1, in771_2;
    wire c771;
    assign in771_1 = {pp88[36]};
    assign in771_2 = {pp89[35]};
    Full_Adder FA_771(s771, c771, in771_1, in771_2, pp87[37]);
    wire[0:0] s772, in772_1, in772_2;
    wire c772;
    assign in772_1 = {pp91[33]};
    assign in772_2 = {pp92[32]};
    Full_Adder FA_772(s772, c772, in772_1, in772_2, pp90[34]);
    wire[0:0] s773, in773_1, in773_2;
    wire c773;
    assign in773_1 = {pp94[30]};
    assign in773_2 = {pp95[29]};
    Full_Adder FA_773(s773, c773, in773_1, in773_2, pp93[31]);
    wire[0:0] s774, in774_1, in774_2;
    wire c774;
    assign in774_1 = {pp97[27]};
    assign in774_2 = {pp98[26]};
    Full_Adder FA_774(s774, c774, in774_1, in774_2, pp96[28]);
    wire[0:0] s775, in775_1, in775_2;
    wire c775;
    assign in775_1 = {pp100[24]};
    assign in775_2 = {pp101[23]};
    Full_Adder FA_775(s775, c775, in775_1, in775_2, pp99[25]);
    wire[0:0] s776, in776_1, in776_2;
    wire c776;
    assign in776_1 = {pp103[21]};
    assign in776_2 = {pp104[20]};
    Full_Adder FA_776(s776, c776, in776_1, in776_2, pp102[22]);
    wire[0:0] s777, in777_1, in777_2;
    wire c777;
    assign in777_1 = {pp106[18]};
    assign in777_2 = {pp107[17]};
    Full_Adder FA_777(s777, c777, in777_1, in777_2, pp105[19]);
    wire[0:0] s778, in778_1, in778_2;
    wire c778;
    assign in778_1 = {pp109[15]};
    assign in778_2 = {pp110[14]};
    Full_Adder FA_778(s778, c778, in778_1, in778_2, pp108[16]);
    wire[0:0] s779, in779_1, in779_2;
    wire c779;
    assign in779_1 = {pp112[12]};
    assign in779_2 = {pp113[11]};
    Full_Adder FA_779(s779, c779, in779_1, in779_2, pp111[13]);
    wire[0:0] s780, in780_1, in780_2;
    wire c780;
    assign in780_1 = {pp114[10]};
    assign in780_2 = {pp115[9]};
    Half_Adder HA_780(s780, c780, in780_1, in780_2);
    wire[0:0] s781, in781_1, in781_2;
    wire c781;
    assign in781_1 = {pp1[124]};
    assign in781_2 = {pp2[123]};
    Full_Adder FA_781(s781, c781, in781_1, in781_2, pp0[125]);
    wire[0:0] s782, in782_1, in782_2;
    wire c782;
    assign in782_1 = {pp4[121]};
    assign in782_2 = {pp5[120]};
    Full_Adder FA_782(s782, c782, in782_1, in782_2, pp3[122]);
    wire[0:0] s783, in783_1, in783_2;
    wire c783;
    assign in783_1 = {pp7[118]};
    assign in783_2 = {pp8[117]};
    Full_Adder FA_783(s783, c783, in783_1, in783_2, pp6[119]);
    wire[0:0] s784, in784_1, in784_2;
    wire c784;
    assign in784_1 = {pp10[115]};
    assign in784_2 = {pp11[114]};
    Full_Adder FA_784(s784, c784, in784_1, in784_2, pp9[116]);
    wire[0:0] s785, in785_1, in785_2;
    wire c785;
    assign in785_1 = {pp13[112]};
    assign in785_2 = {pp14[111]};
    Full_Adder FA_785(s785, c785, in785_1, in785_2, pp12[113]);
    wire[0:0] s786, in786_1, in786_2;
    wire c786;
    assign in786_1 = {pp16[109]};
    assign in786_2 = {pp17[108]};
    Full_Adder FA_786(s786, c786, in786_1, in786_2, pp15[110]);
    wire[0:0] s787, in787_1, in787_2;
    wire c787;
    assign in787_1 = {pp19[106]};
    assign in787_2 = {pp20[105]};
    Full_Adder FA_787(s787, c787, in787_1, in787_2, pp18[107]);
    wire[0:0] s788, in788_1, in788_2;
    wire c788;
    assign in788_1 = {pp22[103]};
    assign in788_2 = {pp23[102]};
    Full_Adder FA_788(s788, c788, in788_1, in788_2, pp21[104]);
    wire[0:0] s789, in789_1, in789_2;
    wire c789;
    assign in789_1 = {pp25[100]};
    assign in789_2 = {pp26[99]};
    Full_Adder FA_789(s789, c789, in789_1, in789_2, pp24[101]);
    wire[0:0] s790, in790_1, in790_2;
    wire c790;
    assign in790_1 = {pp28[97]};
    assign in790_2 = {pp29[96]};
    Full_Adder FA_790(s790, c790, in790_1, in790_2, pp27[98]);
    wire[0:0] s791, in791_1, in791_2;
    wire c791;
    assign in791_1 = {pp31[94]};
    assign in791_2 = {pp32[93]};
    Full_Adder FA_791(s791, c791, in791_1, in791_2, pp30[95]);
    wire[0:0] s792, in792_1, in792_2;
    wire c792;
    assign in792_1 = {pp34[91]};
    assign in792_2 = {pp35[90]};
    Full_Adder FA_792(s792, c792, in792_1, in792_2, pp33[92]);
    wire[0:0] s793, in793_1, in793_2;
    wire c793;
    assign in793_1 = {pp37[88]};
    assign in793_2 = {pp38[87]};
    Full_Adder FA_793(s793, c793, in793_1, in793_2, pp36[89]);
    wire[0:0] s794, in794_1, in794_2;
    wire c794;
    assign in794_1 = {pp40[85]};
    assign in794_2 = {pp41[84]};
    Full_Adder FA_794(s794, c794, in794_1, in794_2, pp39[86]);
    wire[0:0] s795, in795_1, in795_2;
    wire c795;
    assign in795_1 = {pp43[82]};
    assign in795_2 = {pp44[81]};
    Full_Adder FA_795(s795, c795, in795_1, in795_2, pp42[83]);
    wire[0:0] s796, in796_1, in796_2;
    wire c796;
    assign in796_1 = {pp46[79]};
    assign in796_2 = {pp47[78]};
    Full_Adder FA_796(s796, c796, in796_1, in796_2, pp45[80]);
    wire[0:0] s797, in797_1, in797_2;
    wire c797;
    assign in797_1 = {pp49[76]};
    assign in797_2 = {pp50[75]};
    Full_Adder FA_797(s797, c797, in797_1, in797_2, pp48[77]);
    wire[0:0] s798, in798_1, in798_2;
    wire c798;
    assign in798_1 = {pp52[73]};
    assign in798_2 = {pp53[72]};
    Full_Adder FA_798(s798, c798, in798_1, in798_2, pp51[74]);
    wire[0:0] s799, in799_1, in799_2;
    wire c799;
    assign in799_1 = {pp55[70]};
    assign in799_2 = {pp56[69]};
    Full_Adder FA_799(s799, c799, in799_1, in799_2, pp54[71]);
    wire[0:0] s800, in800_1, in800_2;
    wire c800;
    assign in800_1 = {pp58[67]};
    assign in800_2 = {pp59[66]};
    Full_Adder FA_800(s800, c800, in800_1, in800_2, pp57[68]);
    wire[0:0] s801, in801_1, in801_2;
    wire c801;
    assign in801_1 = {pp61[64]};
    assign in801_2 = {pp62[63]};
    Full_Adder FA_801(s801, c801, in801_1, in801_2, pp60[65]);
    wire[0:0] s802, in802_1, in802_2;
    wire c802;
    assign in802_1 = {pp64[61]};
    assign in802_2 = {pp65[60]};
    Full_Adder FA_802(s802, c802, in802_1, in802_2, pp63[62]);
    wire[0:0] s803, in803_1, in803_2;
    wire c803;
    assign in803_1 = {pp67[58]};
    assign in803_2 = {pp68[57]};
    Full_Adder FA_803(s803, c803, in803_1, in803_2, pp66[59]);
    wire[0:0] s804, in804_1, in804_2;
    wire c804;
    assign in804_1 = {pp70[55]};
    assign in804_2 = {pp71[54]};
    Full_Adder FA_804(s804, c804, in804_1, in804_2, pp69[56]);
    wire[0:0] s805, in805_1, in805_2;
    wire c805;
    assign in805_1 = {pp73[52]};
    assign in805_2 = {pp74[51]};
    Full_Adder FA_805(s805, c805, in805_1, in805_2, pp72[53]);
    wire[0:0] s806, in806_1, in806_2;
    wire c806;
    assign in806_1 = {pp76[49]};
    assign in806_2 = {pp77[48]};
    Full_Adder FA_806(s806, c806, in806_1, in806_2, pp75[50]);
    wire[0:0] s807, in807_1, in807_2;
    wire c807;
    assign in807_1 = {pp79[46]};
    assign in807_2 = {pp80[45]};
    Full_Adder FA_807(s807, c807, in807_1, in807_2, pp78[47]);
    wire[0:0] s808, in808_1, in808_2;
    wire c808;
    assign in808_1 = {pp82[43]};
    assign in808_2 = {pp83[42]};
    Full_Adder FA_808(s808, c808, in808_1, in808_2, pp81[44]);
    wire[0:0] s809, in809_1, in809_2;
    wire c809;
    assign in809_1 = {pp85[40]};
    assign in809_2 = {pp86[39]};
    Full_Adder FA_809(s809, c809, in809_1, in809_2, pp84[41]);
    wire[0:0] s810, in810_1, in810_2;
    wire c810;
    assign in810_1 = {pp88[37]};
    assign in810_2 = {pp89[36]};
    Full_Adder FA_810(s810, c810, in810_1, in810_2, pp87[38]);
    wire[0:0] s811, in811_1, in811_2;
    wire c811;
    assign in811_1 = {pp91[34]};
    assign in811_2 = {pp92[33]};
    Full_Adder FA_811(s811, c811, in811_1, in811_2, pp90[35]);
    wire[0:0] s812, in812_1, in812_2;
    wire c812;
    assign in812_1 = {pp94[31]};
    assign in812_2 = {pp95[30]};
    Full_Adder FA_812(s812, c812, in812_1, in812_2, pp93[32]);
    wire[0:0] s813, in813_1, in813_2;
    wire c813;
    assign in813_1 = {pp97[28]};
    assign in813_2 = {pp98[27]};
    Full_Adder FA_813(s813, c813, in813_1, in813_2, pp96[29]);
    wire[0:0] s814, in814_1, in814_2;
    wire c814;
    assign in814_1 = {pp100[25]};
    assign in814_2 = {pp101[24]};
    Full_Adder FA_814(s814, c814, in814_1, in814_2, pp99[26]);
    wire[0:0] s815, in815_1, in815_2;
    wire c815;
    assign in815_1 = {pp103[22]};
    assign in815_2 = {pp104[21]};
    Full_Adder FA_815(s815, c815, in815_1, in815_2, pp102[23]);
    wire[0:0] s816, in816_1, in816_2;
    wire c816;
    assign in816_1 = {pp106[19]};
    assign in816_2 = {pp107[18]};
    Full_Adder FA_816(s816, c816, in816_1, in816_2, pp105[20]);
    wire[0:0] s817, in817_1, in817_2;
    wire c817;
    assign in817_1 = {pp109[16]};
    assign in817_2 = {pp110[15]};
    Full_Adder FA_817(s817, c817, in817_1, in817_2, pp108[17]);
    wire[0:0] s818, in818_1, in818_2;
    wire c818;
    assign in818_1 = {pp112[13]};
    assign in818_2 = {pp113[12]};
    Full_Adder FA_818(s818, c818, in818_1, in818_2, pp111[14]);
    wire[0:0] s819, in819_1, in819_2;
    wire c819;
    assign in819_1 = {pp115[10]};
    assign in819_2 = {pp116[9]};
    Full_Adder FA_819(s819, c819, in819_1, in819_2, pp114[11]);
    wire[0:0] s820, in820_1, in820_2;
    wire c820;
    assign in820_1 = {pp117[8]};
    assign in820_2 = {pp118[7]};
    Half_Adder HA_820(s820, c820, in820_1, in820_2);
    wire[0:0] s821, in821_1, in821_2;
    wire c821;
    assign in821_1 = {pp1[125]};
    assign in821_2 = {pp2[124]};
    Full_Adder FA_821(s821, c821, in821_1, in821_2, pp0[126]);
    wire[0:0] s822, in822_1, in822_2;
    wire c822;
    assign in822_1 = {pp4[122]};
    assign in822_2 = {pp5[121]};
    Full_Adder FA_822(s822, c822, in822_1, in822_2, pp3[123]);
    wire[0:0] s823, in823_1, in823_2;
    wire c823;
    assign in823_1 = {pp7[119]};
    assign in823_2 = {pp8[118]};
    Full_Adder FA_823(s823, c823, in823_1, in823_2, pp6[120]);
    wire[0:0] s824, in824_1, in824_2;
    wire c824;
    assign in824_1 = {pp10[116]};
    assign in824_2 = {pp11[115]};
    Full_Adder FA_824(s824, c824, in824_1, in824_2, pp9[117]);
    wire[0:0] s825, in825_1, in825_2;
    wire c825;
    assign in825_1 = {pp13[113]};
    assign in825_2 = {pp14[112]};
    Full_Adder FA_825(s825, c825, in825_1, in825_2, pp12[114]);
    wire[0:0] s826, in826_1, in826_2;
    wire c826;
    assign in826_1 = {pp16[110]};
    assign in826_2 = {pp17[109]};
    Full_Adder FA_826(s826, c826, in826_1, in826_2, pp15[111]);
    wire[0:0] s827, in827_1, in827_2;
    wire c827;
    assign in827_1 = {pp19[107]};
    assign in827_2 = {pp20[106]};
    Full_Adder FA_827(s827, c827, in827_1, in827_2, pp18[108]);
    wire[0:0] s828, in828_1, in828_2;
    wire c828;
    assign in828_1 = {pp22[104]};
    assign in828_2 = {pp23[103]};
    Full_Adder FA_828(s828, c828, in828_1, in828_2, pp21[105]);
    wire[0:0] s829, in829_1, in829_2;
    wire c829;
    assign in829_1 = {pp25[101]};
    assign in829_2 = {pp26[100]};
    Full_Adder FA_829(s829, c829, in829_1, in829_2, pp24[102]);
    wire[0:0] s830, in830_1, in830_2;
    wire c830;
    assign in830_1 = {pp28[98]};
    assign in830_2 = {pp29[97]};
    Full_Adder FA_830(s830, c830, in830_1, in830_2, pp27[99]);
    wire[0:0] s831, in831_1, in831_2;
    wire c831;
    assign in831_1 = {pp31[95]};
    assign in831_2 = {pp32[94]};
    Full_Adder FA_831(s831, c831, in831_1, in831_2, pp30[96]);
    wire[0:0] s832, in832_1, in832_2;
    wire c832;
    assign in832_1 = {pp34[92]};
    assign in832_2 = {pp35[91]};
    Full_Adder FA_832(s832, c832, in832_1, in832_2, pp33[93]);
    wire[0:0] s833, in833_1, in833_2;
    wire c833;
    assign in833_1 = {pp37[89]};
    assign in833_2 = {pp38[88]};
    Full_Adder FA_833(s833, c833, in833_1, in833_2, pp36[90]);
    wire[0:0] s834, in834_1, in834_2;
    wire c834;
    assign in834_1 = {pp40[86]};
    assign in834_2 = {pp41[85]};
    Full_Adder FA_834(s834, c834, in834_1, in834_2, pp39[87]);
    wire[0:0] s835, in835_1, in835_2;
    wire c835;
    assign in835_1 = {pp43[83]};
    assign in835_2 = {pp44[82]};
    Full_Adder FA_835(s835, c835, in835_1, in835_2, pp42[84]);
    wire[0:0] s836, in836_1, in836_2;
    wire c836;
    assign in836_1 = {pp46[80]};
    assign in836_2 = {pp47[79]};
    Full_Adder FA_836(s836, c836, in836_1, in836_2, pp45[81]);
    wire[0:0] s837, in837_1, in837_2;
    wire c837;
    assign in837_1 = {pp49[77]};
    assign in837_2 = {pp50[76]};
    Full_Adder FA_837(s837, c837, in837_1, in837_2, pp48[78]);
    wire[0:0] s838, in838_1, in838_2;
    wire c838;
    assign in838_1 = {pp52[74]};
    assign in838_2 = {pp53[73]};
    Full_Adder FA_838(s838, c838, in838_1, in838_2, pp51[75]);
    wire[0:0] s839, in839_1, in839_2;
    wire c839;
    assign in839_1 = {pp55[71]};
    assign in839_2 = {pp56[70]};
    Full_Adder FA_839(s839, c839, in839_1, in839_2, pp54[72]);
    wire[0:0] s840, in840_1, in840_2;
    wire c840;
    assign in840_1 = {pp58[68]};
    assign in840_2 = {pp59[67]};
    Full_Adder FA_840(s840, c840, in840_1, in840_2, pp57[69]);
    wire[0:0] s841, in841_1, in841_2;
    wire c841;
    assign in841_1 = {pp61[65]};
    assign in841_2 = {pp62[64]};
    Full_Adder FA_841(s841, c841, in841_1, in841_2, pp60[66]);
    wire[0:0] s842, in842_1, in842_2;
    wire c842;
    assign in842_1 = {pp64[62]};
    assign in842_2 = {pp65[61]};
    Full_Adder FA_842(s842, c842, in842_1, in842_2, pp63[63]);
    wire[0:0] s843, in843_1, in843_2;
    wire c843;
    assign in843_1 = {pp67[59]};
    assign in843_2 = {pp68[58]};
    Full_Adder FA_843(s843, c843, in843_1, in843_2, pp66[60]);
    wire[0:0] s844, in844_1, in844_2;
    wire c844;
    assign in844_1 = {pp70[56]};
    assign in844_2 = {pp71[55]};
    Full_Adder FA_844(s844, c844, in844_1, in844_2, pp69[57]);
    wire[0:0] s845, in845_1, in845_2;
    wire c845;
    assign in845_1 = {pp73[53]};
    assign in845_2 = {pp74[52]};
    Full_Adder FA_845(s845, c845, in845_1, in845_2, pp72[54]);
    wire[0:0] s846, in846_1, in846_2;
    wire c846;
    assign in846_1 = {pp76[50]};
    assign in846_2 = {pp77[49]};
    Full_Adder FA_846(s846, c846, in846_1, in846_2, pp75[51]);
    wire[0:0] s847, in847_1, in847_2;
    wire c847;
    assign in847_1 = {pp79[47]};
    assign in847_2 = {pp80[46]};
    Full_Adder FA_847(s847, c847, in847_1, in847_2, pp78[48]);
    wire[0:0] s848, in848_1, in848_2;
    wire c848;
    assign in848_1 = {pp82[44]};
    assign in848_2 = {pp83[43]};
    Full_Adder FA_848(s848, c848, in848_1, in848_2, pp81[45]);
    wire[0:0] s849, in849_1, in849_2;
    wire c849;
    assign in849_1 = {pp85[41]};
    assign in849_2 = {pp86[40]};
    Full_Adder FA_849(s849, c849, in849_1, in849_2, pp84[42]);
    wire[0:0] s850, in850_1, in850_2;
    wire c850;
    assign in850_1 = {pp88[38]};
    assign in850_2 = {pp89[37]};
    Full_Adder FA_850(s850, c850, in850_1, in850_2, pp87[39]);
    wire[0:0] s851, in851_1, in851_2;
    wire c851;
    assign in851_1 = {pp91[35]};
    assign in851_2 = {pp92[34]};
    Full_Adder FA_851(s851, c851, in851_1, in851_2, pp90[36]);
    wire[0:0] s852, in852_1, in852_2;
    wire c852;
    assign in852_1 = {pp94[32]};
    assign in852_2 = {pp95[31]};
    Full_Adder FA_852(s852, c852, in852_1, in852_2, pp93[33]);
    wire[0:0] s853, in853_1, in853_2;
    wire c853;
    assign in853_1 = {pp97[29]};
    assign in853_2 = {pp98[28]};
    Full_Adder FA_853(s853, c853, in853_1, in853_2, pp96[30]);
    wire[0:0] s854, in854_1, in854_2;
    wire c854;
    assign in854_1 = {pp100[26]};
    assign in854_2 = {pp101[25]};
    Full_Adder FA_854(s854, c854, in854_1, in854_2, pp99[27]);
    wire[0:0] s855, in855_1, in855_2;
    wire c855;
    assign in855_1 = {pp103[23]};
    assign in855_2 = {pp104[22]};
    Full_Adder FA_855(s855, c855, in855_1, in855_2, pp102[24]);
    wire[0:0] s856, in856_1, in856_2;
    wire c856;
    assign in856_1 = {pp106[20]};
    assign in856_2 = {pp107[19]};
    Full_Adder FA_856(s856, c856, in856_1, in856_2, pp105[21]);
    wire[0:0] s857, in857_1, in857_2;
    wire c857;
    assign in857_1 = {pp109[17]};
    assign in857_2 = {pp110[16]};
    Full_Adder FA_857(s857, c857, in857_1, in857_2, pp108[18]);
    wire[0:0] s858, in858_1, in858_2;
    wire c858;
    assign in858_1 = {pp112[14]};
    assign in858_2 = {pp113[13]};
    Full_Adder FA_858(s858, c858, in858_1, in858_2, pp111[15]);
    wire[0:0] s859, in859_1, in859_2;
    wire c859;
    assign in859_1 = {pp115[11]};
    assign in859_2 = {pp116[10]};
    Full_Adder FA_859(s859, c859, in859_1, in859_2, pp114[12]);
    wire[0:0] s860, in860_1, in860_2;
    wire c860;
    assign in860_1 = {pp118[8]};
    assign in860_2 = {pp119[7]};
    Full_Adder FA_860(s860, c860, in860_1, in860_2, pp117[9]);
    wire[0:0] s861, in861_1, in861_2;
    wire c861;
    assign in861_1 = {pp120[6]};
    assign in861_2 = {pp121[5]};
    Half_Adder HA_861(s861, c861, in861_1, in861_2);
    wire[0:0] s862, in862_1, in862_2;
    wire c862;
    assign in862_1 = {pp1[126]};
    assign in862_2 = {pp2[125]};
    Full_Adder FA_862(s862, c862, in862_1, in862_2, pp0[127]);
    wire[0:0] s863, in863_1, in863_2;
    wire c863;
    assign in863_1 = {pp4[123]};
    assign in863_2 = {pp5[122]};
    Full_Adder FA_863(s863, c863, in863_1, in863_2, pp3[124]);
    wire[0:0] s864, in864_1, in864_2;
    wire c864;
    assign in864_1 = {pp7[120]};
    assign in864_2 = {pp8[119]};
    Full_Adder FA_864(s864, c864, in864_1, in864_2, pp6[121]);
    wire[0:0] s865, in865_1, in865_2;
    wire c865;
    assign in865_1 = {pp10[117]};
    assign in865_2 = {pp11[116]};
    Full_Adder FA_865(s865, c865, in865_1, in865_2, pp9[118]);
    wire[0:0] s866, in866_1, in866_2;
    wire c866;
    assign in866_1 = {pp13[114]};
    assign in866_2 = {pp14[113]};
    Full_Adder FA_866(s866, c866, in866_1, in866_2, pp12[115]);
    wire[0:0] s867, in867_1, in867_2;
    wire c867;
    assign in867_1 = {pp16[111]};
    assign in867_2 = {pp17[110]};
    Full_Adder FA_867(s867, c867, in867_1, in867_2, pp15[112]);
    wire[0:0] s868, in868_1, in868_2;
    wire c868;
    assign in868_1 = {pp19[108]};
    assign in868_2 = {pp20[107]};
    Full_Adder FA_868(s868, c868, in868_1, in868_2, pp18[109]);
    wire[0:0] s869, in869_1, in869_2;
    wire c869;
    assign in869_1 = {pp22[105]};
    assign in869_2 = {pp23[104]};
    Full_Adder FA_869(s869, c869, in869_1, in869_2, pp21[106]);
    wire[0:0] s870, in870_1, in870_2;
    wire c870;
    assign in870_1 = {pp25[102]};
    assign in870_2 = {pp26[101]};
    Full_Adder FA_870(s870, c870, in870_1, in870_2, pp24[103]);
    wire[0:0] s871, in871_1, in871_2;
    wire c871;
    assign in871_1 = {pp28[99]};
    assign in871_2 = {pp29[98]};
    Full_Adder FA_871(s871, c871, in871_1, in871_2, pp27[100]);
    wire[0:0] s872, in872_1, in872_2;
    wire c872;
    assign in872_1 = {pp31[96]};
    assign in872_2 = {pp32[95]};
    Full_Adder FA_872(s872, c872, in872_1, in872_2, pp30[97]);
    wire[0:0] s873, in873_1, in873_2;
    wire c873;
    assign in873_1 = {pp34[93]};
    assign in873_2 = {pp35[92]};
    Full_Adder FA_873(s873, c873, in873_1, in873_2, pp33[94]);
    wire[0:0] s874, in874_1, in874_2;
    wire c874;
    assign in874_1 = {pp37[90]};
    assign in874_2 = {pp38[89]};
    Full_Adder FA_874(s874, c874, in874_1, in874_2, pp36[91]);
    wire[0:0] s875, in875_1, in875_2;
    wire c875;
    assign in875_1 = {pp40[87]};
    assign in875_2 = {pp41[86]};
    Full_Adder FA_875(s875, c875, in875_1, in875_2, pp39[88]);
    wire[0:0] s876, in876_1, in876_2;
    wire c876;
    assign in876_1 = {pp43[84]};
    assign in876_2 = {pp44[83]};
    Full_Adder FA_876(s876, c876, in876_1, in876_2, pp42[85]);
    wire[0:0] s877, in877_1, in877_2;
    wire c877;
    assign in877_1 = {pp46[81]};
    assign in877_2 = {pp47[80]};
    Full_Adder FA_877(s877, c877, in877_1, in877_2, pp45[82]);
    wire[0:0] s878, in878_1, in878_2;
    wire c878;
    assign in878_1 = {pp49[78]};
    assign in878_2 = {pp50[77]};
    Full_Adder FA_878(s878, c878, in878_1, in878_2, pp48[79]);
    wire[0:0] s879, in879_1, in879_2;
    wire c879;
    assign in879_1 = {pp52[75]};
    assign in879_2 = {pp53[74]};
    Full_Adder FA_879(s879, c879, in879_1, in879_2, pp51[76]);
    wire[0:0] s880, in880_1, in880_2;
    wire c880;
    assign in880_1 = {pp55[72]};
    assign in880_2 = {pp56[71]};
    Full_Adder FA_880(s880, c880, in880_1, in880_2, pp54[73]);
    wire[0:0] s881, in881_1, in881_2;
    wire c881;
    assign in881_1 = {pp58[69]};
    assign in881_2 = {pp59[68]};
    Full_Adder FA_881(s881, c881, in881_1, in881_2, pp57[70]);
    wire[0:0] s882, in882_1, in882_2;
    wire c882;
    assign in882_1 = {pp61[66]};
    assign in882_2 = {pp62[65]};
    Full_Adder FA_882(s882, c882, in882_1, in882_2, pp60[67]);
    wire[0:0] s883, in883_1, in883_2;
    wire c883;
    assign in883_1 = {pp64[63]};
    assign in883_2 = {pp65[62]};
    Full_Adder FA_883(s883, c883, in883_1, in883_2, pp63[64]);
    wire[0:0] s884, in884_1, in884_2;
    wire c884;
    assign in884_1 = {pp67[60]};
    assign in884_2 = {pp68[59]};
    Full_Adder FA_884(s884, c884, in884_1, in884_2, pp66[61]);
    wire[0:0] s885, in885_1, in885_2;
    wire c885;
    assign in885_1 = {pp70[57]};
    assign in885_2 = {pp71[56]};
    Full_Adder FA_885(s885, c885, in885_1, in885_2, pp69[58]);
    wire[0:0] s886, in886_1, in886_2;
    wire c886;
    assign in886_1 = {pp73[54]};
    assign in886_2 = {pp74[53]};
    Full_Adder FA_886(s886, c886, in886_1, in886_2, pp72[55]);
    wire[0:0] s887, in887_1, in887_2;
    wire c887;
    assign in887_1 = {pp76[51]};
    assign in887_2 = {pp77[50]};
    Full_Adder FA_887(s887, c887, in887_1, in887_2, pp75[52]);
    wire[0:0] s888, in888_1, in888_2;
    wire c888;
    assign in888_1 = {pp79[48]};
    assign in888_2 = {pp80[47]};
    Full_Adder FA_888(s888, c888, in888_1, in888_2, pp78[49]);
    wire[0:0] s889, in889_1, in889_2;
    wire c889;
    assign in889_1 = {pp82[45]};
    assign in889_2 = {pp83[44]};
    Full_Adder FA_889(s889, c889, in889_1, in889_2, pp81[46]);
    wire[0:0] s890, in890_1, in890_2;
    wire c890;
    assign in890_1 = {pp85[42]};
    assign in890_2 = {pp86[41]};
    Full_Adder FA_890(s890, c890, in890_1, in890_2, pp84[43]);
    wire[0:0] s891, in891_1, in891_2;
    wire c891;
    assign in891_1 = {pp88[39]};
    assign in891_2 = {pp89[38]};
    Full_Adder FA_891(s891, c891, in891_1, in891_2, pp87[40]);
    wire[0:0] s892, in892_1, in892_2;
    wire c892;
    assign in892_1 = {pp91[36]};
    assign in892_2 = {pp92[35]};
    Full_Adder FA_892(s892, c892, in892_1, in892_2, pp90[37]);
    wire[0:0] s893, in893_1, in893_2;
    wire c893;
    assign in893_1 = {pp94[33]};
    assign in893_2 = {pp95[32]};
    Full_Adder FA_893(s893, c893, in893_1, in893_2, pp93[34]);
    wire[0:0] s894, in894_1, in894_2;
    wire c894;
    assign in894_1 = {pp97[30]};
    assign in894_2 = {pp98[29]};
    Full_Adder FA_894(s894, c894, in894_1, in894_2, pp96[31]);
    wire[0:0] s895, in895_1, in895_2;
    wire c895;
    assign in895_1 = {pp100[27]};
    assign in895_2 = {pp101[26]};
    Full_Adder FA_895(s895, c895, in895_1, in895_2, pp99[28]);
    wire[0:0] s896, in896_1, in896_2;
    wire c896;
    assign in896_1 = {pp103[24]};
    assign in896_2 = {pp104[23]};
    Full_Adder FA_896(s896, c896, in896_1, in896_2, pp102[25]);
    wire[0:0] s897, in897_1, in897_2;
    wire c897;
    assign in897_1 = {pp106[21]};
    assign in897_2 = {pp107[20]};
    Full_Adder FA_897(s897, c897, in897_1, in897_2, pp105[22]);
    wire[0:0] s898, in898_1, in898_2;
    wire c898;
    assign in898_1 = {pp109[18]};
    assign in898_2 = {pp110[17]};
    Full_Adder FA_898(s898, c898, in898_1, in898_2, pp108[19]);
    wire[0:0] s899, in899_1, in899_2;
    wire c899;
    assign in899_1 = {pp112[15]};
    assign in899_2 = {pp113[14]};
    Full_Adder FA_899(s899, c899, in899_1, in899_2, pp111[16]);
    wire[0:0] s900, in900_1, in900_2;
    wire c900;
    assign in900_1 = {pp115[12]};
    assign in900_2 = {pp116[11]};
    Full_Adder FA_900(s900, c900, in900_1, in900_2, pp114[13]);
    wire[0:0] s901, in901_1, in901_2;
    wire c901;
    assign in901_1 = {pp118[9]};
    assign in901_2 = {pp119[8]};
    Full_Adder FA_901(s901, c901, in901_1, in901_2, pp117[10]);
    wire[0:0] s902, in902_1, in902_2;
    wire c902;
    assign in902_1 = {pp121[6]};
    assign in902_2 = {pp122[5]};
    Full_Adder FA_902(s902, c902, in902_1, in902_2, pp120[7]);
    wire[0:0] s903, in903_1, in903_2;
    wire c903;
    assign in903_1 = {pp123[4]};
    assign in903_2 = {pp124[3]};
    Half_Adder HA_903(s903, c903, in903_1, in903_2);
    wire[0:0] s904, in904_1, in904_2;
    wire c904;
    assign in904_1 = {pp2[126]};
    assign in904_2 = {pp3[125]};
    Full_Adder FA_904(s904, c904, in904_1, in904_2, pp1[127]);
    wire[0:0] s905, in905_1, in905_2;
    wire c905;
    assign in905_1 = {pp5[123]};
    assign in905_2 = {pp6[122]};
    Full_Adder FA_905(s905, c905, in905_1, in905_2, pp4[124]);
    wire[0:0] s906, in906_1, in906_2;
    wire c906;
    assign in906_1 = {pp8[120]};
    assign in906_2 = {pp9[119]};
    Full_Adder FA_906(s906, c906, in906_1, in906_2, pp7[121]);
    wire[0:0] s907, in907_1, in907_2;
    wire c907;
    assign in907_1 = {pp11[117]};
    assign in907_2 = {pp12[116]};
    Full_Adder FA_907(s907, c907, in907_1, in907_2, pp10[118]);
    wire[0:0] s908, in908_1, in908_2;
    wire c908;
    assign in908_1 = {pp14[114]};
    assign in908_2 = {pp15[113]};
    Full_Adder FA_908(s908, c908, in908_1, in908_2, pp13[115]);
    wire[0:0] s909, in909_1, in909_2;
    wire c909;
    assign in909_1 = {pp17[111]};
    assign in909_2 = {pp18[110]};
    Full_Adder FA_909(s909, c909, in909_1, in909_2, pp16[112]);
    wire[0:0] s910, in910_1, in910_2;
    wire c910;
    assign in910_1 = {pp20[108]};
    assign in910_2 = {pp21[107]};
    Full_Adder FA_910(s910, c910, in910_1, in910_2, pp19[109]);
    wire[0:0] s911, in911_1, in911_2;
    wire c911;
    assign in911_1 = {pp23[105]};
    assign in911_2 = {pp24[104]};
    Full_Adder FA_911(s911, c911, in911_1, in911_2, pp22[106]);
    wire[0:0] s912, in912_1, in912_2;
    wire c912;
    assign in912_1 = {pp26[102]};
    assign in912_2 = {pp27[101]};
    Full_Adder FA_912(s912, c912, in912_1, in912_2, pp25[103]);
    wire[0:0] s913, in913_1, in913_2;
    wire c913;
    assign in913_1 = {pp29[99]};
    assign in913_2 = {pp30[98]};
    Full_Adder FA_913(s913, c913, in913_1, in913_2, pp28[100]);
    wire[0:0] s914, in914_1, in914_2;
    wire c914;
    assign in914_1 = {pp32[96]};
    assign in914_2 = {pp33[95]};
    Full_Adder FA_914(s914, c914, in914_1, in914_2, pp31[97]);
    wire[0:0] s915, in915_1, in915_2;
    wire c915;
    assign in915_1 = {pp35[93]};
    assign in915_2 = {pp36[92]};
    Full_Adder FA_915(s915, c915, in915_1, in915_2, pp34[94]);
    wire[0:0] s916, in916_1, in916_2;
    wire c916;
    assign in916_1 = {pp38[90]};
    assign in916_2 = {pp39[89]};
    Full_Adder FA_916(s916, c916, in916_1, in916_2, pp37[91]);
    wire[0:0] s917, in917_1, in917_2;
    wire c917;
    assign in917_1 = {pp41[87]};
    assign in917_2 = {pp42[86]};
    Full_Adder FA_917(s917, c917, in917_1, in917_2, pp40[88]);
    wire[0:0] s918, in918_1, in918_2;
    wire c918;
    assign in918_1 = {pp44[84]};
    assign in918_2 = {pp45[83]};
    Full_Adder FA_918(s918, c918, in918_1, in918_2, pp43[85]);
    wire[0:0] s919, in919_1, in919_2;
    wire c919;
    assign in919_1 = {pp47[81]};
    assign in919_2 = {pp48[80]};
    Full_Adder FA_919(s919, c919, in919_1, in919_2, pp46[82]);
    wire[0:0] s920, in920_1, in920_2;
    wire c920;
    assign in920_1 = {pp50[78]};
    assign in920_2 = {pp51[77]};
    Full_Adder FA_920(s920, c920, in920_1, in920_2, pp49[79]);
    wire[0:0] s921, in921_1, in921_2;
    wire c921;
    assign in921_1 = {pp53[75]};
    assign in921_2 = {pp54[74]};
    Full_Adder FA_921(s921, c921, in921_1, in921_2, pp52[76]);
    wire[0:0] s922, in922_1, in922_2;
    wire c922;
    assign in922_1 = {pp56[72]};
    assign in922_2 = {pp57[71]};
    Full_Adder FA_922(s922, c922, in922_1, in922_2, pp55[73]);
    wire[0:0] s923, in923_1, in923_2;
    wire c923;
    assign in923_1 = {pp59[69]};
    assign in923_2 = {pp60[68]};
    Full_Adder FA_923(s923, c923, in923_1, in923_2, pp58[70]);
    wire[0:0] s924, in924_1, in924_2;
    wire c924;
    assign in924_1 = {pp62[66]};
    assign in924_2 = {pp63[65]};
    Full_Adder FA_924(s924, c924, in924_1, in924_2, pp61[67]);
    wire[0:0] s925, in925_1, in925_2;
    wire c925;
    assign in925_1 = {pp65[63]};
    assign in925_2 = {pp66[62]};
    Full_Adder FA_925(s925, c925, in925_1, in925_2, pp64[64]);
    wire[0:0] s926, in926_1, in926_2;
    wire c926;
    assign in926_1 = {pp68[60]};
    assign in926_2 = {pp69[59]};
    Full_Adder FA_926(s926, c926, in926_1, in926_2, pp67[61]);
    wire[0:0] s927, in927_1, in927_2;
    wire c927;
    assign in927_1 = {pp71[57]};
    assign in927_2 = {pp72[56]};
    Full_Adder FA_927(s927, c927, in927_1, in927_2, pp70[58]);
    wire[0:0] s928, in928_1, in928_2;
    wire c928;
    assign in928_1 = {pp74[54]};
    assign in928_2 = {pp75[53]};
    Full_Adder FA_928(s928, c928, in928_1, in928_2, pp73[55]);
    wire[0:0] s929, in929_1, in929_2;
    wire c929;
    assign in929_1 = {pp77[51]};
    assign in929_2 = {pp78[50]};
    Full_Adder FA_929(s929, c929, in929_1, in929_2, pp76[52]);
    wire[0:0] s930, in930_1, in930_2;
    wire c930;
    assign in930_1 = {pp80[48]};
    assign in930_2 = {pp81[47]};
    Full_Adder FA_930(s930, c930, in930_1, in930_2, pp79[49]);
    wire[0:0] s931, in931_1, in931_2;
    wire c931;
    assign in931_1 = {pp83[45]};
    assign in931_2 = {pp84[44]};
    Full_Adder FA_931(s931, c931, in931_1, in931_2, pp82[46]);
    wire[0:0] s932, in932_1, in932_2;
    wire c932;
    assign in932_1 = {pp86[42]};
    assign in932_2 = {pp87[41]};
    Full_Adder FA_932(s932, c932, in932_1, in932_2, pp85[43]);
    wire[0:0] s933, in933_1, in933_2;
    wire c933;
    assign in933_1 = {pp89[39]};
    assign in933_2 = {pp90[38]};
    Full_Adder FA_933(s933, c933, in933_1, in933_2, pp88[40]);
    wire[0:0] s934, in934_1, in934_2;
    wire c934;
    assign in934_1 = {pp92[36]};
    assign in934_2 = {pp93[35]};
    Full_Adder FA_934(s934, c934, in934_1, in934_2, pp91[37]);
    wire[0:0] s935, in935_1, in935_2;
    wire c935;
    assign in935_1 = {pp95[33]};
    assign in935_2 = {pp96[32]};
    Full_Adder FA_935(s935, c935, in935_1, in935_2, pp94[34]);
    wire[0:0] s936, in936_1, in936_2;
    wire c936;
    assign in936_1 = {pp98[30]};
    assign in936_2 = {pp99[29]};
    Full_Adder FA_936(s936, c936, in936_1, in936_2, pp97[31]);
    wire[0:0] s937, in937_1, in937_2;
    wire c937;
    assign in937_1 = {pp101[27]};
    assign in937_2 = {pp102[26]};
    Full_Adder FA_937(s937, c937, in937_1, in937_2, pp100[28]);
    wire[0:0] s938, in938_1, in938_2;
    wire c938;
    assign in938_1 = {pp104[24]};
    assign in938_2 = {pp105[23]};
    Full_Adder FA_938(s938, c938, in938_1, in938_2, pp103[25]);
    wire[0:0] s939, in939_1, in939_2;
    wire c939;
    assign in939_1 = {pp107[21]};
    assign in939_2 = {pp108[20]};
    Full_Adder FA_939(s939, c939, in939_1, in939_2, pp106[22]);
    wire[0:0] s940, in940_1, in940_2;
    wire c940;
    assign in940_1 = {pp110[18]};
    assign in940_2 = {pp111[17]};
    Full_Adder FA_940(s940, c940, in940_1, in940_2, pp109[19]);
    wire[0:0] s941, in941_1, in941_2;
    wire c941;
    assign in941_1 = {pp113[15]};
    assign in941_2 = {pp114[14]};
    Full_Adder FA_941(s941, c941, in941_1, in941_2, pp112[16]);
    wire[0:0] s942, in942_1, in942_2;
    wire c942;
    assign in942_1 = {pp116[12]};
    assign in942_2 = {pp117[11]};
    Full_Adder FA_942(s942, c942, in942_1, in942_2, pp115[13]);
    wire[0:0] s943, in943_1, in943_2;
    wire c943;
    assign in943_1 = {pp119[9]};
    assign in943_2 = {pp120[8]};
    Full_Adder FA_943(s943, c943, in943_1, in943_2, pp118[10]);
    wire[0:0] s944, in944_1, in944_2;
    wire c944;
    assign in944_1 = {pp122[6]};
    assign in944_2 = {pp123[5]};
    Full_Adder FA_944(s944, c944, in944_1, in944_2, pp121[7]);
    wire[0:0] s945, in945_1, in945_2;
    wire c945;
    assign in945_1 = {pp124[4]};
    assign in945_2 = {pp125[3]};
    Half_Adder HA_945(s945, c945, in945_1, in945_2);
    wire[0:0] s946, in946_1, in946_2;
    wire c946;
    assign in946_1 = {pp3[126]};
    assign in946_2 = {pp4[125]};
    Full_Adder FA_946(s946, c946, in946_1, in946_2, pp2[127]);
    wire[0:0] s947, in947_1, in947_2;
    wire c947;
    assign in947_1 = {pp6[123]};
    assign in947_2 = {pp7[122]};
    Full_Adder FA_947(s947, c947, in947_1, in947_2, pp5[124]);
    wire[0:0] s948, in948_1, in948_2;
    wire c948;
    assign in948_1 = {pp9[120]};
    assign in948_2 = {pp10[119]};
    Full_Adder FA_948(s948, c948, in948_1, in948_2, pp8[121]);
    wire[0:0] s949, in949_1, in949_2;
    wire c949;
    assign in949_1 = {pp12[117]};
    assign in949_2 = {pp13[116]};
    Full_Adder FA_949(s949, c949, in949_1, in949_2, pp11[118]);
    wire[0:0] s950, in950_1, in950_2;
    wire c950;
    assign in950_1 = {pp15[114]};
    assign in950_2 = {pp16[113]};
    Full_Adder FA_950(s950, c950, in950_1, in950_2, pp14[115]);
    wire[0:0] s951, in951_1, in951_2;
    wire c951;
    assign in951_1 = {pp18[111]};
    assign in951_2 = {pp19[110]};
    Full_Adder FA_951(s951, c951, in951_1, in951_2, pp17[112]);
    wire[0:0] s952, in952_1, in952_2;
    wire c952;
    assign in952_1 = {pp21[108]};
    assign in952_2 = {pp22[107]};
    Full_Adder FA_952(s952, c952, in952_1, in952_2, pp20[109]);
    wire[0:0] s953, in953_1, in953_2;
    wire c953;
    assign in953_1 = {pp24[105]};
    assign in953_2 = {pp25[104]};
    Full_Adder FA_953(s953, c953, in953_1, in953_2, pp23[106]);
    wire[0:0] s954, in954_1, in954_2;
    wire c954;
    assign in954_1 = {pp27[102]};
    assign in954_2 = {pp28[101]};
    Full_Adder FA_954(s954, c954, in954_1, in954_2, pp26[103]);
    wire[0:0] s955, in955_1, in955_2;
    wire c955;
    assign in955_1 = {pp30[99]};
    assign in955_2 = {pp31[98]};
    Full_Adder FA_955(s955, c955, in955_1, in955_2, pp29[100]);
    wire[0:0] s956, in956_1, in956_2;
    wire c956;
    assign in956_1 = {pp33[96]};
    assign in956_2 = {pp34[95]};
    Full_Adder FA_956(s956, c956, in956_1, in956_2, pp32[97]);
    wire[0:0] s957, in957_1, in957_2;
    wire c957;
    assign in957_1 = {pp36[93]};
    assign in957_2 = {pp37[92]};
    Full_Adder FA_957(s957, c957, in957_1, in957_2, pp35[94]);
    wire[0:0] s958, in958_1, in958_2;
    wire c958;
    assign in958_1 = {pp39[90]};
    assign in958_2 = {pp40[89]};
    Full_Adder FA_958(s958, c958, in958_1, in958_2, pp38[91]);
    wire[0:0] s959, in959_1, in959_2;
    wire c959;
    assign in959_1 = {pp42[87]};
    assign in959_2 = {pp43[86]};
    Full_Adder FA_959(s959, c959, in959_1, in959_2, pp41[88]);
    wire[0:0] s960, in960_1, in960_2;
    wire c960;
    assign in960_1 = {pp45[84]};
    assign in960_2 = {pp46[83]};
    Full_Adder FA_960(s960, c960, in960_1, in960_2, pp44[85]);
    wire[0:0] s961, in961_1, in961_2;
    wire c961;
    assign in961_1 = {pp48[81]};
    assign in961_2 = {pp49[80]};
    Full_Adder FA_961(s961, c961, in961_1, in961_2, pp47[82]);
    wire[0:0] s962, in962_1, in962_2;
    wire c962;
    assign in962_1 = {pp51[78]};
    assign in962_2 = {pp52[77]};
    Full_Adder FA_962(s962, c962, in962_1, in962_2, pp50[79]);
    wire[0:0] s963, in963_1, in963_2;
    wire c963;
    assign in963_1 = {pp54[75]};
    assign in963_2 = {pp55[74]};
    Full_Adder FA_963(s963, c963, in963_1, in963_2, pp53[76]);
    wire[0:0] s964, in964_1, in964_2;
    wire c964;
    assign in964_1 = {pp57[72]};
    assign in964_2 = {pp58[71]};
    Full_Adder FA_964(s964, c964, in964_1, in964_2, pp56[73]);
    wire[0:0] s965, in965_1, in965_2;
    wire c965;
    assign in965_1 = {pp60[69]};
    assign in965_2 = {pp61[68]};
    Full_Adder FA_965(s965, c965, in965_1, in965_2, pp59[70]);
    wire[0:0] s966, in966_1, in966_2;
    wire c966;
    assign in966_1 = {pp63[66]};
    assign in966_2 = {pp64[65]};
    Full_Adder FA_966(s966, c966, in966_1, in966_2, pp62[67]);
    wire[0:0] s967, in967_1, in967_2;
    wire c967;
    assign in967_1 = {pp66[63]};
    assign in967_2 = {pp67[62]};
    Full_Adder FA_967(s967, c967, in967_1, in967_2, pp65[64]);
    wire[0:0] s968, in968_1, in968_2;
    wire c968;
    assign in968_1 = {pp69[60]};
    assign in968_2 = {pp70[59]};
    Full_Adder FA_968(s968, c968, in968_1, in968_2, pp68[61]);
    wire[0:0] s969, in969_1, in969_2;
    wire c969;
    assign in969_1 = {pp72[57]};
    assign in969_2 = {pp73[56]};
    Full_Adder FA_969(s969, c969, in969_1, in969_2, pp71[58]);
    wire[0:0] s970, in970_1, in970_2;
    wire c970;
    assign in970_1 = {pp75[54]};
    assign in970_2 = {pp76[53]};
    Full_Adder FA_970(s970, c970, in970_1, in970_2, pp74[55]);
    wire[0:0] s971, in971_1, in971_2;
    wire c971;
    assign in971_1 = {pp78[51]};
    assign in971_2 = {pp79[50]};
    Full_Adder FA_971(s971, c971, in971_1, in971_2, pp77[52]);
    wire[0:0] s972, in972_1, in972_2;
    wire c972;
    assign in972_1 = {pp81[48]};
    assign in972_2 = {pp82[47]};
    Full_Adder FA_972(s972, c972, in972_1, in972_2, pp80[49]);
    wire[0:0] s973, in973_1, in973_2;
    wire c973;
    assign in973_1 = {pp84[45]};
    assign in973_2 = {pp85[44]};
    Full_Adder FA_973(s973, c973, in973_1, in973_2, pp83[46]);
    wire[0:0] s974, in974_1, in974_2;
    wire c974;
    assign in974_1 = {pp87[42]};
    assign in974_2 = {pp88[41]};
    Full_Adder FA_974(s974, c974, in974_1, in974_2, pp86[43]);
    wire[0:0] s975, in975_1, in975_2;
    wire c975;
    assign in975_1 = {pp90[39]};
    assign in975_2 = {pp91[38]};
    Full_Adder FA_975(s975, c975, in975_1, in975_2, pp89[40]);
    wire[0:0] s976, in976_1, in976_2;
    wire c976;
    assign in976_1 = {pp93[36]};
    assign in976_2 = {pp94[35]};
    Full_Adder FA_976(s976, c976, in976_1, in976_2, pp92[37]);
    wire[0:0] s977, in977_1, in977_2;
    wire c977;
    assign in977_1 = {pp96[33]};
    assign in977_2 = {pp97[32]};
    Full_Adder FA_977(s977, c977, in977_1, in977_2, pp95[34]);
    wire[0:0] s978, in978_1, in978_2;
    wire c978;
    assign in978_1 = {pp99[30]};
    assign in978_2 = {pp100[29]};
    Full_Adder FA_978(s978, c978, in978_1, in978_2, pp98[31]);
    wire[0:0] s979, in979_1, in979_2;
    wire c979;
    assign in979_1 = {pp102[27]};
    assign in979_2 = {pp103[26]};
    Full_Adder FA_979(s979, c979, in979_1, in979_2, pp101[28]);
    wire[0:0] s980, in980_1, in980_2;
    wire c980;
    assign in980_1 = {pp105[24]};
    assign in980_2 = {pp106[23]};
    Full_Adder FA_980(s980, c980, in980_1, in980_2, pp104[25]);
    wire[0:0] s981, in981_1, in981_2;
    wire c981;
    assign in981_1 = {pp108[21]};
    assign in981_2 = {pp109[20]};
    Full_Adder FA_981(s981, c981, in981_1, in981_2, pp107[22]);
    wire[0:0] s982, in982_1, in982_2;
    wire c982;
    assign in982_1 = {pp111[18]};
    assign in982_2 = {pp112[17]};
    Full_Adder FA_982(s982, c982, in982_1, in982_2, pp110[19]);
    wire[0:0] s983, in983_1, in983_2;
    wire c983;
    assign in983_1 = {pp114[15]};
    assign in983_2 = {pp115[14]};
    Full_Adder FA_983(s983, c983, in983_1, in983_2, pp113[16]);
    wire[0:0] s984, in984_1, in984_2;
    wire c984;
    assign in984_1 = {pp117[12]};
    assign in984_2 = {pp118[11]};
    Full_Adder FA_984(s984, c984, in984_1, in984_2, pp116[13]);
    wire[0:0] s985, in985_1, in985_2;
    wire c985;
    assign in985_1 = {pp120[9]};
    assign in985_2 = {pp121[8]};
    Full_Adder FA_985(s985, c985, in985_1, in985_2, pp119[10]);
    wire[0:0] s986, in986_1, in986_2;
    wire c986;
    assign in986_1 = {pp123[6]};
    assign in986_2 = {pp124[5]};
    Full_Adder FA_986(s986, c986, in986_1, in986_2, pp122[7]);
    wire[0:0] s987, in987_1, in987_2;
    wire c987;
    assign in987_1 = {pp4[126]};
    assign in987_2 = {pp5[125]};
    Full_Adder FA_987(s987, c987, in987_1, in987_2, pp3[127]);
    wire[0:0] s988, in988_1, in988_2;
    wire c988;
    assign in988_1 = {pp7[123]};
    assign in988_2 = {pp8[122]};
    Full_Adder FA_988(s988, c988, in988_1, in988_2, pp6[124]);
    wire[0:0] s989, in989_1, in989_2;
    wire c989;
    assign in989_1 = {pp10[120]};
    assign in989_2 = {pp11[119]};
    Full_Adder FA_989(s989, c989, in989_1, in989_2, pp9[121]);
    wire[0:0] s990, in990_1, in990_2;
    wire c990;
    assign in990_1 = {pp13[117]};
    assign in990_2 = {pp14[116]};
    Full_Adder FA_990(s990, c990, in990_1, in990_2, pp12[118]);
    wire[0:0] s991, in991_1, in991_2;
    wire c991;
    assign in991_1 = {pp16[114]};
    assign in991_2 = {pp17[113]};
    Full_Adder FA_991(s991, c991, in991_1, in991_2, pp15[115]);
    wire[0:0] s992, in992_1, in992_2;
    wire c992;
    assign in992_1 = {pp19[111]};
    assign in992_2 = {pp20[110]};
    Full_Adder FA_992(s992, c992, in992_1, in992_2, pp18[112]);
    wire[0:0] s993, in993_1, in993_2;
    wire c993;
    assign in993_1 = {pp22[108]};
    assign in993_2 = {pp23[107]};
    Full_Adder FA_993(s993, c993, in993_1, in993_2, pp21[109]);
    wire[0:0] s994, in994_1, in994_2;
    wire c994;
    assign in994_1 = {pp25[105]};
    assign in994_2 = {pp26[104]};
    Full_Adder FA_994(s994, c994, in994_1, in994_2, pp24[106]);
    wire[0:0] s995, in995_1, in995_2;
    wire c995;
    assign in995_1 = {pp28[102]};
    assign in995_2 = {pp29[101]};
    Full_Adder FA_995(s995, c995, in995_1, in995_2, pp27[103]);
    wire[0:0] s996, in996_1, in996_2;
    wire c996;
    assign in996_1 = {pp31[99]};
    assign in996_2 = {pp32[98]};
    Full_Adder FA_996(s996, c996, in996_1, in996_2, pp30[100]);
    wire[0:0] s997, in997_1, in997_2;
    wire c997;
    assign in997_1 = {pp34[96]};
    assign in997_2 = {pp35[95]};
    Full_Adder FA_997(s997, c997, in997_1, in997_2, pp33[97]);
    wire[0:0] s998, in998_1, in998_2;
    wire c998;
    assign in998_1 = {pp37[93]};
    assign in998_2 = {pp38[92]};
    Full_Adder FA_998(s998, c998, in998_1, in998_2, pp36[94]);
    wire[0:0] s999, in999_1, in999_2;
    wire c999;
    assign in999_1 = {pp40[90]};
    assign in999_2 = {pp41[89]};
    Full_Adder FA_999(s999, c999, in999_1, in999_2, pp39[91]);
    wire[0:0] s1000, in1000_1, in1000_2;
    wire c1000;
    assign in1000_1 = {pp43[87]};
    assign in1000_2 = {pp44[86]};
    Full_Adder FA_1000(s1000, c1000, in1000_1, in1000_2, pp42[88]);
    wire[0:0] s1001, in1001_1, in1001_2;
    wire c1001;
    assign in1001_1 = {pp46[84]};
    assign in1001_2 = {pp47[83]};
    Full_Adder FA_1001(s1001, c1001, in1001_1, in1001_2, pp45[85]);
    wire[0:0] s1002, in1002_1, in1002_2;
    wire c1002;
    assign in1002_1 = {pp49[81]};
    assign in1002_2 = {pp50[80]};
    Full_Adder FA_1002(s1002, c1002, in1002_1, in1002_2, pp48[82]);
    wire[0:0] s1003, in1003_1, in1003_2;
    wire c1003;
    assign in1003_1 = {pp52[78]};
    assign in1003_2 = {pp53[77]};
    Full_Adder FA_1003(s1003, c1003, in1003_1, in1003_2, pp51[79]);
    wire[0:0] s1004, in1004_1, in1004_2;
    wire c1004;
    assign in1004_1 = {pp55[75]};
    assign in1004_2 = {pp56[74]};
    Full_Adder FA_1004(s1004, c1004, in1004_1, in1004_2, pp54[76]);
    wire[0:0] s1005, in1005_1, in1005_2;
    wire c1005;
    assign in1005_1 = {pp58[72]};
    assign in1005_2 = {pp59[71]};
    Full_Adder FA_1005(s1005, c1005, in1005_1, in1005_2, pp57[73]);
    wire[0:0] s1006, in1006_1, in1006_2;
    wire c1006;
    assign in1006_1 = {pp61[69]};
    assign in1006_2 = {pp62[68]};
    Full_Adder FA_1006(s1006, c1006, in1006_1, in1006_2, pp60[70]);
    wire[0:0] s1007, in1007_1, in1007_2;
    wire c1007;
    assign in1007_1 = {pp64[66]};
    assign in1007_2 = {pp65[65]};
    Full_Adder FA_1007(s1007, c1007, in1007_1, in1007_2, pp63[67]);
    wire[0:0] s1008, in1008_1, in1008_2;
    wire c1008;
    assign in1008_1 = {pp67[63]};
    assign in1008_2 = {pp68[62]};
    Full_Adder FA_1008(s1008, c1008, in1008_1, in1008_2, pp66[64]);
    wire[0:0] s1009, in1009_1, in1009_2;
    wire c1009;
    assign in1009_1 = {pp70[60]};
    assign in1009_2 = {pp71[59]};
    Full_Adder FA_1009(s1009, c1009, in1009_1, in1009_2, pp69[61]);
    wire[0:0] s1010, in1010_1, in1010_2;
    wire c1010;
    assign in1010_1 = {pp73[57]};
    assign in1010_2 = {pp74[56]};
    Full_Adder FA_1010(s1010, c1010, in1010_1, in1010_2, pp72[58]);
    wire[0:0] s1011, in1011_1, in1011_2;
    wire c1011;
    assign in1011_1 = {pp76[54]};
    assign in1011_2 = {pp77[53]};
    Full_Adder FA_1011(s1011, c1011, in1011_1, in1011_2, pp75[55]);
    wire[0:0] s1012, in1012_1, in1012_2;
    wire c1012;
    assign in1012_1 = {pp79[51]};
    assign in1012_2 = {pp80[50]};
    Full_Adder FA_1012(s1012, c1012, in1012_1, in1012_2, pp78[52]);
    wire[0:0] s1013, in1013_1, in1013_2;
    wire c1013;
    assign in1013_1 = {pp82[48]};
    assign in1013_2 = {pp83[47]};
    Full_Adder FA_1013(s1013, c1013, in1013_1, in1013_2, pp81[49]);
    wire[0:0] s1014, in1014_1, in1014_2;
    wire c1014;
    assign in1014_1 = {pp85[45]};
    assign in1014_2 = {pp86[44]};
    Full_Adder FA_1014(s1014, c1014, in1014_1, in1014_2, pp84[46]);
    wire[0:0] s1015, in1015_1, in1015_2;
    wire c1015;
    assign in1015_1 = {pp88[42]};
    assign in1015_2 = {pp89[41]};
    Full_Adder FA_1015(s1015, c1015, in1015_1, in1015_2, pp87[43]);
    wire[0:0] s1016, in1016_1, in1016_2;
    wire c1016;
    assign in1016_1 = {pp91[39]};
    assign in1016_2 = {pp92[38]};
    Full_Adder FA_1016(s1016, c1016, in1016_1, in1016_2, pp90[40]);
    wire[0:0] s1017, in1017_1, in1017_2;
    wire c1017;
    assign in1017_1 = {pp94[36]};
    assign in1017_2 = {pp95[35]};
    Full_Adder FA_1017(s1017, c1017, in1017_1, in1017_2, pp93[37]);
    wire[0:0] s1018, in1018_1, in1018_2;
    wire c1018;
    assign in1018_1 = {pp97[33]};
    assign in1018_2 = {pp98[32]};
    Full_Adder FA_1018(s1018, c1018, in1018_1, in1018_2, pp96[34]);
    wire[0:0] s1019, in1019_1, in1019_2;
    wire c1019;
    assign in1019_1 = {pp100[30]};
    assign in1019_2 = {pp101[29]};
    Full_Adder FA_1019(s1019, c1019, in1019_1, in1019_2, pp99[31]);
    wire[0:0] s1020, in1020_1, in1020_2;
    wire c1020;
    assign in1020_1 = {pp103[27]};
    assign in1020_2 = {pp104[26]};
    Full_Adder FA_1020(s1020, c1020, in1020_1, in1020_2, pp102[28]);
    wire[0:0] s1021, in1021_1, in1021_2;
    wire c1021;
    assign in1021_1 = {pp106[24]};
    assign in1021_2 = {pp107[23]};
    Full_Adder FA_1021(s1021, c1021, in1021_1, in1021_2, pp105[25]);
    wire[0:0] s1022, in1022_1, in1022_2;
    wire c1022;
    assign in1022_1 = {pp109[21]};
    assign in1022_2 = {pp110[20]};
    Full_Adder FA_1022(s1022, c1022, in1022_1, in1022_2, pp108[22]);
    wire[0:0] s1023, in1023_1, in1023_2;
    wire c1023;
    assign in1023_1 = {pp112[18]};
    assign in1023_2 = {pp113[17]};
    Full_Adder FA_1023(s1023, c1023, in1023_1, in1023_2, pp111[19]);
    wire[0:0] s1024, in1024_1, in1024_2;
    wire c1024;
    assign in1024_1 = {pp115[15]};
    assign in1024_2 = {pp116[14]};
    Full_Adder FA_1024(s1024, c1024, in1024_1, in1024_2, pp114[16]);
    wire[0:0] s1025, in1025_1, in1025_2;
    wire c1025;
    assign in1025_1 = {pp118[12]};
    assign in1025_2 = {pp119[11]};
    Full_Adder FA_1025(s1025, c1025, in1025_1, in1025_2, pp117[13]);
    wire[0:0] s1026, in1026_1, in1026_2;
    wire c1026;
    assign in1026_1 = {pp121[9]};
    assign in1026_2 = {pp122[8]};
    Full_Adder FA_1026(s1026, c1026, in1026_1, in1026_2, pp120[10]);
    wire[0:0] s1027, in1027_1, in1027_2;
    wire c1027;
    assign in1027_1 = {pp5[126]};
    assign in1027_2 = {pp6[125]};
    Full_Adder FA_1027(s1027, c1027, in1027_1, in1027_2, pp4[127]);
    wire[0:0] s1028, in1028_1, in1028_2;
    wire c1028;
    assign in1028_1 = {pp8[123]};
    assign in1028_2 = {pp9[122]};
    Full_Adder FA_1028(s1028, c1028, in1028_1, in1028_2, pp7[124]);
    wire[0:0] s1029, in1029_1, in1029_2;
    wire c1029;
    assign in1029_1 = {pp11[120]};
    assign in1029_2 = {pp12[119]};
    Full_Adder FA_1029(s1029, c1029, in1029_1, in1029_2, pp10[121]);
    wire[0:0] s1030, in1030_1, in1030_2;
    wire c1030;
    assign in1030_1 = {pp14[117]};
    assign in1030_2 = {pp15[116]};
    Full_Adder FA_1030(s1030, c1030, in1030_1, in1030_2, pp13[118]);
    wire[0:0] s1031, in1031_1, in1031_2;
    wire c1031;
    assign in1031_1 = {pp17[114]};
    assign in1031_2 = {pp18[113]};
    Full_Adder FA_1031(s1031, c1031, in1031_1, in1031_2, pp16[115]);
    wire[0:0] s1032, in1032_1, in1032_2;
    wire c1032;
    assign in1032_1 = {pp20[111]};
    assign in1032_2 = {pp21[110]};
    Full_Adder FA_1032(s1032, c1032, in1032_1, in1032_2, pp19[112]);
    wire[0:0] s1033, in1033_1, in1033_2;
    wire c1033;
    assign in1033_1 = {pp23[108]};
    assign in1033_2 = {pp24[107]};
    Full_Adder FA_1033(s1033, c1033, in1033_1, in1033_2, pp22[109]);
    wire[0:0] s1034, in1034_1, in1034_2;
    wire c1034;
    assign in1034_1 = {pp26[105]};
    assign in1034_2 = {pp27[104]};
    Full_Adder FA_1034(s1034, c1034, in1034_1, in1034_2, pp25[106]);
    wire[0:0] s1035, in1035_1, in1035_2;
    wire c1035;
    assign in1035_1 = {pp29[102]};
    assign in1035_2 = {pp30[101]};
    Full_Adder FA_1035(s1035, c1035, in1035_1, in1035_2, pp28[103]);
    wire[0:0] s1036, in1036_1, in1036_2;
    wire c1036;
    assign in1036_1 = {pp32[99]};
    assign in1036_2 = {pp33[98]};
    Full_Adder FA_1036(s1036, c1036, in1036_1, in1036_2, pp31[100]);
    wire[0:0] s1037, in1037_1, in1037_2;
    wire c1037;
    assign in1037_1 = {pp35[96]};
    assign in1037_2 = {pp36[95]};
    Full_Adder FA_1037(s1037, c1037, in1037_1, in1037_2, pp34[97]);
    wire[0:0] s1038, in1038_1, in1038_2;
    wire c1038;
    assign in1038_1 = {pp38[93]};
    assign in1038_2 = {pp39[92]};
    Full_Adder FA_1038(s1038, c1038, in1038_1, in1038_2, pp37[94]);
    wire[0:0] s1039, in1039_1, in1039_2;
    wire c1039;
    assign in1039_1 = {pp41[90]};
    assign in1039_2 = {pp42[89]};
    Full_Adder FA_1039(s1039, c1039, in1039_1, in1039_2, pp40[91]);
    wire[0:0] s1040, in1040_1, in1040_2;
    wire c1040;
    assign in1040_1 = {pp44[87]};
    assign in1040_2 = {pp45[86]};
    Full_Adder FA_1040(s1040, c1040, in1040_1, in1040_2, pp43[88]);
    wire[0:0] s1041, in1041_1, in1041_2;
    wire c1041;
    assign in1041_1 = {pp47[84]};
    assign in1041_2 = {pp48[83]};
    Full_Adder FA_1041(s1041, c1041, in1041_1, in1041_2, pp46[85]);
    wire[0:0] s1042, in1042_1, in1042_2;
    wire c1042;
    assign in1042_1 = {pp50[81]};
    assign in1042_2 = {pp51[80]};
    Full_Adder FA_1042(s1042, c1042, in1042_1, in1042_2, pp49[82]);
    wire[0:0] s1043, in1043_1, in1043_2;
    wire c1043;
    assign in1043_1 = {pp53[78]};
    assign in1043_2 = {pp54[77]};
    Full_Adder FA_1043(s1043, c1043, in1043_1, in1043_2, pp52[79]);
    wire[0:0] s1044, in1044_1, in1044_2;
    wire c1044;
    assign in1044_1 = {pp56[75]};
    assign in1044_2 = {pp57[74]};
    Full_Adder FA_1044(s1044, c1044, in1044_1, in1044_2, pp55[76]);
    wire[0:0] s1045, in1045_1, in1045_2;
    wire c1045;
    assign in1045_1 = {pp59[72]};
    assign in1045_2 = {pp60[71]};
    Full_Adder FA_1045(s1045, c1045, in1045_1, in1045_2, pp58[73]);
    wire[0:0] s1046, in1046_1, in1046_2;
    wire c1046;
    assign in1046_1 = {pp62[69]};
    assign in1046_2 = {pp63[68]};
    Full_Adder FA_1046(s1046, c1046, in1046_1, in1046_2, pp61[70]);
    wire[0:0] s1047, in1047_1, in1047_2;
    wire c1047;
    assign in1047_1 = {pp65[66]};
    assign in1047_2 = {pp66[65]};
    Full_Adder FA_1047(s1047, c1047, in1047_1, in1047_2, pp64[67]);
    wire[0:0] s1048, in1048_1, in1048_2;
    wire c1048;
    assign in1048_1 = {pp68[63]};
    assign in1048_2 = {pp69[62]};
    Full_Adder FA_1048(s1048, c1048, in1048_1, in1048_2, pp67[64]);
    wire[0:0] s1049, in1049_1, in1049_2;
    wire c1049;
    assign in1049_1 = {pp71[60]};
    assign in1049_2 = {pp72[59]};
    Full_Adder FA_1049(s1049, c1049, in1049_1, in1049_2, pp70[61]);
    wire[0:0] s1050, in1050_1, in1050_2;
    wire c1050;
    assign in1050_1 = {pp74[57]};
    assign in1050_2 = {pp75[56]};
    Full_Adder FA_1050(s1050, c1050, in1050_1, in1050_2, pp73[58]);
    wire[0:0] s1051, in1051_1, in1051_2;
    wire c1051;
    assign in1051_1 = {pp77[54]};
    assign in1051_2 = {pp78[53]};
    Full_Adder FA_1051(s1051, c1051, in1051_1, in1051_2, pp76[55]);
    wire[0:0] s1052, in1052_1, in1052_2;
    wire c1052;
    assign in1052_1 = {pp80[51]};
    assign in1052_2 = {pp81[50]};
    Full_Adder FA_1052(s1052, c1052, in1052_1, in1052_2, pp79[52]);
    wire[0:0] s1053, in1053_1, in1053_2;
    wire c1053;
    assign in1053_1 = {pp83[48]};
    assign in1053_2 = {pp84[47]};
    Full_Adder FA_1053(s1053, c1053, in1053_1, in1053_2, pp82[49]);
    wire[0:0] s1054, in1054_1, in1054_2;
    wire c1054;
    assign in1054_1 = {pp86[45]};
    assign in1054_2 = {pp87[44]};
    Full_Adder FA_1054(s1054, c1054, in1054_1, in1054_2, pp85[46]);
    wire[0:0] s1055, in1055_1, in1055_2;
    wire c1055;
    assign in1055_1 = {pp89[42]};
    assign in1055_2 = {pp90[41]};
    Full_Adder FA_1055(s1055, c1055, in1055_1, in1055_2, pp88[43]);
    wire[0:0] s1056, in1056_1, in1056_2;
    wire c1056;
    assign in1056_1 = {pp92[39]};
    assign in1056_2 = {pp93[38]};
    Full_Adder FA_1056(s1056, c1056, in1056_1, in1056_2, pp91[40]);
    wire[0:0] s1057, in1057_1, in1057_2;
    wire c1057;
    assign in1057_1 = {pp95[36]};
    assign in1057_2 = {pp96[35]};
    Full_Adder FA_1057(s1057, c1057, in1057_1, in1057_2, pp94[37]);
    wire[0:0] s1058, in1058_1, in1058_2;
    wire c1058;
    assign in1058_1 = {pp98[33]};
    assign in1058_2 = {pp99[32]};
    Full_Adder FA_1058(s1058, c1058, in1058_1, in1058_2, pp97[34]);
    wire[0:0] s1059, in1059_1, in1059_2;
    wire c1059;
    assign in1059_1 = {pp101[30]};
    assign in1059_2 = {pp102[29]};
    Full_Adder FA_1059(s1059, c1059, in1059_1, in1059_2, pp100[31]);
    wire[0:0] s1060, in1060_1, in1060_2;
    wire c1060;
    assign in1060_1 = {pp104[27]};
    assign in1060_2 = {pp105[26]};
    Full_Adder FA_1060(s1060, c1060, in1060_1, in1060_2, pp103[28]);
    wire[0:0] s1061, in1061_1, in1061_2;
    wire c1061;
    assign in1061_1 = {pp107[24]};
    assign in1061_2 = {pp108[23]};
    Full_Adder FA_1061(s1061, c1061, in1061_1, in1061_2, pp106[25]);
    wire[0:0] s1062, in1062_1, in1062_2;
    wire c1062;
    assign in1062_1 = {pp110[21]};
    assign in1062_2 = {pp111[20]};
    Full_Adder FA_1062(s1062, c1062, in1062_1, in1062_2, pp109[22]);
    wire[0:0] s1063, in1063_1, in1063_2;
    wire c1063;
    assign in1063_1 = {pp113[18]};
    assign in1063_2 = {pp114[17]};
    Full_Adder FA_1063(s1063, c1063, in1063_1, in1063_2, pp112[19]);
    wire[0:0] s1064, in1064_1, in1064_2;
    wire c1064;
    assign in1064_1 = {pp116[15]};
    assign in1064_2 = {pp117[14]};
    Full_Adder FA_1064(s1064, c1064, in1064_1, in1064_2, pp115[16]);
    wire[0:0] s1065, in1065_1, in1065_2;
    wire c1065;
    assign in1065_1 = {pp119[12]};
    assign in1065_2 = {pp120[11]};
    Full_Adder FA_1065(s1065, c1065, in1065_1, in1065_2, pp118[13]);
    wire[0:0] s1066, in1066_1, in1066_2;
    wire c1066;
    assign in1066_1 = {pp6[126]};
    assign in1066_2 = {pp7[125]};
    Full_Adder FA_1066(s1066, c1066, in1066_1, in1066_2, pp5[127]);
    wire[0:0] s1067, in1067_1, in1067_2;
    wire c1067;
    assign in1067_1 = {pp9[123]};
    assign in1067_2 = {pp10[122]};
    Full_Adder FA_1067(s1067, c1067, in1067_1, in1067_2, pp8[124]);
    wire[0:0] s1068, in1068_1, in1068_2;
    wire c1068;
    assign in1068_1 = {pp12[120]};
    assign in1068_2 = {pp13[119]};
    Full_Adder FA_1068(s1068, c1068, in1068_1, in1068_2, pp11[121]);
    wire[0:0] s1069, in1069_1, in1069_2;
    wire c1069;
    assign in1069_1 = {pp15[117]};
    assign in1069_2 = {pp16[116]};
    Full_Adder FA_1069(s1069, c1069, in1069_1, in1069_2, pp14[118]);
    wire[0:0] s1070, in1070_1, in1070_2;
    wire c1070;
    assign in1070_1 = {pp18[114]};
    assign in1070_2 = {pp19[113]};
    Full_Adder FA_1070(s1070, c1070, in1070_1, in1070_2, pp17[115]);
    wire[0:0] s1071, in1071_1, in1071_2;
    wire c1071;
    assign in1071_1 = {pp21[111]};
    assign in1071_2 = {pp22[110]};
    Full_Adder FA_1071(s1071, c1071, in1071_1, in1071_2, pp20[112]);
    wire[0:0] s1072, in1072_1, in1072_2;
    wire c1072;
    assign in1072_1 = {pp24[108]};
    assign in1072_2 = {pp25[107]};
    Full_Adder FA_1072(s1072, c1072, in1072_1, in1072_2, pp23[109]);
    wire[0:0] s1073, in1073_1, in1073_2;
    wire c1073;
    assign in1073_1 = {pp27[105]};
    assign in1073_2 = {pp28[104]};
    Full_Adder FA_1073(s1073, c1073, in1073_1, in1073_2, pp26[106]);
    wire[0:0] s1074, in1074_1, in1074_2;
    wire c1074;
    assign in1074_1 = {pp30[102]};
    assign in1074_2 = {pp31[101]};
    Full_Adder FA_1074(s1074, c1074, in1074_1, in1074_2, pp29[103]);
    wire[0:0] s1075, in1075_1, in1075_2;
    wire c1075;
    assign in1075_1 = {pp33[99]};
    assign in1075_2 = {pp34[98]};
    Full_Adder FA_1075(s1075, c1075, in1075_1, in1075_2, pp32[100]);
    wire[0:0] s1076, in1076_1, in1076_2;
    wire c1076;
    assign in1076_1 = {pp36[96]};
    assign in1076_2 = {pp37[95]};
    Full_Adder FA_1076(s1076, c1076, in1076_1, in1076_2, pp35[97]);
    wire[0:0] s1077, in1077_1, in1077_2;
    wire c1077;
    assign in1077_1 = {pp39[93]};
    assign in1077_2 = {pp40[92]};
    Full_Adder FA_1077(s1077, c1077, in1077_1, in1077_2, pp38[94]);
    wire[0:0] s1078, in1078_1, in1078_2;
    wire c1078;
    assign in1078_1 = {pp42[90]};
    assign in1078_2 = {pp43[89]};
    Full_Adder FA_1078(s1078, c1078, in1078_1, in1078_2, pp41[91]);
    wire[0:0] s1079, in1079_1, in1079_2;
    wire c1079;
    assign in1079_1 = {pp45[87]};
    assign in1079_2 = {pp46[86]};
    Full_Adder FA_1079(s1079, c1079, in1079_1, in1079_2, pp44[88]);
    wire[0:0] s1080, in1080_1, in1080_2;
    wire c1080;
    assign in1080_1 = {pp48[84]};
    assign in1080_2 = {pp49[83]};
    Full_Adder FA_1080(s1080, c1080, in1080_1, in1080_2, pp47[85]);
    wire[0:0] s1081, in1081_1, in1081_2;
    wire c1081;
    assign in1081_1 = {pp51[81]};
    assign in1081_2 = {pp52[80]};
    Full_Adder FA_1081(s1081, c1081, in1081_1, in1081_2, pp50[82]);
    wire[0:0] s1082, in1082_1, in1082_2;
    wire c1082;
    assign in1082_1 = {pp54[78]};
    assign in1082_2 = {pp55[77]};
    Full_Adder FA_1082(s1082, c1082, in1082_1, in1082_2, pp53[79]);
    wire[0:0] s1083, in1083_1, in1083_2;
    wire c1083;
    assign in1083_1 = {pp57[75]};
    assign in1083_2 = {pp58[74]};
    Full_Adder FA_1083(s1083, c1083, in1083_1, in1083_2, pp56[76]);
    wire[0:0] s1084, in1084_1, in1084_2;
    wire c1084;
    assign in1084_1 = {pp60[72]};
    assign in1084_2 = {pp61[71]};
    Full_Adder FA_1084(s1084, c1084, in1084_1, in1084_2, pp59[73]);
    wire[0:0] s1085, in1085_1, in1085_2;
    wire c1085;
    assign in1085_1 = {pp63[69]};
    assign in1085_2 = {pp64[68]};
    Full_Adder FA_1085(s1085, c1085, in1085_1, in1085_2, pp62[70]);
    wire[0:0] s1086, in1086_1, in1086_2;
    wire c1086;
    assign in1086_1 = {pp66[66]};
    assign in1086_2 = {pp67[65]};
    Full_Adder FA_1086(s1086, c1086, in1086_1, in1086_2, pp65[67]);
    wire[0:0] s1087, in1087_1, in1087_2;
    wire c1087;
    assign in1087_1 = {pp69[63]};
    assign in1087_2 = {pp70[62]};
    Full_Adder FA_1087(s1087, c1087, in1087_1, in1087_2, pp68[64]);
    wire[0:0] s1088, in1088_1, in1088_2;
    wire c1088;
    assign in1088_1 = {pp72[60]};
    assign in1088_2 = {pp73[59]};
    Full_Adder FA_1088(s1088, c1088, in1088_1, in1088_2, pp71[61]);
    wire[0:0] s1089, in1089_1, in1089_2;
    wire c1089;
    assign in1089_1 = {pp75[57]};
    assign in1089_2 = {pp76[56]};
    Full_Adder FA_1089(s1089, c1089, in1089_1, in1089_2, pp74[58]);
    wire[0:0] s1090, in1090_1, in1090_2;
    wire c1090;
    assign in1090_1 = {pp78[54]};
    assign in1090_2 = {pp79[53]};
    Full_Adder FA_1090(s1090, c1090, in1090_1, in1090_2, pp77[55]);
    wire[0:0] s1091, in1091_1, in1091_2;
    wire c1091;
    assign in1091_1 = {pp81[51]};
    assign in1091_2 = {pp82[50]};
    Full_Adder FA_1091(s1091, c1091, in1091_1, in1091_2, pp80[52]);
    wire[0:0] s1092, in1092_1, in1092_2;
    wire c1092;
    assign in1092_1 = {pp84[48]};
    assign in1092_2 = {pp85[47]};
    Full_Adder FA_1092(s1092, c1092, in1092_1, in1092_2, pp83[49]);
    wire[0:0] s1093, in1093_1, in1093_2;
    wire c1093;
    assign in1093_1 = {pp87[45]};
    assign in1093_2 = {pp88[44]};
    Full_Adder FA_1093(s1093, c1093, in1093_1, in1093_2, pp86[46]);
    wire[0:0] s1094, in1094_1, in1094_2;
    wire c1094;
    assign in1094_1 = {pp90[42]};
    assign in1094_2 = {pp91[41]};
    Full_Adder FA_1094(s1094, c1094, in1094_1, in1094_2, pp89[43]);
    wire[0:0] s1095, in1095_1, in1095_2;
    wire c1095;
    assign in1095_1 = {pp93[39]};
    assign in1095_2 = {pp94[38]};
    Full_Adder FA_1095(s1095, c1095, in1095_1, in1095_2, pp92[40]);
    wire[0:0] s1096, in1096_1, in1096_2;
    wire c1096;
    assign in1096_1 = {pp96[36]};
    assign in1096_2 = {pp97[35]};
    Full_Adder FA_1096(s1096, c1096, in1096_1, in1096_2, pp95[37]);
    wire[0:0] s1097, in1097_1, in1097_2;
    wire c1097;
    assign in1097_1 = {pp99[33]};
    assign in1097_2 = {pp100[32]};
    Full_Adder FA_1097(s1097, c1097, in1097_1, in1097_2, pp98[34]);
    wire[0:0] s1098, in1098_1, in1098_2;
    wire c1098;
    assign in1098_1 = {pp102[30]};
    assign in1098_2 = {pp103[29]};
    Full_Adder FA_1098(s1098, c1098, in1098_1, in1098_2, pp101[31]);
    wire[0:0] s1099, in1099_1, in1099_2;
    wire c1099;
    assign in1099_1 = {pp105[27]};
    assign in1099_2 = {pp106[26]};
    Full_Adder FA_1099(s1099, c1099, in1099_1, in1099_2, pp104[28]);
    wire[0:0] s1100, in1100_1, in1100_2;
    wire c1100;
    assign in1100_1 = {pp108[24]};
    assign in1100_2 = {pp109[23]};
    Full_Adder FA_1100(s1100, c1100, in1100_1, in1100_2, pp107[25]);
    wire[0:0] s1101, in1101_1, in1101_2;
    wire c1101;
    assign in1101_1 = {pp111[21]};
    assign in1101_2 = {pp112[20]};
    Full_Adder FA_1101(s1101, c1101, in1101_1, in1101_2, pp110[22]);
    wire[0:0] s1102, in1102_1, in1102_2;
    wire c1102;
    assign in1102_1 = {pp114[18]};
    assign in1102_2 = {pp115[17]};
    Full_Adder FA_1102(s1102, c1102, in1102_1, in1102_2, pp113[19]);
    wire[0:0] s1103, in1103_1, in1103_2;
    wire c1103;
    assign in1103_1 = {pp117[15]};
    assign in1103_2 = {pp118[14]};
    Full_Adder FA_1103(s1103, c1103, in1103_1, in1103_2, pp116[16]);
    wire[0:0] s1104, in1104_1, in1104_2;
    wire c1104;
    assign in1104_1 = {pp7[126]};
    assign in1104_2 = {pp8[125]};
    Full_Adder FA_1104(s1104, c1104, in1104_1, in1104_2, pp6[127]);
    wire[0:0] s1105, in1105_1, in1105_2;
    wire c1105;
    assign in1105_1 = {pp10[123]};
    assign in1105_2 = {pp11[122]};
    Full_Adder FA_1105(s1105, c1105, in1105_1, in1105_2, pp9[124]);
    wire[0:0] s1106, in1106_1, in1106_2;
    wire c1106;
    assign in1106_1 = {pp13[120]};
    assign in1106_2 = {pp14[119]};
    Full_Adder FA_1106(s1106, c1106, in1106_1, in1106_2, pp12[121]);
    wire[0:0] s1107, in1107_1, in1107_2;
    wire c1107;
    assign in1107_1 = {pp16[117]};
    assign in1107_2 = {pp17[116]};
    Full_Adder FA_1107(s1107, c1107, in1107_1, in1107_2, pp15[118]);
    wire[0:0] s1108, in1108_1, in1108_2;
    wire c1108;
    assign in1108_1 = {pp19[114]};
    assign in1108_2 = {pp20[113]};
    Full_Adder FA_1108(s1108, c1108, in1108_1, in1108_2, pp18[115]);
    wire[0:0] s1109, in1109_1, in1109_2;
    wire c1109;
    assign in1109_1 = {pp22[111]};
    assign in1109_2 = {pp23[110]};
    Full_Adder FA_1109(s1109, c1109, in1109_1, in1109_2, pp21[112]);
    wire[0:0] s1110, in1110_1, in1110_2;
    wire c1110;
    assign in1110_1 = {pp25[108]};
    assign in1110_2 = {pp26[107]};
    Full_Adder FA_1110(s1110, c1110, in1110_1, in1110_2, pp24[109]);
    wire[0:0] s1111, in1111_1, in1111_2;
    wire c1111;
    assign in1111_1 = {pp28[105]};
    assign in1111_2 = {pp29[104]};
    Full_Adder FA_1111(s1111, c1111, in1111_1, in1111_2, pp27[106]);
    wire[0:0] s1112, in1112_1, in1112_2;
    wire c1112;
    assign in1112_1 = {pp31[102]};
    assign in1112_2 = {pp32[101]};
    Full_Adder FA_1112(s1112, c1112, in1112_1, in1112_2, pp30[103]);
    wire[0:0] s1113, in1113_1, in1113_2;
    wire c1113;
    assign in1113_1 = {pp34[99]};
    assign in1113_2 = {pp35[98]};
    Full_Adder FA_1113(s1113, c1113, in1113_1, in1113_2, pp33[100]);
    wire[0:0] s1114, in1114_1, in1114_2;
    wire c1114;
    assign in1114_1 = {pp37[96]};
    assign in1114_2 = {pp38[95]};
    Full_Adder FA_1114(s1114, c1114, in1114_1, in1114_2, pp36[97]);
    wire[0:0] s1115, in1115_1, in1115_2;
    wire c1115;
    assign in1115_1 = {pp40[93]};
    assign in1115_2 = {pp41[92]};
    Full_Adder FA_1115(s1115, c1115, in1115_1, in1115_2, pp39[94]);
    wire[0:0] s1116, in1116_1, in1116_2;
    wire c1116;
    assign in1116_1 = {pp43[90]};
    assign in1116_2 = {pp44[89]};
    Full_Adder FA_1116(s1116, c1116, in1116_1, in1116_2, pp42[91]);
    wire[0:0] s1117, in1117_1, in1117_2;
    wire c1117;
    assign in1117_1 = {pp46[87]};
    assign in1117_2 = {pp47[86]};
    Full_Adder FA_1117(s1117, c1117, in1117_1, in1117_2, pp45[88]);
    wire[0:0] s1118, in1118_1, in1118_2;
    wire c1118;
    assign in1118_1 = {pp49[84]};
    assign in1118_2 = {pp50[83]};
    Full_Adder FA_1118(s1118, c1118, in1118_1, in1118_2, pp48[85]);
    wire[0:0] s1119, in1119_1, in1119_2;
    wire c1119;
    assign in1119_1 = {pp52[81]};
    assign in1119_2 = {pp53[80]};
    Full_Adder FA_1119(s1119, c1119, in1119_1, in1119_2, pp51[82]);
    wire[0:0] s1120, in1120_1, in1120_2;
    wire c1120;
    assign in1120_1 = {pp55[78]};
    assign in1120_2 = {pp56[77]};
    Full_Adder FA_1120(s1120, c1120, in1120_1, in1120_2, pp54[79]);
    wire[0:0] s1121, in1121_1, in1121_2;
    wire c1121;
    assign in1121_1 = {pp58[75]};
    assign in1121_2 = {pp59[74]};
    Full_Adder FA_1121(s1121, c1121, in1121_1, in1121_2, pp57[76]);
    wire[0:0] s1122, in1122_1, in1122_2;
    wire c1122;
    assign in1122_1 = {pp61[72]};
    assign in1122_2 = {pp62[71]};
    Full_Adder FA_1122(s1122, c1122, in1122_1, in1122_2, pp60[73]);
    wire[0:0] s1123, in1123_1, in1123_2;
    wire c1123;
    assign in1123_1 = {pp64[69]};
    assign in1123_2 = {pp65[68]};
    Full_Adder FA_1123(s1123, c1123, in1123_1, in1123_2, pp63[70]);
    wire[0:0] s1124, in1124_1, in1124_2;
    wire c1124;
    assign in1124_1 = {pp67[66]};
    assign in1124_2 = {pp68[65]};
    Full_Adder FA_1124(s1124, c1124, in1124_1, in1124_2, pp66[67]);
    wire[0:0] s1125, in1125_1, in1125_2;
    wire c1125;
    assign in1125_1 = {pp70[63]};
    assign in1125_2 = {pp71[62]};
    Full_Adder FA_1125(s1125, c1125, in1125_1, in1125_2, pp69[64]);
    wire[0:0] s1126, in1126_1, in1126_2;
    wire c1126;
    assign in1126_1 = {pp73[60]};
    assign in1126_2 = {pp74[59]};
    Full_Adder FA_1126(s1126, c1126, in1126_1, in1126_2, pp72[61]);
    wire[0:0] s1127, in1127_1, in1127_2;
    wire c1127;
    assign in1127_1 = {pp76[57]};
    assign in1127_2 = {pp77[56]};
    Full_Adder FA_1127(s1127, c1127, in1127_1, in1127_2, pp75[58]);
    wire[0:0] s1128, in1128_1, in1128_2;
    wire c1128;
    assign in1128_1 = {pp79[54]};
    assign in1128_2 = {pp80[53]};
    Full_Adder FA_1128(s1128, c1128, in1128_1, in1128_2, pp78[55]);
    wire[0:0] s1129, in1129_1, in1129_2;
    wire c1129;
    assign in1129_1 = {pp82[51]};
    assign in1129_2 = {pp83[50]};
    Full_Adder FA_1129(s1129, c1129, in1129_1, in1129_2, pp81[52]);
    wire[0:0] s1130, in1130_1, in1130_2;
    wire c1130;
    assign in1130_1 = {pp85[48]};
    assign in1130_2 = {pp86[47]};
    Full_Adder FA_1130(s1130, c1130, in1130_1, in1130_2, pp84[49]);
    wire[0:0] s1131, in1131_1, in1131_2;
    wire c1131;
    assign in1131_1 = {pp88[45]};
    assign in1131_2 = {pp89[44]};
    Full_Adder FA_1131(s1131, c1131, in1131_1, in1131_2, pp87[46]);
    wire[0:0] s1132, in1132_1, in1132_2;
    wire c1132;
    assign in1132_1 = {pp91[42]};
    assign in1132_2 = {pp92[41]};
    Full_Adder FA_1132(s1132, c1132, in1132_1, in1132_2, pp90[43]);
    wire[0:0] s1133, in1133_1, in1133_2;
    wire c1133;
    assign in1133_1 = {pp94[39]};
    assign in1133_2 = {pp95[38]};
    Full_Adder FA_1133(s1133, c1133, in1133_1, in1133_2, pp93[40]);
    wire[0:0] s1134, in1134_1, in1134_2;
    wire c1134;
    assign in1134_1 = {pp97[36]};
    assign in1134_2 = {pp98[35]};
    Full_Adder FA_1134(s1134, c1134, in1134_1, in1134_2, pp96[37]);
    wire[0:0] s1135, in1135_1, in1135_2;
    wire c1135;
    assign in1135_1 = {pp100[33]};
    assign in1135_2 = {pp101[32]};
    Full_Adder FA_1135(s1135, c1135, in1135_1, in1135_2, pp99[34]);
    wire[0:0] s1136, in1136_1, in1136_2;
    wire c1136;
    assign in1136_1 = {pp103[30]};
    assign in1136_2 = {pp104[29]};
    Full_Adder FA_1136(s1136, c1136, in1136_1, in1136_2, pp102[31]);
    wire[0:0] s1137, in1137_1, in1137_2;
    wire c1137;
    assign in1137_1 = {pp106[27]};
    assign in1137_2 = {pp107[26]};
    Full_Adder FA_1137(s1137, c1137, in1137_1, in1137_2, pp105[28]);
    wire[0:0] s1138, in1138_1, in1138_2;
    wire c1138;
    assign in1138_1 = {pp109[24]};
    assign in1138_2 = {pp110[23]};
    Full_Adder FA_1138(s1138, c1138, in1138_1, in1138_2, pp108[25]);
    wire[0:0] s1139, in1139_1, in1139_2;
    wire c1139;
    assign in1139_1 = {pp112[21]};
    assign in1139_2 = {pp113[20]};
    Full_Adder FA_1139(s1139, c1139, in1139_1, in1139_2, pp111[22]);
    wire[0:0] s1140, in1140_1, in1140_2;
    wire c1140;
    assign in1140_1 = {pp115[18]};
    assign in1140_2 = {pp116[17]};
    Full_Adder FA_1140(s1140, c1140, in1140_1, in1140_2, pp114[19]);
    wire[0:0] s1141, in1141_1, in1141_2;
    wire c1141;
    assign in1141_1 = {pp8[126]};
    assign in1141_2 = {pp9[125]};
    Full_Adder FA_1141(s1141, c1141, in1141_1, in1141_2, pp7[127]);
    wire[0:0] s1142, in1142_1, in1142_2;
    wire c1142;
    assign in1142_1 = {pp11[123]};
    assign in1142_2 = {pp12[122]};
    Full_Adder FA_1142(s1142, c1142, in1142_1, in1142_2, pp10[124]);
    wire[0:0] s1143, in1143_1, in1143_2;
    wire c1143;
    assign in1143_1 = {pp14[120]};
    assign in1143_2 = {pp15[119]};
    Full_Adder FA_1143(s1143, c1143, in1143_1, in1143_2, pp13[121]);
    wire[0:0] s1144, in1144_1, in1144_2;
    wire c1144;
    assign in1144_1 = {pp17[117]};
    assign in1144_2 = {pp18[116]};
    Full_Adder FA_1144(s1144, c1144, in1144_1, in1144_2, pp16[118]);
    wire[0:0] s1145, in1145_1, in1145_2;
    wire c1145;
    assign in1145_1 = {pp20[114]};
    assign in1145_2 = {pp21[113]};
    Full_Adder FA_1145(s1145, c1145, in1145_1, in1145_2, pp19[115]);
    wire[0:0] s1146, in1146_1, in1146_2;
    wire c1146;
    assign in1146_1 = {pp23[111]};
    assign in1146_2 = {pp24[110]};
    Full_Adder FA_1146(s1146, c1146, in1146_1, in1146_2, pp22[112]);
    wire[0:0] s1147, in1147_1, in1147_2;
    wire c1147;
    assign in1147_1 = {pp26[108]};
    assign in1147_2 = {pp27[107]};
    Full_Adder FA_1147(s1147, c1147, in1147_1, in1147_2, pp25[109]);
    wire[0:0] s1148, in1148_1, in1148_2;
    wire c1148;
    assign in1148_1 = {pp29[105]};
    assign in1148_2 = {pp30[104]};
    Full_Adder FA_1148(s1148, c1148, in1148_1, in1148_2, pp28[106]);
    wire[0:0] s1149, in1149_1, in1149_2;
    wire c1149;
    assign in1149_1 = {pp32[102]};
    assign in1149_2 = {pp33[101]};
    Full_Adder FA_1149(s1149, c1149, in1149_1, in1149_2, pp31[103]);
    wire[0:0] s1150, in1150_1, in1150_2;
    wire c1150;
    assign in1150_1 = {pp35[99]};
    assign in1150_2 = {pp36[98]};
    Full_Adder FA_1150(s1150, c1150, in1150_1, in1150_2, pp34[100]);
    wire[0:0] s1151, in1151_1, in1151_2;
    wire c1151;
    assign in1151_1 = {pp38[96]};
    assign in1151_2 = {pp39[95]};
    Full_Adder FA_1151(s1151, c1151, in1151_1, in1151_2, pp37[97]);
    wire[0:0] s1152, in1152_1, in1152_2;
    wire c1152;
    assign in1152_1 = {pp41[93]};
    assign in1152_2 = {pp42[92]};
    Full_Adder FA_1152(s1152, c1152, in1152_1, in1152_2, pp40[94]);
    wire[0:0] s1153, in1153_1, in1153_2;
    wire c1153;
    assign in1153_1 = {pp44[90]};
    assign in1153_2 = {pp45[89]};
    Full_Adder FA_1153(s1153, c1153, in1153_1, in1153_2, pp43[91]);
    wire[0:0] s1154, in1154_1, in1154_2;
    wire c1154;
    assign in1154_1 = {pp47[87]};
    assign in1154_2 = {pp48[86]};
    Full_Adder FA_1154(s1154, c1154, in1154_1, in1154_2, pp46[88]);
    wire[0:0] s1155, in1155_1, in1155_2;
    wire c1155;
    assign in1155_1 = {pp50[84]};
    assign in1155_2 = {pp51[83]};
    Full_Adder FA_1155(s1155, c1155, in1155_1, in1155_2, pp49[85]);
    wire[0:0] s1156, in1156_1, in1156_2;
    wire c1156;
    assign in1156_1 = {pp53[81]};
    assign in1156_2 = {pp54[80]};
    Full_Adder FA_1156(s1156, c1156, in1156_1, in1156_2, pp52[82]);
    wire[0:0] s1157, in1157_1, in1157_2;
    wire c1157;
    assign in1157_1 = {pp56[78]};
    assign in1157_2 = {pp57[77]};
    Full_Adder FA_1157(s1157, c1157, in1157_1, in1157_2, pp55[79]);
    wire[0:0] s1158, in1158_1, in1158_2;
    wire c1158;
    assign in1158_1 = {pp59[75]};
    assign in1158_2 = {pp60[74]};
    Full_Adder FA_1158(s1158, c1158, in1158_1, in1158_2, pp58[76]);
    wire[0:0] s1159, in1159_1, in1159_2;
    wire c1159;
    assign in1159_1 = {pp62[72]};
    assign in1159_2 = {pp63[71]};
    Full_Adder FA_1159(s1159, c1159, in1159_1, in1159_2, pp61[73]);
    wire[0:0] s1160, in1160_1, in1160_2;
    wire c1160;
    assign in1160_1 = {pp65[69]};
    assign in1160_2 = {pp66[68]};
    Full_Adder FA_1160(s1160, c1160, in1160_1, in1160_2, pp64[70]);
    wire[0:0] s1161, in1161_1, in1161_2;
    wire c1161;
    assign in1161_1 = {pp68[66]};
    assign in1161_2 = {pp69[65]};
    Full_Adder FA_1161(s1161, c1161, in1161_1, in1161_2, pp67[67]);
    wire[0:0] s1162, in1162_1, in1162_2;
    wire c1162;
    assign in1162_1 = {pp71[63]};
    assign in1162_2 = {pp72[62]};
    Full_Adder FA_1162(s1162, c1162, in1162_1, in1162_2, pp70[64]);
    wire[0:0] s1163, in1163_1, in1163_2;
    wire c1163;
    assign in1163_1 = {pp74[60]};
    assign in1163_2 = {pp75[59]};
    Full_Adder FA_1163(s1163, c1163, in1163_1, in1163_2, pp73[61]);
    wire[0:0] s1164, in1164_1, in1164_2;
    wire c1164;
    assign in1164_1 = {pp77[57]};
    assign in1164_2 = {pp78[56]};
    Full_Adder FA_1164(s1164, c1164, in1164_1, in1164_2, pp76[58]);
    wire[0:0] s1165, in1165_1, in1165_2;
    wire c1165;
    assign in1165_1 = {pp80[54]};
    assign in1165_2 = {pp81[53]};
    Full_Adder FA_1165(s1165, c1165, in1165_1, in1165_2, pp79[55]);
    wire[0:0] s1166, in1166_1, in1166_2;
    wire c1166;
    assign in1166_1 = {pp83[51]};
    assign in1166_2 = {pp84[50]};
    Full_Adder FA_1166(s1166, c1166, in1166_1, in1166_2, pp82[52]);
    wire[0:0] s1167, in1167_1, in1167_2;
    wire c1167;
    assign in1167_1 = {pp86[48]};
    assign in1167_2 = {pp87[47]};
    Full_Adder FA_1167(s1167, c1167, in1167_1, in1167_2, pp85[49]);
    wire[0:0] s1168, in1168_1, in1168_2;
    wire c1168;
    assign in1168_1 = {pp89[45]};
    assign in1168_2 = {pp90[44]};
    Full_Adder FA_1168(s1168, c1168, in1168_1, in1168_2, pp88[46]);
    wire[0:0] s1169, in1169_1, in1169_2;
    wire c1169;
    assign in1169_1 = {pp92[42]};
    assign in1169_2 = {pp93[41]};
    Full_Adder FA_1169(s1169, c1169, in1169_1, in1169_2, pp91[43]);
    wire[0:0] s1170, in1170_1, in1170_2;
    wire c1170;
    assign in1170_1 = {pp95[39]};
    assign in1170_2 = {pp96[38]};
    Full_Adder FA_1170(s1170, c1170, in1170_1, in1170_2, pp94[40]);
    wire[0:0] s1171, in1171_1, in1171_2;
    wire c1171;
    assign in1171_1 = {pp98[36]};
    assign in1171_2 = {pp99[35]};
    Full_Adder FA_1171(s1171, c1171, in1171_1, in1171_2, pp97[37]);
    wire[0:0] s1172, in1172_1, in1172_2;
    wire c1172;
    assign in1172_1 = {pp101[33]};
    assign in1172_2 = {pp102[32]};
    Full_Adder FA_1172(s1172, c1172, in1172_1, in1172_2, pp100[34]);
    wire[0:0] s1173, in1173_1, in1173_2;
    wire c1173;
    assign in1173_1 = {pp104[30]};
    assign in1173_2 = {pp105[29]};
    Full_Adder FA_1173(s1173, c1173, in1173_1, in1173_2, pp103[31]);
    wire[0:0] s1174, in1174_1, in1174_2;
    wire c1174;
    assign in1174_1 = {pp107[27]};
    assign in1174_2 = {pp108[26]};
    Full_Adder FA_1174(s1174, c1174, in1174_1, in1174_2, pp106[28]);
    wire[0:0] s1175, in1175_1, in1175_2;
    wire c1175;
    assign in1175_1 = {pp110[24]};
    assign in1175_2 = {pp111[23]};
    Full_Adder FA_1175(s1175, c1175, in1175_1, in1175_2, pp109[25]);
    wire[0:0] s1176, in1176_1, in1176_2;
    wire c1176;
    assign in1176_1 = {pp113[21]};
    assign in1176_2 = {pp114[20]};
    Full_Adder FA_1176(s1176, c1176, in1176_1, in1176_2, pp112[22]);
    wire[0:0] s1177, in1177_1, in1177_2;
    wire c1177;
    assign in1177_1 = {pp9[126]};
    assign in1177_2 = {pp10[125]};
    Full_Adder FA_1177(s1177, c1177, in1177_1, in1177_2, pp8[127]);
    wire[0:0] s1178, in1178_1, in1178_2;
    wire c1178;
    assign in1178_1 = {pp12[123]};
    assign in1178_2 = {pp13[122]};
    Full_Adder FA_1178(s1178, c1178, in1178_1, in1178_2, pp11[124]);
    wire[0:0] s1179, in1179_1, in1179_2;
    wire c1179;
    assign in1179_1 = {pp15[120]};
    assign in1179_2 = {pp16[119]};
    Full_Adder FA_1179(s1179, c1179, in1179_1, in1179_2, pp14[121]);
    wire[0:0] s1180, in1180_1, in1180_2;
    wire c1180;
    assign in1180_1 = {pp18[117]};
    assign in1180_2 = {pp19[116]};
    Full_Adder FA_1180(s1180, c1180, in1180_1, in1180_2, pp17[118]);
    wire[0:0] s1181, in1181_1, in1181_2;
    wire c1181;
    assign in1181_1 = {pp21[114]};
    assign in1181_2 = {pp22[113]};
    Full_Adder FA_1181(s1181, c1181, in1181_1, in1181_2, pp20[115]);
    wire[0:0] s1182, in1182_1, in1182_2;
    wire c1182;
    assign in1182_1 = {pp24[111]};
    assign in1182_2 = {pp25[110]};
    Full_Adder FA_1182(s1182, c1182, in1182_1, in1182_2, pp23[112]);
    wire[0:0] s1183, in1183_1, in1183_2;
    wire c1183;
    assign in1183_1 = {pp27[108]};
    assign in1183_2 = {pp28[107]};
    Full_Adder FA_1183(s1183, c1183, in1183_1, in1183_2, pp26[109]);
    wire[0:0] s1184, in1184_1, in1184_2;
    wire c1184;
    assign in1184_1 = {pp30[105]};
    assign in1184_2 = {pp31[104]};
    Full_Adder FA_1184(s1184, c1184, in1184_1, in1184_2, pp29[106]);
    wire[0:0] s1185, in1185_1, in1185_2;
    wire c1185;
    assign in1185_1 = {pp33[102]};
    assign in1185_2 = {pp34[101]};
    Full_Adder FA_1185(s1185, c1185, in1185_1, in1185_2, pp32[103]);
    wire[0:0] s1186, in1186_1, in1186_2;
    wire c1186;
    assign in1186_1 = {pp36[99]};
    assign in1186_2 = {pp37[98]};
    Full_Adder FA_1186(s1186, c1186, in1186_1, in1186_2, pp35[100]);
    wire[0:0] s1187, in1187_1, in1187_2;
    wire c1187;
    assign in1187_1 = {pp39[96]};
    assign in1187_2 = {pp40[95]};
    Full_Adder FA_1187(s1187, c1187, in1187_1, in1187_2, pp38[97]);
    wire[0:0] s1188, in1188_1, in1188_2;
    wire c1188;
    assign in1188_1 = {pp42[93]};
    assign in1188_2 = {pp43[92]};
    Full_Adder FA_1188(s1188, c1188, in1188_1, in1188_2, pp41[94]);
    wire[0:0] s1189, in1189_1, in1189_2;
    wire c1189;
    assign in1189_1 = {pp45[90]};
    assign in1189_2 = {pp46[89]};
    Full_Adder FA_1189(s1189, c1189, in1189_1, in1189_2, pp44[91]);
    wire[0:0] s1190, in1190_1, in1190_2;
    wire c1190;
    assign in1190_1 = {pp48[87]};
    assign in1190_2 = {pp49[86]};
    Full_Adder FA_1190(s1190, c1190, in1190_1, in1190_2, pp47[88]);
    wire[0:0] s1191, in1191_1, in1191_2;
    wire c1191;
    assign in1191_1 = {pp51[84]};
    assign in1191_2 = {pp52[83]};
    Full_Adder FA_1191(s1191, c1191, in1191_1, in1191_2, pp50[85]);
    wire[0:0] s1192, in1192_1, in1192_2;
    wire c1192;
    assign in1192_1 = {pp54[81]};
    assign in1192_2 = {pp55[80]};
    Full_Adder FA_1192(s1192, c1192, in1192_1, in1192_2, pp53[82]);
    wire[0:0] s1193, in1193_1, in1193_2;
    wire c1193;
    assign in1193_1 = {pp57[78]};
    assign in1193_2 = {pp58[77]};
    Full_Adder FA_1193(s1193, c1193, in1193_1, in1193_2, pp56[79]);
    wire[0:0] s1194, in1194_1, in1194_2;
    wire c1194;
    assign in1194_1 = {pp60[75]};
    assign in1194_2 = {pp61[74]};
    Full_Adder FA_1194(s1194, c1194, in1194_1, in1194_2, pp59[76]);
    wire[0:0] s1195, in1195_1, in1195_2;
    wire c1195;
    assign in1195_1 = {pp63[72]};
    assign in1195_2 = {pp64[71]};
    Full_Adder FA_1195(s1195, c1195, in1195_1, in1195_2, pp62[73]);
    wire[0:0] s1196, in1196_1, in1196_2;
    wire c1196;
    assign in1196_1 = {pp66[69]};
    assign in1196_2 = {pp67[68]};
    Full_Adder FA_1196(s1196, c1196, in1196_1, in1196_2, pp65[70]);
    wire[0:0] s1197, in1197_1, in1197_2;
    wire c1197;
    assign in1197_1 = {pp69[66]};
    assign in1197_2 = {pp70[65]};
    Full_Adder FA_1197(s1197, c1197, in1197_1, in1197_2, pp68[67]);
    wire[0:0] s1198, in1198_1, in1198_2;
    wire c1198;
    assign in1198_1 = {pp72[63]};
    assign in1198_2 = {pp73[62]};
    Full_Adder FA_1198(s1198, c1198, in1198_1, in1198_2, pp71[64]);
    wire[0:0] s1199, in1199_1, in1199_2;
    wire c1199;
    assign in1199_1 = {pp75[60]};
    assign in1199_2 = {pp76[59]};
    Full_Adder FA_1199(s1199, c1199, in1199_1, in1199_2, pp74[61]);
    wire[0:0] s1200, in1200_1, in1200_2;
    wire c1200;
    assign in1200_1 = {pp78[57]};
    assign in1200_2 = {pp79[56]};
    Full_Adder FA_1200(s1200, c1200, in1200_1, in1200_2, pp77[58]);
    wire[0:0] s1201, in1201_1, in1201_2;
    wire c1201;
    assign in1201_1 = {pp81[54]};
    assign in1201_2 = {pp82[53]};
    Full_Adder FA_1201(s1201, c1201, in1201_1, in1201_2, pp80[55]);
    wire[0:0] s1202, in1202_1, in1202_2;
    wire c1202;
    assign in1202_1 = {pp84[51]};
    assign in1202_2 = {pp85[50]};
    Full_Adder FA_1202(s1202, c1202, in1202_1, in1202_2, pp83[52]);
    wire[0:0] s1203, in1203_1, in1203_2;
    wire c1203;
    assign in1203_1 = {pp87[48]};
    assign in1203_2 = {pp88[47]};
    Full_Adder FA_1203(s1203, c1203, in1203_1, in1203_2, pp86[49]);
    wire[0:0] s1204, in1204_1, in1204_2;
    wire c1204;
    assign in1204_1 = {pp90[45]};
    assign in1204_2 = {pp91[44]};
    Full_Adder FA_1204(s1204, c1204, in1204_1, in1204_2, pp89[46]);
    wire[0:0] s1205, in1205_1, in1205_2;
    wire c1205;
    assign in1205_1 = {pp93[42]};
    assign in1205_2 = {pp94[41]};
    Full_Adder FA_1205(s1205, c1205, in1205_1, in1205_2, pp92[43]);
    wire[0:0] s1206, in1206_1, in1206_2;
    wire c1206;
    assign in1206_1 = {pp96[39]};
    assign in1206_2 = {pp97[38]};
    Full_Adder FA_1206(s1206, c1206, in1206_1, in1206_2, pp95[40]);
    wire[0:0] s1207, in1207_1, in1207_2;
    wire c1207;
    assign in1207_1 = {pp99[36]};
    assign in1207_2 = {pp100[35]};
    Full_Adder FA_1207(s1207, c1207, in1207_1, in1207_2, pp98[37]);
    wire[0:0] s1208, in1208_1, in1208_2;
    wire c1208;
    assign in1208_1 = {pp102[33]};
    assign in1208_2 = {pp103[32]};
    Full_Adder FA_1208(s1208, c1208, in1208_1, in1208_2, pp101[34]);
    wire[0:0] s1209, in1209_1, in1209_2;
    wire c1209;
    assign in1209_1 = {pp105[30]};
    assign in1209_2 = {pp106[29]};
    Full_Adder FA_1209(s1209, c1209, in1209_1, in1209_2, pp104[31]);
    wire[0:0] s1210, in1210_1, in1210_2;
    wire c1210;
    assign in1210_1 = {pp108[27]};
    assign in1210_2 = {pp109[26]};
    Full_Adder FA_1210(s1210, c1210, in1210_1, in1210_2, pp107[28]);
    wire[0:0] s1211, in1211_1, in1211_2;
    wire c1211;
    assign in1211_1 = {pp111[24]};
    assign in1211_2 = {pp112[23]};
    Full_Adder FA_1211(s1211, c1211, in1211_1, in1211_2, pp110[25]);
    wire[0:0] s1212, in1212_1, in1212_2;
    wire c1212;
    assign in1212_1 = {pp10[126]};
    assign in1212_2 = {pp11[125]};
    Full_Adder FA_1212(s1212, c1212, in1212_1, in1212_2, pp9[127]);
    wire[0:0] s1213, in1213_1, in1213_2;
    wire c1213;
    assign in1213_1 = {pp13[123]};
    assign in1213_2 = {pp14[122]};
    Full_Adder FA_1213(s1213, c1213, in1213_1, in1213_2, pp12[124]);
    wire[0:0] s1214, in1214_1, in1214_2;
    wire c1214;
    assign in1214_1 = {pp16[120]};
    assign in1214_2 = {pp17[119]};
    Full_Adder FA_1214(s1214, c1214, in1214_1, in1214_2, pp15[121]);
    wire[0:0] s1215, in1215_1, in1215_2;
    wire c1215;
    assign in1215_1 = {pp19[117]};
    assign in1215_2 = {pp20[116]};
    Full_Adder FA_1215(s1215, c1215, in1215_1, in1215_2, pp18[118]);
    wire[0:0] s1216, in1216_1, in1216_2;
    wire c1216;
    assign in1216_1 = {pp22[114]};
    assign in1216_2 = {pp23[113]};
    Full_Adder FA_1216(s1216, c1216, in1216_1, in1216_2, pp21[115]);
    wire[0:0] s1217, in1217_1, in1217_2;
    wire c1217;
    assign in1217_1 = {pp25[111]};
    assign in1217_2 = {pp26[110]};
    Full_Adder FA_1217(s1217, c1217, in1217_1, in1217_2, pp24[112]);
    wire[0:0] s1218, in1218_1, in1218_2;
    wire c1218;
    assign in1218_1 = {pp28[108]};
    assign in1218_2 = {pp29[107]};
    Full_Adder FA_1218(s1218, c1218, in1218_1, in1218_2, pp27[109]);
    wire[0:0] s1219, in1219_1, in1219_2;
    wire c1219;
    assign in1219_1 = {pp31[105]};
    assign in1219_2 = {pp32[104]};
    Full_Adder FA_1219(s1219, c1219, in1219_1, in1219_2, pp30[106]);
    wire[0:0] s1220, in1220_1, in1220_2;
    wire c1220;
    assign in1220_1 = {pp34[102]};
    assign in1220_2 = {pp35[101]};
    Full_Adder FA_1220(s1220, c1220, in1220_1, in1220_2, pp33[103]);
    wire[0:0] s1221, in1221_1, in1221_2;
    wire c1221;
    assign in1221_1 = {pp37[99]};
    assign in1221_2 = {pp38[98]};
    Full_Adder FA_1221(s1221, c1221, in1221_1, in1221_2, pp36[100]);
    wire[0:0] s1222, in1222_1, in1222_2;
    wire c1222;
    assign in1222_1 = {pp40[96]};
    assign in1222_2 = {pp41[95]};
    Full_Adder FA_1222(s1222, c1222, in1222_1, in1222_2, pp39[97]);
    wire[0:0] s1223, in1223_1, in1223_2;
    wire c1223;
    assign in1223_1 = {pp43[93]};
    assign in1223_2 = {pp44[92]};
    Full_Adder FA_1223(s1223, c1223, in1223_1, in1223_2, pp42[94]);
    wire[0:0] s1224, in1224_1, in1224_2;
    wire c1224;
    assign in1224_1 = {pp46[90]};
    assign in1224_2 = {pp47[89]};
    Full_Adder FA_1224(s1224, c1224, in1224_1, in1224_2, pp45[91]);
    wire[0:0] s1225, in1225_1, in1225_2;
    wire c1225;
    assign in1225_1 = {pp49[87]};
    assign in1225_2 = {pp50[86]};
    Full_Adder FA_1225(s1225, c1225, in1225_1, in1225_2, pp48[88]);
    wire[0:0] s1226, in1226_1, in1226_2;
    wire c1226;
    assign in1226_1 = {pp52[84]};
    assign in1226_2 = {pp53[83]};
    Full_Adder FA_1226(s1226, c1226, in1226_1, in1226_2, pp51[85]);
    wire[0:0] s1227, in1227_1, in1227_2;
    wire c1227;
    assign in1227_1 = {pp55[81]};
    assign in1227_2 = {pp56[80]};
    Full_Adder FA_1227(s1227, c1227, in1227_1, in1227_2, pp54[82]);
    wire[0:0] s1228, in1228_1, in1228_2;
    wire c1228;
    assign in1228_1 = {pp58[78]};
    assign in1228_2 = {pp59[77]};
    Full_Adder FA_1228(s1228, c1228, in1228_1, in1228_2, pp57[79]);
    wire[0:0] s1229, in1229_1, in1229_2;
    wire c1229;
    assign in1229_1 = {pp61[75]};
    assign in1229_2 = {pp62[74]};
    Full_Adder FA_1229(s1229, c1229, in1229_1, in1229_2, pp60[76]);
    wire[0:0] s1230, in1230_1, in1230_2;
    wire c1230;
    assign in1230_1 = {pp64[72]};
    assign in1230_2 = {pp65[71]};
    Full_Adder FA_1230(s1230, c1230, in1230_1, in1230_2, pp63[73]);
    wire[0:0] s1231, in1231_1, in1231_2;
    wire c1231;
    assign in1231_1 = {pp67[69]};
    assign in1231_2 = {pp68[68]};
    Full_Adder FA_1231(s1231, c1231, in1231_1, in1231_2, pp66[70]);
    wire[0:0] s1232, in1232_1, in1232_2;
    wire c1232;
    assign in1232_1 = {pp70[66]};
    assign in1232_2 = {pp71[65]};
    Full_Adder FA_1232(s1232, c1232, in1232_1, in1232_2, pp69[67]);
    wire[0:0] s1233, in1233_1, in1233_2;
    wire c1233;
    assign in1233_1 = {pp73[63]};
    assign in1233_2 = {pp74[62]};
    Full_Adder FA_1233(s1233, c1233, in1233_1, in1233_2, pp72[64]);
    wire[0:0] s1234, in1234_1, in1234_2;
    wire c1234;
    assign in1234_1 = {pp76[60]};
    assign in1234_2 = {pp77[59]};
    Full_Adder FA_1234(s1234, c1234, in1234_1, in1234_2, pp75[61]);
    wire[0:0] s1235, in1235_1, in1235_2;
    wire c1235;
    assign in1235_1 = {pp79[57]};
    assign in1235_2 = {pp80[56]};
    Full_Adder FA_1235(s1235, c1235, in1235_1, in1235_2, pp78[58]);
    wire[0:0] s1236, in1236_1, in1236_2;
    wire c1236;
    assign in1236_1 = {pp82[54]};
    assign in1236_2 = {pp83[53]};
    Full_Adder FA_1236(s1236, c1236, in1236_1, in1236_2, pp81[55]);
    wire[0:0] s1237, in1237_1, in1237_2;
    wire c1237;
    assign in1237_1 = {pp85[51]};
    assign in1237_2 = {pp86[50]};
    Full_Adder FA_1237(s1237, c1237, in1237_1, in1237_2, pp84[52]);
    wire[0:0] s1238, in1238_1, in1238_2;
    wire c1238;
    assign in1238_1 = {pp88[48]};
    assign in1238_2 = {pp89[47]};
    Full_Adder FA_1238(s1238, c1238, in1238_1, in1238_2, pp87[49]);
    wire[0:0] s1239, in1239_1, in1239_2;
    wire c1239;
    assign in1239_1 = {pp91[45]};
    assign in1239_2 = {pp92[44]};
    Full_Adder FA_1239(s1239, c1239, in1239_1, in1239_2, pp90[46]);
    wire[0:0] s1240, in1240_1, in1240_2;
    wire c1240;
    assign in1240_1 = {pp94[42]};
    assign in1240_2 = {pp95[41]};
    Full_Adder FA_1240(s1240, c1240, in1240_1, in1240_2, pp93[43]);
    wire[0:0] s1241, in1241_1, in1241_2;
    wire c1241;
    assign in1241_1 = {pp97[39]};
    assign in1241_2 = {pp98[38]};
    Full_Adder FA_1241(s1241, c1241, in1241_1, in1241_2, pp96[40]);
    wire[0:0] s1242, in1242_1, in1242_2;
    wire c1242;
    assign in1242_1 = {pp100[36]};
    assign in1242_2 = {pp101[35]};
    Full_Adder FA_1242(s1242, c1242, in1242_1, in1242_2, pp99[37]);
    wire[0:0] s1243, in1243_1, in1243_2;
    wire c1243;
    assign in1243_1 = {pp103[33]};
    assign in1243_2 = {pp104[32]};
    Full_Adder FA_1243(s1243, c1243, in1243_1, in1243_2, pp102[34]);
    wire[0:0] s1244, in1244_1, in1244_2;
    wire c1244;
    assign in1244_1 = {pp106[30]};
    assign in1244_2 = {pp107[29]};
    Full_Adder FA_1244(s1244, c1244, in1244_1, in1244_2, pp105[31]);
    wire[0:0] s1245, in1245_1, in1245_2;
    wire c1245;
    assign in1245_1 = {pp109[27]};
    assign in1245_2 = {pp110[26]};
    Full_Adder FA_1245(s1245, c1245, in1245_1, in1245_2, pp108[28]);
    wire[0:0] s1246, in1246_1, in1246_2;
    wire c1246;
    assign in1246_1 = {pp11[126]};
    assign in1246_2 = {pp12[125]};
    Full_Adder FA_1246(s1246, c1246, in1246_1, in1246_2, pp10[127]);
    wire[0:0] s1247, in1247_1, in1247_2;
    wire c1247;
    assign in1247_1 = {pp14[123]};
    assign in1247_2 = {pp15[122]};
    Full_Adder FA_1247(s1247, c1247, in1247_1, in1247_2, pp13[124]);
    wire[0:0] s1248, in1248_1, in1248_2;
    wire c1248;
    assign in1248_1 = {pp17[120]};
    assign in1248_2 = {pp18[119]};
    Full_Adder FA_1248(s1248, c1248, in1248_1, in1248_2, pp16[121]);
    wire[0:0] s1249, in1249_1, in1249_2;
    wire c1249;
    assign in1249_1 = {pp20[117]};
    assign in1249_2 = {pp21[116]};
    Full_Adder FA_1249(s1249, c1249, in1249_1, in1249_2, pp19[118]);
    wire[0:0] s1250, in1250_1, in1250_2;
    wire c1250;
    assign in1250_1 = {pp23[114]};
    assign in1250_2 = {pp24[113]};
    Full_Adder FA_1250(s1250, c1250, in1250_1, in1250_2, pp22[115]);
    wire[0:0] s1251, in1251_1, in1251_2;
    wire c1251;
    assign in1251_1 = {pp26[111]};
    assign in1251_2 = {pp27[110]};
    Full_Adder FA_1251(s1251, c1251, in1251_1, in1251_2, pp25[112]);
    wire[0:0] s1252, in1252_1, in1252_2;
    wire c1252;
    assign in1252_1 = {pp29[108]};
    assign in1252_2 = {pp30[107]};
    Full_Adder FA_1252(s1252, c1252, in1252_1, in1252_2, pp28[109]);
    wire[0:0] s1253, in1253_1, in1253_2;
    wire c1253;
    assign in1253_1 = {pp32[105]};
    assign in1253_2 = {pp33[104]};
    Full_Adder FA_1253(s1253, c1253, in1253_1, in1253_2, pp31[106]);
    wire[0:0] s1254, in1254_1, in1254_2;
    wire c1254;
    assign in1254_1 = {pp35[102]};
    assign in1254_2 = {pp36[101]};
    Full_Adder FA_1254(s1254, c1254, in1254_1, in1254_2, pp34[103]);
    wire[0:0] s1255, in1255_1, in1255_2;
    wire c1255;
    assign in1255_1 = {pp38[99]};
    assign in1255_2 = {pp39[98]};
    Full_Adder FA_1255(s1255, c1255, in1255_1, in1255_2, pp37[100]);
    wire[0:0] s1256, in1256_1, in1256_2;
    wire c1256;
    assign in1256_1 = {pp41[96]};
    assign in1256_2 = {pp42[95]};
    Full_Adder FA_1256(s1256, c1256, in1256_1, in1256_2, pp40[97]);
    wire[0:0] s1257, in1257_1, in1257_2;
    wire c1257;
    assign in1257_1 = {pp44[93]};
    assign in1257_2 = {pp45[92]};
    Full_Adder FA_1257(s1257, c1257, in1257_1, in1257_2, pp43[94]);
    wire[0:0] s1258, in1258_1, in1258_2;
    wire c1258;
    assign in1258_1 = {pp47[90]};
    assign in1258_2 = {pp48[89]};
    Full_Adder FA_1258(s1258, c1258, in1258_1, in1258_2, pp46[91]);
    wire[0:0] s1259, in1259_1, in1259_2;
    wire c1259;
    assign in1259_1 = {pp50[87]};
    assign in1259_2 = {pp51[86]};
    Full_Adder FA_1259(s1259, c1259, in1259_1, in1259_2, pp49[88]);
    wire[0:0] s1260, in1260_1, in1260_2;
    wire c1260;
    assign in1260_1 = {pp53[84]};
    assign in1260_2 = {pp54[83]};
    Full_Adder FA_1260(s1260, c1260, in1260_1, in1260_2, pp52[85]);
    wire[0:0] s1261, in1261_1, in1261_2;
    wire c1261;
    assign in1261_1 = {pp56[81]};
    assign in1261_2 = {pp57[80]};
    Full_Adder FA_1261(s1261, c1261, in1261_1, in1261_2, pp55[82]);
    wire[0:0] s1262, in1262_1, in1262_2;
    wire c1262;
    assign in1262_1 = {pp59[78]};
    assign in1262_2 = {pp60[77]};
    Full_Adder FA_1262(s1262, c1262, in1262_1, in1262_2, pp58[79]);
    wire[0:0] s1263, in1263_1, in1263_2;
    wire c1263;
    assign in1263_1 = {pp62[75]};
    assign in1263_2 = {pp63[74]};
    Full_Adder FA_1263(s1263, c1263, in1263_1, in1263_2, pp61[76]);
    wire[0:0] s1264, in1264_1, in1264_2;
    wire c1264;
    assign in1264_1 = {pp65[72]};
    assign in1264_2 = {pp66[71]};
    Full_Adder FA_1264(s1264, c1264, in1264_1, in1264_2, pp64[73]);
    wire[0:0] s1265, in1265_1, in1265_2;
    wire c1265;
    assign in1265_1 = {pp68[69]};
    assign in1265_2 = {pp69[68]};
    Full_Adder FA_1265(s1265, c1265, in1265_1, in1265_2, pp67[70]);
    wire[0:0] s1266, in1266_1, in1266_2;
    wire c1266;
    assign in1266_1 = {pp71[66]};
    assign in1266_2 = {pp72[65]};
    Full_Adder FA_1266(s1266, c1266, in1266_1, in1266_2, pp70[67]);
    wire[0:0] s1267, in1267_1, in1267_2;
    wire c1267;
    assign in1267_1 = {pp74[63]};
    assign in1267_2 = {pp75[62]};
    Full_Adder FA_1267(s1267, c1267, in1267_1, in1267_2, pp73[64]);
    wire[0:0] s1268, in1268_1, in1268_2;
    wire c1268;
    assign in1268_1 = {pp77[60]};
    assign in1268_2 = {pp78[59]};
    Full_Adder FA_1268(s1268, c1268, in1268_1, in1268_2, pp76[61]);
    wire[0:0] s1269, in1269_1, in1269_2;
    wire c1269;
    assign in1269_1 = {pp80[57]};
    assign in1269_2 = {pp81[56]};
    Full_Adder FA_1269(s1269, c1269, in1269_1, in1269_2, pp79[58]);
    wire[0:0] s1270, in1270_1, in1270_2;
    wire c1270;
    assign in1270_1 = {pp83[54]};
    assign in1270_2 = {pp84[53]};
    Full_Adder FA_1270(s1270, c1270, in1270_1, in1270_2, pp82[55]);
    wire[0:0] s1271, in1271_1, in1271_2;
    wire c1271;
    assign in1271_1 = {pp86[51]};
    assign in1271_2 = {pp87[50]};
    Full_Adder FA_1271(s1271, c1271, in1271_1, in1271_2, pp85[52]);
    wire[0:0] s1272, in1272_1, in1272_2;
    wire c1272;
    assign in1272_1 = {pp89[48]};
    assign in1272_2 = {pp90[47]};
    Full_Adder FA_1272(s1272, c1272, in1272_1, in1272_2, pp88[49]);
    wire[0:0] s1273, in1273_1, in1273_2;
    wire c1273;
    assign in1273_1 = {pp92[45]};
    assign in1273_2 = {pp93[44]};
    Full_Adder FA_1273(s1273, c1273, in1273_1, in1273_2, pp91[46]);
    wire[0:0] s1274, in1274_1, in1274_2;
    wire c1274;
    assign in1274_1 = {pp95[42]};
    assign in1274_2 = {pp96[41]};
    Full_Adder FA_1274(s1274, c1274, in1274_1, in1274_2, pp94[43]);
    wire[0:0] s1275, in1275_1, in1275_2;
    wire c1275;
    assign in1275_1 = {pp98[39]};
    assign in1275_2 = {pp99[38]};
    Full_Adder FA_1275(s1275, c1275, in1275_1, in1275_2, pp97[40]);
    wire[0:0] s1276, in1276_1, in1276_2;
    wire c1276;
    assign in1276_1 = {pp101[36]};
    assign in1276_2 = {pp102[35]};
    Full_Adder FA_1276(s1276, c1276, in1276_1, in1276_2, pp100[37]);
    wire[0:0] s1277, in1277_1, in1277_2;
    wire c1277;
    assign in1277_1 = {pp104[33]};
    assign in1277_2 = {pp105[32]};
    Full_Adder FA_1277(s1277, c1277, in1277_1, in1277_2, pp103[34]);
    wire[0:0] s1278, in1278_1, in1278_2;
    wire c1278;
    assign in1278_1 = {pp107[30]};
    assign in1278_2 = {pp108[29]};
    Full_Adder FA_1278(s1278, c1278, in1278_1, in1278_2, pp106[31]);
    wire[0:0] s1279, in1279_1, in1279_2;
    wire c1279;
    assign in1279_1 = {pp12[126]};
    assign in1279_2 = {pp13[125]};
    Full_Adder FA_1279(s1279, c1279, in1279_1, in1279_2, pp11[127]);
    wire[0:0] s1280, in1280_1, in1280_2;
    wire c1280;
    assign in1280_1 = {pp15[123]};
    assign in1280_2 = {pp16[122]};
    Full_Adder FA_1280(s1280, c1280, in1280_1, in1280_2, pp14[124]);
    wire[0:0] s1281, in1281_1, in1281_2;
    wire c1281;
    assign in1281_1 = {pp18[120]};
    assign in1281_2 = {pp19[119]};
    Full_Adder FA_1281(s1281, c1281, in1281_1, in1281_2, pp17[121]);
    wire[0:0] s1282, in1282_1, in1282_2;
    wire c1282;
    assign in1282_1 = {pp21[117]};
    assign in1282_2 = {pp22[116]};
    Full_Adder FA_1282(s1282, c1282, in1282_1, in1282_2, pp20[118]);
    wire[0:0] s1283, in1283_1, in1283_2;
    wire c1283;
    assign in1283_1 = {pp24[114]};
    assign in1283_2 = {pp25[113]};
    Full_Adder FA_1283(s1283, c1283, in1283_1, in1283_2, pp23[115]);
    wire[0:0] s1284, in1284_1, in1284_2;
    wire c1284;
    assign in1284_1 = {pp27[111]};
    assign in1284_2 = {pp28[110]};
    Full_Adder FA_1284(s1284, c1284, in1284_1, in1284_2, pp26[112]);
    wire[0:0] s1285, in1285_1, in1285_2;
    wire c1285;
    assign in1285_1 = {pp30[108]};
    assign in1285_2 = {pp31[107]};
    Full_Adder FA_1285(s1285, c1285, in1285_1, in1285_2, pp29[109]);
    wire[0:0] s1286, in1286_1, in1286_2;
    wire c1286;
    assign in1286_1 = {pp33[105]};
    assign in1286_2 = {pp34[104]};
    Full_Adder FA_1286(s1286, c1286, in1286_1, in1286_2, pp32[106]);
    wire[0:0] s1287, in1287_1, in1287_2;
    wire c1287;
    assign in1287_1 = {pp36[102]};
    assign in1287_2 = {pp37[101]};
    Full_Adder FA_1287(s1287, c1287, in1287_1, in1287_2, pp35[103]);
    wire[0:0] s1288, in1288_1, in1288_2;
    wire c1288;
    assign in1288_1 = {pp39[99]};
    assign in1288_2 = {pp40[98]};
    Full_Adder FA_1288(s1288, c1288, in1288_1, in1288_2, pp38[100]);
    wire[0:0] s1289, in1289_1, in1289_2;
    wire c1289;
    assign in1289_1 = {pp42[96]};
    assign in1289_2 = {pp43[95]};
    Full_Adder FA_1289(s1289, c1289, in1289_1, in1289_2, pp41[97]);
    wire[0:0] s1290, in1290_1, in1290_2;
    wire c1290;
    assign in1290_1 = {pp45[93]};
    assign in1290_2 = {pp46[92]};
    Full_Adder FA_1290(s1290, c1290, in1290_1, in1290_2, pp44[94]);
    wire[0:0] s1291, in1291_1, in1291_2;
    wire c1291;
    assign in1291_1 = {pp48[90]};
    assign in1291_2 = {pp49[89]};
    Full_Adder FA_1291(s1291, c1291, in1291_1, in1291_2, pp47[91]);
    wire[0:0] s1292, in1292_1, in1292_2;
    wire c1292;
    assign in1292_1 = {pp51[87]};
    assign in1292_2 = {pp52[86]};
    Full_Adder FA_1292(s1292, c1292, in1292_1, in1292_2, pp50[88]);
    wire[0:0] s1293, in1293_1, in1293_2;
    wire c1293;
    assign in1293_1 = {pp54[84]};
    assign in1293_2 = {pp55[83]};
    Full_Adder FA_1293(s1293, c1293, in1293_1, in1293_2, pp53[85]);
    wire[0:0] s1294, in1294_1, in1294_2;
    wire c1294;
    assign in1294_1 = {pp57[81]};
    assign in1294_2 = {pp58[80]};
    Full_Adder FA_1294(s1294, c1294, in1294_1, in1294_2, pp56[82]);
    wire[0:0] s1295, in1295_1, in1295_2;
    wire c1295;
    assign in1295_1 = {pp60[78]};
    assign in1295_2 = {pp61[77]};
    Full_Adder FA_1295(s1295, c1295, in1295_1, in1295_2, pp59[79]);
    wire[0:0] s1296, in1296_1, in1296_2;
    wire c1296;
    assign in1296_1 = {pp63[75]};
    assign in1296_2 = {pp64[74]};
    Full_Adder FA_1296(s1296, c1296, in1296_1, in1296_2, pp62[76]);
    wire[0:0] s1297, in1297_1, in1297_2;
    wire c1297;
    assign in1297_1 = {pp66[72]};
    assign in1297_2 = {pp67[71]};
    Full_Adder FA_1297(s1297, c1297, in1297_1, in1297_2, pp65[73]);
    wire[0:0] s1298, in1298_1, in1298_2;
    wire c1298;
    assign in1298_1 = {pp69[69]};
    assign in1298_2 = {pp70[68]};
    Full_Adder FA_1298(s1298, c1298, in1298_1, in1298_2, pp68[70]);
    wire[0:0] s1299, in1299_1, in1299_2;
    wire c1299;
    assign in1299_1 = {pp72[66]};
    assign in1299_2 = {pp73[65]};
    Full_Adder FA_1299(s1299, c1299, in1299_1, in1299_2, pp71[67]);
    wire[0:0] s1300, in1300_1, in1300_2;
    wire c1300;
    assign in1300_1 = {pp75[63]};
    assign in1300_2 = {pp76[62]};
    Full_Adder FA_1300(s1300, c1300, in1300_1, in1300_2, pp74[64]);
    wire[0:0] s1301, in1301_1, in1301_2;
    wire c1301;
    assign in1301_1 = {pp78[60]};
    assign in1301_2 = {pp79[59]};
    Full_Adder FA_1301(s1301, c1301, in1301_1, in1301_2, pp77[61]);
    wire[0:0] s1302, in1302_1, in1302_2;
    wire c1302;
    assign in1302_1 = {pp81[57]};
    assign in1302_2 = {pp82[56]};
    Full_Adder FA_1302(s1302, c1302, in1302_1, in1302_2, pp80[58]);
    wire[0:0] s1303, in1303_1, in1303_2;
    wire c1303;
    assign in1303_1 = {pp84[54]};
    assign in1303_2 = {pp85[53]};
    Full_Adder FA_1303(s1303, c1303, in1303_1, in1303_2, pp83[55]);
    wire[0:0] s1304, in1304_1, in1304_2;
    wire c1304;
    assign in1304_1 = {pp87[51]};
    assign in1304_2 = {pp88[50]};
    Full_Adder FA_1304(s1304, c1304, in1304_1, in1304_2, pp86[52]);
    wire[0:0] s1305, in1305_1, in1305_2;
    wire c1305;
    assign in1305_1 = {pp90[48]};
    assign in1305_2 = {pp91[47]};
    Full_Adder FA_1305(s1305, c1305, in1305_1, in1305_2, pp89[49]);
    wire[0:0] s1306, in1306_1, in1306_2;
    wire c1306;
    assign in1306_1 = {pp93[45]};
    assign in1306_2 = {pp94[44]};
    Full_Adder FA_1306(s1306, c1306, in1306_1, in1306_2, pp92[46]);
    wire[0:0] s1307, in1307_1, in1307_2;
    wire c1307;
    assign in1307_1 = {pp96[42]};
    assign in1307_2 = {pp97[41]};
    Full_Adder FA_1307(s1307, c1307, in1307_1, in1307_2, pp95[43]);
    wire[0:0] s1308, in1308_1, in1308_2;
    wire c1308;
    assign in1308_1 = {pp99[39]};
    assign in1308_2 = {pp100[38]};
    Full_Adder FA_1308(s1308, c1308, in1308_1, in1308_2, pp98[40]);
    wire[0:0] s1309, in1309_1, in1309_2;
    wire c1309;
    assign in1309_1 = {pp102[36]};
    assign in1309_2 = {pp103[35]};
    Full_Adder FA_1309(s1309, c1309, in1309_1, in1309_2, pp101[37]);
    wire[0:0] s1310, in1310_1, in1310_2;
    wire c1310;
    assign in1310_1 = {pp105[33]};
    assign in1310_2 = {pp106[32]};
    Full_Adder FA_1310(s1310, c1310, in1310_1, in1310_2, pp104[34]);
    wire[0:0] s1311, in1311_1, in1311_2;
    wire c1311;
    assign in1311_1 = {pp13[126]};
    assign in1311_2 = {pp14[125]};
    Full_Adder FA_1311(s1311, c1311, in1311_1, in1311_2, pp12[127]);
    wire[0:0] s1312, in1312_1, in1312_2;
    wire c1312;
    assign in1312_1 = {pp16[123]};
    assign in1312_2 = {pp17[122]};
    Full_Adder FA_1312(s1312, c1312, in1312_1, in1312_2, pp15[124]);
    wire[0:0] s1313, in1313_1, in1313_2;
    wire c1313;
    assign in1313_1 = {pp19[120]};
    assign in1313_2 = {pp20[119]};
    Full_Adder FA_1313(s1313, c1313, in1313_1, in1313_2, pp18[121]);
    wire[0:0] s1314, in1314_1, in1314_2;
    wire c1314;
    assign in1314_1 = {pp22[117]};
    assign in1314_2 = {pp23[116]};
    Full_Adder FA_1314(s1314, c1314, in1314_1, in1314_2, pp21[118]);
    wire[0:0] s1315, in1315_1, in1315_2;
    wire c1315;
    assign in1315_1 = {pp25[114]};
    assign in1315_2 = {pp26[113]};
    Full_Adder FA_1315(s1315, c1315, in1315_1, in1315_2, pp24[115]);
    wire[0:0] s1316, in1316_1, in1316_2;
    wire c1316;
    assign in1316_1 = {pp28[111]};
    assign in1316_2 = {pp29[110]};
    Full_Adder FA_1316(s1316, c1316, in1316_1, in1316_2, pp27[112]);
    wire[0:0] s1317, in1317_1, in1317_2;
    wire c1317;
    assign in1317_1 = {pp31[108]};
    assign in1317_2 = {pp32[107]};
    Full_Adder FA_1317(s1317, c1317, in1317_1, in1317_2, pp30[109]);
    wire[0:0] s1318, in1318_1, in1318_2;
    wire c1318;
    assign in1318_1 = {pp34[105]};
    assign in1318_2 = {pp35[104]};
    Full_Adder FA_1318(s1318, c1318, in1318_1, in1318_2, pp33[106]);
    wire[0:0] s1319, in1319_1, in1319_2;
    wire c1319;
    assign in1319_1 = {pp37[102]};
    assign in1319_2 = {pp38[101]};
    Full_Adder FA_1319(s1319, c1319, in1319_1, in1319_2, pp36[103]);
    wire[0:0] s1320, in1320_1, in1320_2;
    wire c1320;
    assign in1320_1 = {pp40[99]};
    assign in1320_2 = {pp41[98]};
    Full_Adder FA_1320(s1320, c1320, in1320_1, in1320_2, pp39[100]);
    wire[0:0] s1321, in1321_1, in1321_2;
    wire c1321;
    assign in1321_1 = {pp43[96]};
    assign in1321_2 = {pp44[95]};
    Full_Adder FA_1321(s1321, c1321, in1321_1, in1321_2, pp42[97]);
    wire[0:0] s1322, in1322_1, in1322_2;
    wire c1322;
    assign in1322_1 = {pp46[93]};
    assign in1322_2 = {pp47[92]};
    Full_Adder FA_1322(s1322, c1322, in1322_1, in1322_2, pp45[94]);
    wire[0:0] s1323, in1323_1, in1323_2;
    wire c1323;
    assign in1323_1 = {pp49[90]};
    assign in1323_2 = {pp50[89]};
    Full_Adder FA_1323(s1323, c1323, in1323_1, in1323_2, pp48[91]);
    wire[0:0] s1324, in1324_1, in1324_2;
    wire c1324;
    assign in1324_1 = {pp52[87]};
    assign in1324_2 = {pp53[86]};
    Full_Adder FA_1324(s1324, c1324, in1324_1, in1324_2, pp51[88]);
    wire[0:0] s1325, in1325_1, in1325_2;
    wire c1325;
    assign in1325_1 = {pp55[84]};
    assign in1325_2 = {pp56[83]};
    Full_Adder FA_1325(s1325, c1325, in1325_1, in1325_2, pp54[85]);
    wire[0:0] s1326, in1326_1, in1326_2;
    wire c1326;
    assign in1326_1 = {pp58[81]};
    assign in1326_2 = {pp59[80]};
    Full_Adder FA_1326(s1326, c1326, in1326_1, in1326_2, pp57[82]);
    wire[0:0] s1327, in1327_1, in1327_2;
    wire c1327;
    assign in1327_1 = {pp61[78]};
    assign in1327_2 = {pp62[77]};
    Full_Adder FA_1327(s1327, c1327, in1327_1, in1327_2, pp60[79]);
    wire[0:0] s1328, in1328_1, in1328_2;
    wire c1328;
    assign in1328_1 = {pp64[75]};
    assign in1328_2 = {pp65[74]};
    Full_Adder FA_1328(s1328, c1328, in1328_1, in1328_2, pp63[76]);
    wire[0:0] s1329, in1329_1, in1329_2;
    wire c1329;
    assign in1329_1 = {pp67[72]};
    assign in1329_2 = {pp68[71]};
    Full_Adder FA_1329(s1329, c1329, in1329_1, in1329_2, pp66[73]);
    wire[0:0] s1330, in1330_1, in1330_2;
    wire c1330;
    assign in1330_1 = {pp70[69]};
    assign in1330_2 = {pp71[68]};
    Full_Adder FA_1330(s1330, c1330, in1330_1, in1330_2, pp69[70]);
    wire[0:0] s1331, in1331_1, in1331_2;
    wire c1331;
    assign in1331_1 = {pp73[66]};
    assign in1331_2 = {pp74[65]};
    Full_Adder FA_1331(s1331, c1331, in1331_1, in1331_2, pp72[67]);
    wire[0:0] s1332, in1332_1, in1332_2;
    wire c1332;
    assign in1332_1 = {pp76[63]};
    assign in1332_2 = {pp77[62]};
    Full_Adder FA_1332(s1332, c1332, in1332_1, in1332_2, pp75[64]);
    wire[0:0] s1333, in1333_1, in1333_2;
    wire c1333;
    assign in1333_1 = {pp79[60]};
    assign in1333_2 = {pp80[59]};
    Full_Adder FA_1333(s1333, c1333, in1333_1, in1333_2, pp78[61]);
    wire[0:0] s1334, in1334_1, in1334_2;
    wire c1334;
    assign in1334_1 = {pp82[57]};
    assign in1334_2 = {pp83[56]};
    Full_Adder FA_1334(s1334, c1334, in1334_1, in1334_2, pp81[58]);
    wire[0:0] s1335, in1335_1, in1335_2;
    wire c1335;
    assign in1335_1 = {pp85[54]};
    assign in1335_2 = {pp86[53]};
    Full_Adder FA_1335(s1335, c1335, in1335_1, in1335_2, pp84[55]);
    wire[0:0] s1336, in1336_1, in1336_2;
    wire c1336;
    assign in1336_1 = {pp88[51]};
    assign in1336_2 = {pp89[50]};
    Full_Adder FA_1336(s1336, c1336, in1336_1, in1336_2, pp87[52]);
    wire[0:0] s1337, in1337_1, in1337_2;
    wire c1337;
    assign in1337_1 = {pp91[48]};
    assign in1337_2 = {pp92[47]};
    Full_Adder FA_1337(s1337, c1337, in1337_1, in1337_2, pp90[49]);
    wire[0:0] s1338, in1338_1, in1338_2;
    wire c1338;
    assign in1338_1 = {pp94[45]};
    assign in1338_2 = {pp95[44]};
    Full_Adder FA_1338(s1338, c1338, in1338_1, in1338_2, pp93[46]);
    wire[0:0] s1339, in1339_1, in1339_2;
    wire c1339;
    assign in1339_1 = {pp97[42]};
    assign in1339_2 = {pp98[41]};
    Full_Adder FA_1339(s1339, c1339, in1339_1, in1339_2, pp96[43]);
    wire[0:0] s1340, in1340_1, in1340_2;
    wire c1340;
    assign in1340_1 = {pp100[39]};
    assign in1340_2 = {pp101[38]};
    Full_Adder FA_1340(s1340, c1340, in1340_1, in1340_2, pp99[40]);
    wire[0:0] s1341, in1341_1, in1341_2;
    wire c1341;
    assign in1341_1 = {pp103[36]};
    assign in1341_2 = {pp104[35]};
    Full_Adder FA_1341(s1341, c1341, in1341_1, in1341_2, pp102[37]);
    wire[0:0] s1342, in1342_1, in1342_2;
    wire c1342;
    assign in1342_1 = {pp14[126]};
    assign in1342_2 = {pp15[125]};
    Full_Adder FA_1342(s1342, c1342, in1342_1, in1342_2, pp13[127]);
    wire[0:0] s1343, in1343_1, in1343_2;
    wire c1343;
    assign in1343_1 = {pp17[123]};
    assign in1343_2 = {pp18[122]};
    Full_Adder FA_1343(s1343, c1343, in1343_1, in1343_2, pp16[124]);
    wire[0:0] s1344, in1344_1, in1344_2;
    wire c1344;
    assign in1344_1 = {pp20[120]};
    assign in1344_2 = {pp21[119]};
    Full_Adder FA_1344(s1344, c1344, in1344_1, in1344_2, pp19[121]);
    wire[0:0] s1345, in1345_1, in1345_2;
    wire c1345;
    assign in1345_1 = {pp23[117]};
    assign in1345_2 = {pp24[116]};
    Full_Adder FA_1345(s1345, c1345, in1345_1, in1345_2, pp22[118]);
    wire[0:0] s1346, in1346_1, in1346_2;
    wire c1346;
    assign in1346_1 = {pp26[114]};
    assign in1346_2 = {pp27[113]};
    Full_Adder FA_1346(s1346, c1346, in1346_1, in1346_2, pp25[115]);
    wire[0:0] s1347, in1347_1, in1347_2;
    wire c1347;
    assign in1347_1 = {pp29[111]};
    assign in1347_2 = {pp30[110]};
    Full_Adder FA_1347(s1347, c1347, in1347_1, in1347_2, pp28[112]);
    wire[0:0] s1348, in1348_1, in1348_2;
    wire c1348;
    assign in1348_1 = {pp32[108]};
    assign in1348_2 = {pp33[107]};
    Full_Adder FA_1348(s1348, c1348, in1348_1, in1348_2, pp31[109]);
    wire[0:0] s1349, in1349_1, in1349_2;
    wire c1349;
    assign in1349_1 = {pp35[105]};
    assign in1349_2 = {pp36[104]};
    Full_Adder FA_1349(s1349, c1349, in1349_1, in1349_2, pp34[106]);
    wire[0:0] s1350, in1350_1, in1350_2;
    wire c1350;
    assign in1350_1 = {pp38[102]};
    assign in1350_2 = {pp39[101]};
    Full_Adder FA_1350(s1350, c1350, in1350_1, in1350_2, pp37[103]);
    wire[0:0] s1351, in1351_1, in1351_2;
    wire c1351;
    assign in1351_1 = {pp41[99]};
    assign in1351_2 = {pp42[98]};
    Full_Adder FA_1351(s1351, c1351, in1351_1, in1351_2, pp40[100]);
    wire[0:0] s1352, in1352_1, in1352_2;
    wire c1352;
    assign in1352_1 = {pp44[96]};
    assign in1352_2 = {pp45[95]};
    Full_Adder FA_1352(s1352, c1352, in1352_1, in1352_2, pp43[97]);
    wire[0:0] s1353, in1353_1, in1353_2;
    wire c1353;
    assign in1353_1 = {pp47[93]};
    assign in1353_2 = {pp48[92]};
    Full_Adder FA_1353(s1353, c1353, in1353_1, in1353_2, pp46[94]);
    wire[0:0] s1354, in1354_1, in1354_2;
    wire c1354;
    assign in1354_1 = {pp50[90]};
    assign in1354_2 = {pp51[89]};
    Full_Adder FA_1354(s1354, c1354, in1354_1, in1354_2, pp49[91]);
    wire[0:0] s1355, in1355_1, in1355_2;
    wire c1355;
    assign in1355_1 = {pp53[87]};
    assign in1355_2 = {pp54[86]};
    Full_Adder FA_1355(s1355, c1355, in1355_1, in1355_2, pp52[88]);
    wire[0:0] s1356, in1356_1, in1356_2;
    wire c1356;
    assign in1356_1 = {pp56[84]};
    assign in1356_2 = {pp57[83]};
    Full_Adder FA_1356(s1356, c1356, in1356_1, in1356_2, pp55[85]);
    wire[0:0] s1357, in1357_1, in1357_2;
    wire c1357;
    assign in1357_1 = {pp59[81]};
    assign in1357_2 = {pp60[80]};
    Full_Adder FA_1357(s1357, c1357, in1357_1, in1357_2, pp58[82]);
    wire[0:0] s1358, in1358_1, in1358_2;
    wire c1358;
    assign in1358_1 = {pp62[78]};
    assign in1358_2 = {pp63[77]};
    Full_Adder FA_1358(s1358, c1358, in1358_1, in1358_2, pp61[79]);
    wire[0:0] s1359, in1359_1, in1359_2;
    wire c1359;
    assign in1359_1 = {pp65[75]};
    assign in1359_2 = {pp66[74]};
    Full_Adder FA_1359(s1359, c1359, in1359_1, in1359_2, pp64[76]);
    wire[0:0] s1360, in1360_1, in1360_2;
    wire c1360;
    assign in1360_1 = {pp68[72]};
    assign in1360_2 = {pp69[71]};
    Full_Adder FA_1360(s1360, c1360, in1360_1, in1360_2, pp67[73]);
    wire[0:0] s1361, in1361_1, in1361_2;
    wire c1361;
    assign in1361_1 = {pp71[69]};
    assign in1361_2 = {pp72[68]};
    Full_Adder FA_1361(s1361, c1361, in1361_1, in1361_2, pp70[70]);
    wire[0:0] s1362, in1362_1, in1362_2;
    wire c1362;
    assign in1362_1 = {pp74[66]};
    assign in1362_2 = {pp75[65]};
    Full_Adder FA_1362(s1362, c1362, in1362_1, in1362_2, pp73[67]);
    wire[0:0] s1363, in1363_1, in1363_2;
    wire c1363;
    assign in1363_1 = {pp77[63]};
    assign in1363_2 = {pp78[62]};
    Full_Adder FA_1363(s1363, c1363, in1363_1, in1363_2, pp76[64]);
    wire[0:0] s1364, in1364_1, in1364_2;
    wire c1364;
    assign in1364_1 = {pp80[60]};
    assign in1364_2 = {pp81[59]};
    Full_Adder FA_1364(s1364, c1364, in1364_1, in1364_2, pp79[61]);
    wire[0:0] s1365, in1365_1, in1365_2;
    wire c1365;
    assign in1365_1 = {pp83[57]};
    assign in1365_2 = {pp84[56]};
    Full_Adder FA_1365(s1365, c1365, in1365_1, in1365_2, pp82[58]);
    wire[0:0] s1366, in1366_1, in1366_2;
    wire c1366;
    assign in1366_1 = {pp86[54]};
    assign in1366_2 = {pp87[53]};
    Full_Adder FA_1366(s1366, c1366, in1366_1, in1366_2, pp85[55]);
    wire[0:0] s1367, in1367_1, in1367_2;
    wire c1367;
    assign in1367_1 = {pp89[51]};
    assign in1367_2 = {pp90[50]};
    Full_Adder FA_1367(s1367, c1367, in1367_1, in1367_2, pp88[52]);
    wire[0:0] s1368, in1368_1, in1368_2;
    wire c1368;
    assign in1368_1 = {pp92[48]};
    assign in1368_2 = {pp93[47]};
    Full_Adder FA_1368(s1368, c1368, in1368_1, in1368_2, pp91[49]);
    wire[0:0] s1369, in1369_1, in1369_2;
    wire c1369;
    assign in1369_1 = {pp95[45]};
    assign in1369_2 = {pp96[44]};
    Full_Adder FA_1369(s1369, c1369, in1369_1, in1369_2, pp94[46]);
    wire[0:0] s1370, in1370_1, in1370_2;
    wire c1370;
    assign in1370_1 = {pp98[42]};
    assign in1370_2 = {pp99[41]};
    Full_Adder FA_1370(s1370, c1370, in1370_1, in1370_2, pp97[43]);
    wire[0:0] s1371, in1371_1, in1371_2;
    wire c1371;
    assign in1371_1 = {pp101[39]};
    assign in1371_2 = {pp102[38]};
    Full_Adder FA_1371(s1371, c1371, in1371_1, in1371_2, pp100[40]);
    wire[0:0] s1372, in1372_1, in1372_2;
    wire c1372;
    assign in1372_1 = {pp15[126]};
    assign in1372_2 = {pp16[125]};
    Full_Adder FA_1372(s1372, c1372, in1372_1, in1372_2, pp14[127]);
    wire[0:0] s1373, in1373_1, in1373_2;
    wire c1373;
    assign in1373_1 = {pp18[123]};
    assign in1373_2 = {pp19[122]};
    Full_Adder FA_1373(s1373, c1373, in1373_1, in1373_2, pp17[124]);
    wire[0:0] s1374, in1374_1, in1374_2;
    wire c1374;
    assign in1374_1 = {pp21[120]};
    assign in1374_2 = {pp22[119]};
    Full_Adder FA_1374(s1374, c1374, in1374_1, in1374_2, pp20[121]);
    wire[0:0] s1375, in1375_1, in1375_2;
    wire c1375;
    assign in1375_1 = {pp24[117]};
    assign in1375_2 = {pp25[116]};
    Full_Adder FA_1375(s1375, c1375, in1375_1, in1375_2, pp23[118]);
    wire[0:0] s1376, in1376_1, in1376_2;
    wire c1376;
    assign in1376_1 = {pp27[114]};
    assign in1376_2 = {pp28[113]};
    Full_Adder FA_1376(s1376, c1376, in1376_1, in1376_2, pp26[115]);
    wire[0:0] s1377, in1377_1, in1377_2;
    wire c1377;
    assign in1377_1 = {pp30[111]};
    assign in1377_2 = {pp31[110]};
    Full_Adder FA_1377(s1377, c1377, in1377_1, in1377_2, pp29[112]);
    wire[0:0] s1378, in1378_1, in1378_2;
    wire c1378;
    assign in1378_1 = {pp33[108]};
    assign in1378_2 = {pp34[107]};
    Full_Adder FA_1378(s1378, c1378, in1378_1, in1378_2, pp32[109]);
    wire[0:0] s1379, in1379_1, in1379_2;
    wire c1379;
    assign in1379_1 = {pp36[105]};
    assign in1379_2 = {pp37[104]};
    Full_Adder FA_1379(s1379, c1379, in1379_1, in1379_2, pp35[106]);
    wire[0:0] s1380, in1380_1, in1380_2;
    wire c1380;
    assign in1380_1 = {pp39[102]};
    assign in1380_2 = {pp40[101]};
    Full_Adder FA_1380(s1380, c1380, in1380_1, in1380_2, pp38[103]);
    wire[0:0] s1381, in1381_1, in1381_2;
    wire c1381;
    assign in1381_1 = {pp42[99]};
    assign in1381_2 = {pp43[98]};
    Full_Adder FA_1381(s1381, c1381, in1381_1, in1381_2, pp41[100]);
    wire[0:0] s1382, in1382_1, in1382_2;
    wire c1382;
    assign in1382_1 = {pp45[96]};
    assign in1382_2 = {pp46[95]};
    Full_Adder FA_1382(s1382, c1382, in1382_1, in1382_2, pp44[97]);
    wire[0:0] s1383, in1383_1, in1383_2;
    wire c1383;
    assign in1383_1 = {pp48[93]};
    assign in1383_2 = {pp49[92]};
    Full_Adder FA_1383(s1383, c1383, in1383_1, in1383_2, pp47[94]);
    wire[0:0] s1384, in1384_1, in1384_2;
    wire c1384;
    assign in1384_1 = {pp51[90]};
    assign in1384_2 = {pp52[89]};
    Full_Adder FA_1384(s1384, c1384, in1384_1, in1384_2, pp50[91]);
    wire[0:0] s1385, in1385_1, in1385_2;
    wire c1385;
    assign in1385_1 = {pp54[87]};
    assign in1385_2 = {pp55[86]};
    Full_Adder FA_1385(s1385, c1385, in1385_1, in1385_2, pp53[88]);
    wire[0:0] s1386, in1386_1, in1386_2;
    wire c1386;
    assign in1386_1 = {pp57[84]};
    assign in1386_2 = {pp58[83]};
    Full_Adder FA_1386(s1386, c1386, in1386_1, in1386_2, pp56[85]);
    wire[0:0] s1387, in1387_1, in1387_2;
    wire c1387;
    assign in1387_1 = {pp60[81]};
    assign in1387_2 = {pp61[80]};
    Full_Adder FA_1387(s1387, c1387, in1387_1, in1387_2, pp59[82]);
    wire[0:0] s1388, in1388_1, in1388_2;
    wire c1388;
    assign in1388_1 = {pp63[78]};
    assign in1388_2 = {pp64[77]};
    Full_Adder FA_1388(s1388, c1388, in1388_1, in1388_2, pp62[79]);
    wire[0:0] s1389, in1389_1, in1389_2;
    wire c1389;
    assign in1389_1 = {pp66[75]};
    assign in1389_2 = {pp67[74]};
    Full_Adder FA_1389(s1389, c1389, in1389_1, in1389_2, pp65[76]);
    wire[0:0] s1390, in1390_1, in1390_2;
    wire c1390;
    assign in1390_1 = {pp69[72]};
    assign in1390_2 = {pp70[71]};
    Full_Adder FA_1390(s1390, c1390, in1390_1, in1390_2, pp68[73]);
    wire[0:0] s1391, in1391_1, in1391_2;
    wire c1391;
    assign in1391_1 = {pp72[69]};
    assign in1391_2 = {pp73[68]};
    Full_Adder FA_1391(s1391, c1391, in1391_1, in1391_2, pp71[70]);
    wire[0:0] s1392, in1392_1, in1392_2;
    wire c1392;
    assign in1392_1 = {pp75[66]};
    assign in1392_2 = {pp76[65]};
    Full_Adder FA_1392(s1392, c1392, in1392_1, in1392_2, pp74[67]);
    wire[0:0] s1393, in1393_1, in1393_2;
    wire c1393;
    assign in1393_1 = {pp78[63]};
    assign in1393_2 = {pp79[62]};
    Full_Adder FA_1393(s1393, c1393, in1393_1, in1393_2, pp77[64]);
    wire[0:0] s1394, in1394_1, in1394_2;
    wire c1394;
    assign in1394_1 = {pp81[60]};
    assign in1394_2 = {pp82[59]};
    Full_Adder FA_1394(s1394, c1394, in1394_1, in1394_2, pp80[61]);
    wire[0:0] s1395, in1395_1, in1395_2;
    wire c1395;
    assign in1395_1 = {pp84[57]};
    assign in1395_2 = {pp85[56]};
    Full_Adder FA_1395(s1395, c1395, in1395_1, in1395_2, pp83[58]);
    wire[0:0] s1396, in1396_1, in1396_2;
    wire c1396;
    assign in1396_1 = {pp87[54]};
    assign in1396_2 = {pp88[53]};
    Full_Adder FA_1396(s1396, c1396, in1396_1, in1396_2, pp86[55]);
    wire[0:0] s1397, in1397_1, in1397_2;
    wire c1397;
    assign in1397_1 = {pp90[51]};
    assign in1397_2 = {pp91[50]};
    Full_Adder FA_1397(s1397, c1397, in1397_1, in1397_2, pp89[52]);
    wire[0:0] s1398, in1398_1, in1398_2;
    wire c1398;
    assign in1398_1 = {pp93[48]};
    assign in1398_2 = {pp94[47]};
    Full_Adder FA_1398(s1398, c1398, in1398_1, in1398_2, pp92[49]);
    wire[0:0] s1399, in1399_1, in1399_2;
    wire c1399;
    assign in1399_1 = {pp96[45]};
    assign in1399_2 = {pp97[44]};
    Full_Adder FA_1399(s1399, c1399, in1399_1, in1399_2, pp95[46]);
    wire[0:0] s1400, in1400_1, in1400_2;
    wire c1400;
    assign in1400_1 = {pp99[42]};
    assign in1400_2 = {pp100[41]};
    Full_Adder FA_1400(s1400, c1400, in1400_1, in1400_2, pp98[43]);
    wire[0:0] s1401, in1401_1, in1401_2;
    wire c1401;
    assign in1401_1 = {pp16[126]};
    assign in1401_2 = {pp17[125]};
    Full_Adder FA_1401(s1401, c1401, in1401_1, in1401_2, pp15[127]);
    wire[0:0] s1402, in1402_1, in1402_2;
    wire c1402;
    assign in1402_1 = {pp19[123]};
    assign in1402_2 = {pp20[122]};
    Full_Adder FA_1402(s1402, c1402, in1402_1, in1402_2, pp18[124]);
    wire[0:0] s1403, in1403_1, in1403_2;
    wire c1403;
    assign in1403_1 = {pp22[120]};
    assign in1403_2 = {pp23[119]};
    Full_Adder FA_1403(s1403, c1403, in1403_1, in1403_2, pp21[121]);
    wire[0:0] s1404, in1404_1, in1404_2;
    wire c1404;
    assign in1404_1 = {pp25[117]};
    assign in1404_2 = {pp26[116]};
    Full_Adder FA_1404(s1404, c1404, in1404_1, in1404_2, pp24[118]);
    wire[0:0] s1405, in1405_1, in1405_2;
    wire c1405;
    assign in1405_1 = {pp28[114]};
    assign in1405_2 = {pp29[113]};
    Full_Adder FA_1405(s1405, c1405, in1405_1, in1405_2, pp27[115]);
    wire[0:0] s1406, in1406_1, in1406_2;
    wire c1406;
    assign in1406_1 = {pp31[111]};
    assign in1406_2 = {pp32[110]};
    Full_Adder FA_1406(s1406, c1406, in1406_1, in1406_2, pp30[112]);
    wire[0:0] s1407, in1407_1, in1407_2;
    wire c1407;
    assign in1407_1 = {pp34[108]};
    assign in1407_2 = {pp35[107]};
    Full_Adder FA_1407(s1407, c1407, in1407_1, in1407_2, pp33[109]);
    wire[0:0] s1408, in1408_1, in1408_2;
    wire c1408;
    assign in1408_1 = {pp37[105]};
    assign in1408_2 = {pp38[104]};
    Full_Adder FA_1408(s1408, c1408, in1408_1, in1408_2, pp36[106]);
    wire[0:0] s1409, in1409_1, in1409_2;
    wire c1409;
    assign in1409_1 = {pp40[102]};
    assign in1409_2 = {pp41[101]};
    Full_Adder FA_1409(s1409, c1409, in1409_1, in1409_2, pp39[103]);
    wire[0:0] s1410, in1410_1, in1410_2;
    wire c1410;
    assign in1410_1 = {pp43[99]};
    assign in1410_2 = {pp44[98]};
    Full_Adder FA_1410(s1410, c1410, in1410_1, in1410_2, pp42[100]);
    wire[0:0] s1411, in1411_1, in1411_2;
    wire c1411;
    assign in1411_1 = {pp46[96]};
    assign in1411_2 = {pp47[95]};
    Full_Adder FA_1411(s1411, c1411, in1411_1, in1411_2, pp45[97]);
    wire[0:0] s1412, in1412_1, in1412_2;
    wire c1412;
    assign in1412_1 = {pp49[93]};
    assign in1412_2 = {pp50[92]};
    Full_Adder FA_1412(s1412, c1412, in1412_1, in1412_2, pp48[94]);
    wire[0:0] s1413, in1413_1, in1413_2;
    wire c1413;
    assign in1413_1 = {pp52[90]};
    assign in1413_2 = {pp53[89]};
    Full_Adder FA_1413(s1413, c1413, in1413_1, in1413_2, pp51[91]);
    wire[0:0] s1414, in1414_1, in1414_2;
    wire c1414;
    assign in1414_1 = {pp55[87]};
    assign in1414_2 = {pp56[86]};
    Full_Adder FA_1414(s1414, c1414, in1414_1, in1414_2, pp54[88]);
    wire[0:0] s1415, in1415_1, in1415_2;
    wire c1415;
    assign in1415_1 = {pp58[84]};
    assign in1415_2 = {pp59[83]};
    Full_Adder FA_1415(s1415, c1415, in1415_1, in1415_2, pp57[85]);
    wire[0:0] s1416, in1416_1, in1416_2;
    wire c1416;
    assign in1416_1 = {pp61[81]};
    assign in1416_2 = {pp62[80]};
    Full_Adder FA_1416(s1416, c1416, in1416_1, in1416_2, pp60[82]);
    wire[0:0] s1417, in1417_1, in1417_2;
    wire c1417;
    assign in1417_1 = {pp64[78]};
    assign in1417_2 = {pp65[77]};
    Full_Adder FA_1417(s1417, c1417, in1417_1, in1417_2, pp63[79]);
    wire[0:0] s1418, in1418_1, in1418_2;
    wire c1418;
    assign in1418_1 = {pp67[75]};
    assign in1418_2 = {pp68[74]};
    Full_Adder FA_1418(s1418, c1418, in1418_1, in1418_2, pp66[76]);
    wire[0:0] s1419, in1419_1, in1419_2;
    wire c1419;
    assign in1419_1 = {pp70[72]};
    assign in1419_2 = {pp71[71]};
    Full_Adder FA_1419(s1419, c1419, in1419_1, in1419_2, pp69[73]);
    wire[0:0] s1420, in1420_1, in1420_2;
    wire c1420;
    assign in1420_1 = {pp73[69]};
    assign in1420_2 = {pp74[68]};
    Full_Adder FA_1420(s1420, c1420, in1420_1, in1420_2, pp72[70]);
    wire[0:0] s1421, in1421_1, in1421_2;
    wire c1421;
    assign in1421_1 = {pp76[66]};
    assign in1421_2 = {pp77[65]};
    Full_Adder FA_1421(s1421, c1421, in1421_1, in1421_2, pp75[67]);
    wire[0:0] s1422, in1422_1, in1422_2;
    wire c1422;
    assign in1422_1 = {pp79[63]};
    assign in1422_2 = {pp80[62]};
    Full_Adder FA_1422(s1422, c1422, in1422_1, in1422_2, pp78[64]);
    wire[0:0] s1423, in1423_1, in1423_2;
    wire c1423;
    assign in1423_1 = {pp82[60]};
    assign in1423_2 = {pp83[59]};
    Full_Adder FA_1423(s1423, c1423, in1423_1, in1423_2, pp81[61]);
    wire[0:0] s1424, in1424_1, in1424_2;
    wire c1424;
    assign in1424_1 = {pp85[57]};
    assign in1424_2 = {pp86[56]};
    Full_Adder FA_1424(s1424, c1424, in1424_1, in1424_2, pp84[58]);
    wire[0:0] s1425, in1425_1, in1425_2;
    wire c1425;
    assign in1425_1 = {pp88[54]};
    assign in1425_2 = {pp89[53]};
    Full_Adder FA_1425(s1425, c1425, in1425_1, in1425_2, pp87[55]);
    wire[0:0] s1426, in1426_1, in1426_2;
    wire c1426;
    assign in1426_1 = {pp91[51]};
    assign in1426_2 = {pp92[50]};
    Full_Adder FA_1426(s1426, c1426, in1426_1, in1426_2, pp90[52]);
    wire[0:0] s1427, in1427_1, in1427_2;
    wire c1427;
    assign in1427_1 = {pp94[48]};
    assign in1427_2 = {pp95[47]};
    Full_Adder FA_1427(s1427, c1427, in1427_1, in1427_2, pp93[49]);
    wire[0:0] s1428, in1428_1, in1428_2;
    wire c1428;
    assign in1428_1 = {pp97[45]};
    assign in1428_2 = {pp98[44]};
    Full_Adder FA_1428(s1428, c1428, in1428_1, in1428_2, pp96[46]);
    wire[0:0] s1429, in1429_1, in1429_2;
    wire c1429;
    assign in1429_1 = {pp17[126]};
    assign in1429_2 = {pp18[125]};
    Full_Adder FA_1429(s1429, c1429, in1429_1, in1429_2, pp16[127]);
    wire[0:0] s1430, in1430_1, in1430_2;
    wire c1430;
    assign in1430_1 = {pp20[123]};
    assign in1430_2 = {pp21[122]};
    Full_Adder FA_1430(s1430, c1430, in1430_1, in1430_2, pp19[124]);
    wire[0:0] s1431, in1431_1, in1431_2;
    wire c1431;
    assign in1431_1 = {pp23[120]};
    assign in1431_2 = {pp24[119]};
    Full_Adder FA_1431(s1431, c1431, in1431_1, in1431_2, pp22[121]);
    wire[0:0] s1432, in1432_1, in1432_2;
    wire c1432;
    assign in1432_1 = {pp26[117]};
    assign in1432_2 = {pp27[116]};
    Full_Adder FA_1432(s1432, c1432, in1432_1, in1432_2, pp25[118]);
    wire[0:0] s1433, in1433_1, in1433_2;
    wire c1433;
    assign in1433_1 = {pp29[114]};
    assign in1433_2 = {pp30[113]};
    Full_Adder FA_1433(s1433, c1433, in1433_1, in1433_2, pp28[115]);
    wire[0:0] s1434, in1434_1, in1434_2;
    wire c1434;
    assign in1434_1 = {pp32[111]};
    assign in1434_2 = {pp33[110]};
    Full_Adder FA_1434(s1434, c1434, in1434_1, in1434_2, pp31[112]);
    wire[0:0] s1435, in1435_1, in1435_2;
    wire c1435;
    assign in1435_1 = {pp35[108]};
    assign in1435_2 = {pp36[107]};
    Full_Adder FA_1435(s1435, c1435, in1435_1, in1435_2, pp34[109]);
    wire[0:0] s1436, in1436_1, in1436_2;
    wire c1436;
    assign in1436_1 = {pp38[105]};
    assign in1436_2 = {pp39[104]};
    Full_Adder FA_1436(s1436, c1436, in1436_1, in1436_2, pp37[106]);
    wire[0:0] s1437, in1437_1, in1437_2;
    wire c1437;
    assign in1437_1 = {pp41[102]};
    assign in1437_2 = {pp42[101]};
    Full_Adder FA_1437(s1437, c1437, in1437_1, in1437_2, pp40[103]);
    wire[0:0] s1438, in1438_1, in1438_2;
    wire c1438;
    assign in1438_1 = {pp44[99]};
    assign in1438_2 = {pp45[98]};
    Full_Adder FA_1438(s1438, c1438, in1438_1, in1438_2, pp43[100]);
    wire[0:0] s1439, in1439_1, in1439_2;
    wire c1439;
    assign in1439_1 = {pp47[96]};
    assign in1439_2 = {pp48[95]};
    Full_Adder FA_1439(s1439, c1439, in1439_1, in1439_2, pp46[97]);
    wire[0:0] s1440, in1440_1, in1440_2;
    wire c1440;
    assign in1440_1 = {pp50[93]};
    assign in1440_2 = {pp51[92]};
    Full_Adder FA_1440(s1440, c1440, in1440_1, in1440_2, pp49[94]);
    wire[0:0] s1441, in1441_1, in1441_2;
    wire c1441;
    assign in1441_1 = {pp53[90]};
    assign in1441_2 = {pp54[89]};
    Full_Adder FA_1441(s1441, c1441, in1441_1, in1441_2, pp52[91]);
    wire[0:0] s1442, in1442_1, in1442_2;
    wire c1442;
    assign in1442_1 = {pp56[87]};
    assign in1442_2 = {pp57[86]};
    Full_Adder FA_1442(s1442, c1442, in1442_1, in1442_2, pp55[88]);
    wire[0:0] s1443, in1443_1, in1443_2;
    wire c1443;
    assign in1443_1 = {pp59[84]};
    assign in1443_2 = {pp60[83]};
    Full_Adder FA_1443(s1443, c1443, in1443_1, in1443_2, pp58[85]);
    wire[0:0] s1444, in1444_1, in1444_2;
    wire c1444;
    assign in1444_1 = {pp62[81]};
    assign in1444_2 = {pp63[80]};
    Full_Adder FA_1444(s1444, c1444, in1444_1, in1444_2, pp61[82]);
    wire[0:0] s1445, in1445_1, in1445_2;
    wire c1445;
    assign in1445_1 = {pp65[78]};
    assign in1445_2 = {pp66[77]};
    Full_Adder FA_1445(s1445, c1445, in1445_1, in1445_2, pp64[79]);
    wire[0:0] s1446, in1446_1, in1446_2;
    wire c1446;
    assign in1446_1 = {pp68[75]};
    assign in1446_2 = {pp69[74]};
    Full_Adder FA_1446(s1446, c1446, in1446_1, in1446_2, pp67[76]);
    wire[0:0] s1447, in1447_1, in1447_2;
    wire c1447;
    assign in1447_1 = {pp71[72]};
    assign in1447_2 = {pp72[71]};
    Full_Adder FA_1447(s1447, c1447, in1447_1, in1447_2, pp70[73]);
    wire[0:0] s1448, in1448_1, in1448_2;
    wire c1448;
    assign in1448_1 = {pp74[69]};
    assign in1448_2 = {pp75[68]};
    Full_Adder FA_1448(s1448, c1448, in1448_1, in1448_2, pp73[70]);
    wire[0:0] s1449, in1449_1, in1449_2;
    wire c1449;
    assign in1449_1 = {pp77[66]};
    assign in1449_2 = {pp78[65]};
    Full_Adder FA_1449(s1449, c1449, in1449_1, in1449_2, pp76[67]);
    wire[0:0] s1450, in1450_1, in1450_2;
    wire c1450;
    assign in1450_1 = {pp80[63]};
    assign in1450_2 = {pp81[62]};
    Full_Adder FA_1450(s1450, c1450, in1450_1, in1450_2, pp79[64]);
    wire[0:0] s1451, in1451_1, in1451_2;
    wire c1451;
    assign in1451_1 = {pp83[60]};
    assign in1451_2 = {pp84[59]};
    Full_Adder FA_1451(s1451, c1451, in1451_1, in1451_2, pp82[61]);
    wire[0:0] s1452, in1452_1, in1452_2;
    wire c1452;
    assign in1452_1 = {pp86[57]};
    assign in1452_2 = {pp87[56]};
    Full_Adder FA_1452(s1452, c1452, in1452_1, in1452_2, pp85[58]);
    wire[0:0] s1453, in1453_1, in1453_2;
    wire c1453;
    assign in1453_1 = {pp89[54]};
    assign in1453_2 = {pp90[53]};
    Full_Adder FA_1453(s1453, c1453, in1453_1, in1453_2, pp88[55]);
    wire[0:0] s1454, in1454_1, in1454_2;
    wire c1454;
    assign in1454_1 = {pp92[51]};
    assign in1454_2 = {pp93[50]};
    Full_Adder FA_1454(s1454, c1454, in1454_1, in1454_2, pp91[52]);
    wire[0:0] s1455, in1455_1, in1455_2;
    wire c1455;
    assign in1455_1 = {pp95[48]};
    assign in1455_2 = {pp96[47]};
    Full_Adder FA_1455(s1455, c1455, in1455_1, in1455_2, pp94[49]);
    wire[0:0] s1456, in1456_1, in1456_2;
    wire c1456;
    assign in1456_1 = {pp18[126]};
    assign in1456_2 = {pp19[125]};
    Full_Adder FA_1456(s1456, c1456, in1456_1, in1456_2, pp17[127]);
    wire[0:0] s1457, in1457_1, in1457_2;
    wire c1457;
    assign in1457_1 = {pp21[123]};
    assign in1457_2 = {pp22[122]};
    Full_Adder FA_1457(s1457, c1457, in1457_1, in1457_2, pp20[124]);
    wire[0:0] s1458, in1458_1, in1458_2;
    wire c1458;
    assign in1458_1 = {pp24[120]};
    assign in1458_2 = {pp25[119]};
    Full_Adder FA_1458(s1458, c1458, in1458_1, in1458_2, pp23[121]);
    wire[0:0] s1459, in1459_1, in1459_2;
    wire c1459;
    assign in1459_1 = {pp27[117]};
    assign in1459_2 = {pp28[116]};
    Full_Adder FA_1459(s1459, c1459, in1459_1, in1459_2, pp26[118]);
    wire[0:0] s1460, in1460_1, in1460_2;
    wire c1460;
    assign in1460_1 = {pp30[114]};
    assign in1460_2 = {pp31[113]};
    Full_Adder FA_1460(s1460, c1460, in1460_1, in1460_2, pp29[115]);
    wire[0:0] s1461, in1461_1, in1461_2;
    wire c1461;
    assign in1461_1 = {pp33[111]};
    assign in1461_2 = {pp34[110]};
    Full_Adder FA_1461(s1461, c1461, in1461_1, in1461_2, pp32[112]);
    wire[0:0] s1462, in1462_1, in1462_2;
    wire c1462;
    assign in1462_1 = {pp36[108]};
    assign in1462_2 = {pp37[107]};
    Full_Adder FA_1462(s1462, c1462, in1462_1, in1462_2, pp35[109]);
    wire[0:0] s1463, in1463_1, in1463_2;
    wire c1463;
    assign in1463_1 = {pp39[105]};
    assign in1463_2 = {pp40[104]};
    Full_Adder FA_1463(s1463, c1463, in1463_1, in1463_2, pp38[106]);
    wire[0:0] s1464, in1464_1, in1464_2;
    wire c1464;
    assign in1464_1 = {pp42[102]};
    assign in1464_2 = {pp43[101]};
    Full_Adder FA_1464(s1464, c1464, in1464_1, in1464_2, pp41[103]);
    wire[0:0] s1465, in1465_1, in1465_2;
    wire c1465;
    assign in1465_1 = {pp45[99]};
    assign in1465_2 = {pp46[98]};
    Full_Adder FA_1465(s1465, c1465, in1465_1, in1465_2, pp44[100]);
    wire[0:0] s1466, in1466_1, in1466_2;
    wire c1466;
    assign in1466_1 = {pp48[96]};
    assign in1466_2 = {pp49[95]};
    Full_Adder FA_1466(s1466, c1466, in1466_1, in1466_2, pp47[97]);
    wire[0:0] s1467, in1467_1, in1467_2;
    wire c1467;
    assign in1467_1 = {pp51[93]};
    assign in1467_2 = {pp52[92]};
    Full_Adder FA_1467(s1467, c1467, in1467_1, in1467_2, pp50[94]);
    wire[0:0] s1468, in1468_1, in1468_2;
    wire c1468;
    assign in1468_1 = {pp54[90]};
    assign in1468_2 = {pp55[89]};
    Full_Adder FA_1468(s1468, c1468, in1468_1, in1468_2, pp53[91]);
    wire[0:0] s1469, in1469_1, in1469_2;
    wire c1469;
    assign in1469_1 = {pp57[87]};
    assign in1469_2 = {pp58[86]};
    Full_Adder FA_1469(s1469, c1469, in1469_1, in1469_2, pp56[88]);
    wire[0:0] s1470, in1470_1, in1470_2;
    wire c1470;
    assign in1470_1 = {pp60[84]};
    assign in1470_2 = {pp61[83]};
    Full_Adder FA_1470(s1470, c1470, in1470_1, in1470_2, pp59[85]);
    wire[0:0] s1471, in1471_1, in1471_2;
    wire c1471;
    assign in1471_1 = {pp63[81]};
    assign in1471_2 = {pp64[80]};
    Full_Adder FA_1471(s1471, c1471, in1471_1, in1471_2, pp62[82]);
    wire[0:0] s1472, in1472_1, in1472_2;
    wire c1472;
    assign in1472_1 = {pp66[78]};
    assign in1472_2 = {pp67[77]};
    Full_Adder FA_1472(s1472, c1472, in1472_1, in1472_2, pp65[79]);
    wire[0:0] s1473, in1473_1, in1473_2;
    wire c1473;
    assign in1473_1 = {pp69[75]};
    assign in1473_2 = {pp70[74]};
    Full_Adder FA_1473(s1473, c1473, in1473_1, in1473_2, pp68[76]);
    wire[0:0] s1474, in1474_1, in1474_2;
    wire c1474;
    assign in1474_1 = {pp72[72]};
    assign in1474_2 = {pp73[71]};
    Full_Adder FA_1474(s1474, c1474, in1474_1, in1474_2, pp71[73]);
    wire[0:0] s1475, in1475_1, in1475_2;
    wire c1475;
    assign in1475_1 = {pp75[69]};
    assign in1475_2 = {pp76[68]};
    Full_Adder FA_1475(s1475, c1475, in1475_1, in1475_2, pp74[70]);
    wire[0:0] s1476, in1476_1, in1476_2;
    wire c1476;
    assign in1476_1 = {pp78[66]};
    assign in1476_2 = {pp79[65]};
    Full_Adder FA_1476(s1476, c1476, in1476_1, in1476_2, pp77[67]);
    wire[0:0] s1477, in1477_1, in1477_2;
    wire c1477;
    assign in1477_1 = {pp81[63]};
    assign in1477_2 = {pp82[62]};
    Full_Adder FA_1477(s1477, c1477, in1477_1, in1477_2, pp80[64]);
    wire[0:0] s1478, in1478_1, in1478_2;
    wire c1478;
    assign in1478_1 = {pp84[60]};
    assign in1478_2 = {pp85[59]};
    Full_Adder FA_1478(s1478, c1478, in1478_1, in1478_2, pp83[61]);
    wire[0:0] s1479, in1479_1, in1479_2;
    wire c1479;
    assign in1479_1 = {pp87[57]};
    assign in1479_2 = {pp88[56]};
    Full_Adder FA_1479(s1479, c1479, in1479_1, in1479_2, pp86[58]);
    wire[0:0] s1480, in1480_1, in1480_2;
    wire c1480;
    assign in1480_1 = {pp90[54]};
    assign in1480_2 = {pp91[53]};
    Full_Adder FA_1480(s1480, c1480, in1480_1, in1480_2, pp89[55]);
    wire[0:0] s1481, in1481_1, in1481_2;
    wire c1481;
    assign in1481_1 = {pp93[51]};
    assign in1481_2 = {pp94[50]};
    Full_Adder FA_1481(s1481, c1481, in1481_1, in1481_2, pp92[52]);
    wire[0:0] s1482, in1482_1, in1482_2;
    wire c1482;
    assign in1482_1 = {pp19[126]};
    assign in1482_2 = {pp20[125]};
    Full_Adder FA_1482(s1482, c1482, in1482_1, in1482_2, pp18[127]);
    wire[0:0] s1483, in1483_1, in1483_2;
    wire c1483;
    assign in1483_1 = {pp22[123]};
    assign in1483_2 = {pp23[122]};
    Full_Adder FA_1483(s1483, c1483, in1483_1, in1483_2, pp21[124]);
    wire[0:0] s1484, in1484_1, in1484_2;
    wire c1484;
    assign in1484_1 = {pp25[120]};
    assign in1484_2 = {pp26[119]};
    Full_Adder FA_1484(s1484, c1484, in1484_1, in1484_2, pp24[121]);
    wire[0:0] s1485, in1485_1, in1485_2;
    wire c1485;
    assign in1485_1 = {pp28[117]};
    assign in1485_2 = {pp29[116]};
    Full_Adder FA_1485(s1485, c1485, in1485_1, in1485_2, pp27[118]);
    wire[0:0] s1486, in1486_1, in1486_2;
    wire c1486;
    assign in1486_1 = {pp31[114]};
    assign in1486_2 = {pp32[113]};
    Full_Adder FA_1486(s1486, c1486, in1486_1, in1486_2, pp30[115]);
    wire[0:0] s1487, in1487_1, in1487_2;
    wire c1487;
    assign in1487_1 = {pp34[111]};
    assign in1487_2 = {pp35[110]};
    Full_Adder FA_1487(s1487, c1487, in1487_1, in1487_2, pp33[112]);
    wire[0:0] s1488, in1488_1, in1488_2;
    wire c1488;
    assign in1488_1 = {pp37[108]};
    assign in1488_2 = {pp38[107]};
    Full_Adder FA_1488(s1488, c1488, in1488_1, in1488_2, pp36[109]);
    wire[0:0] s1489, in1489_1, in1489_2;
    wire c1489;
    assign in1489_1 = {pp40[105]};
    assign in1489_2 = {pp41[104]};
    Full_Adder FA_1489(s1489, c1489, in1489_1, in1489_2, pp39[106]);
    wire[0:0] s1490, in1490_1, in1490_2;
    wire c1490;
    assign in1490_1 = {pp43[102]};
    assign in1490_2 = {pp44[101]};
    Full_Adder FA_1490(s1490, c1490, in1490_1, in1490_2, pp42[103]);
    wire[0:0] s1491, in1491_1, in1491_2;
    wire c1491;
    assign in1491_1 = {pp46[99]};
    assign in1491_2 = {pp47[98]};
    Full_Adder FA_1491(s1491, c1491, in1491_1, in1491_2, pp45[100]);
    wire[0:0] s1492, in1492_1, in1492_2;
    wire c1492;
    assign in1492_1 = {pp49[96]};
    assign in1492_2 = {pp50[95]};
    Full_Adder FA_1492(s1492, c1492, in1492_1, in1492_2, pp48[97]);
    wire[0:0] s1493, in1493_1, in1493_2;
    wire c1493;
    assign in1493_1 = {pp52[93]};
    assign in1493_2 = {pp53[92]};
    Full_Adder FA_1493(s1493, c1493, in1493_1, in1493_2, pp51[94]);
    wire[0:0] s1494, in1494_1, in1494_2;
    wire c1494;
    assign in1494_1 = {pp55[90]};
    assign in1494_2 = {pp56[89]};
    Full_Adder FA_1494(s1494, c1494, in1494_1, in1494_2, pp54[91]);
    wire[0:0] s1495, in1495_1, in1495_2;
    wire c1495;
    assign in1495_1 = {pp58[87]};
    assign in1495_2 = {pp59[86]};
    Full_Adder FA_1495(s1495, c1495, in1495_1, in1495_2, pp57[88]);
    wire[0:0] s1496, in1496_1, in1496_2;
    wire c1496;
    assign in1496_1 = {pp61[84]};
    assign in1496_2 = {pp62[83]};
    Full_Adder FA_1496(s1496, c1496, in1496_1, in1496_2, pp60[85]);
    wire[0:0] s1497, in1497_1, in1497_2;
    wire c1497;
    assign in1497_1 = {pp64[81]};
    assign in1497_2 = {pp65[80]};
    Full_Adder FA_1497(s1497, c1497, in1497_1, in1497_2, pp63[82]);
    wire[0:0] s1498, in1498_1, in1498_2;
    wire c1498;
    assign in1498_1 = {pp67[78]};
    assign in1498_2 = {pp68[77]};
    Full_Adder FA_1498(s1498, c1498, in1498_1, in1498_2, pp66[79]);
    wire[0:0] s1499, in1499_1, in1499_2;
    wire c1499;
    assign in1499_1 = {pp70[75]};
    assign in1499_2 = {pp71[74]};
    Full_Adder FA_1499(s1499, c1499, in1499_1, in1499_2, pp69[76]);
    wire[0:0] s1500, in1500_1, in1500_2;
    wire c1500;
    assign in1500_1 = {pp73[72]};
    assign in1500_2 = {pp74[71]};
    Full_Adder FA_1500(s1500, c1500, in1500_1, in1500_2, pp72[73]);
    wire[0:0] s1501, in1501_1, in1501_2;
    wire c1501;
    assign in1501_1 = {pp76[69]};
    assign in1501_2 = {pp77[68]};
    Full_Adder FA_1501(s1501, c1501, in1501_1, in1501_2, pp75[70]);
    wire[0:0] s1502, in1502_1, in1502_2;
    wire c1502;
    assign in1502_1 = {pp79[66]};
    assign in1502_2 = {pp80[65]};
    Full_Adder FA_1502(s1502, c1502, in1502_1, in1502_2, pp78[67]);
    wire[0:0] s1503, in1503_1, in1503_2;
    wire c1503;
    assign in1503_1 = {pp82[63]};
    assign in1503_2 = {pp83[62]};
    Full_Adder FA_1503(s1503, c1503, in1503_1, in1503_2, pp81[64]);
    wire[0:0] s1504, in1504_1, in1504_2;
    wire c1504;
    assign in1504_1 = {pp85[60]};
    assign in1504_2 = {pp86[59]};
    Full_Adder FA_1504(s1504, c1504, in1504_1, in1504_2, pp84[61]);
    wire[0:0] s1505, in1505_1, in1505_2;
    wire c1505;
    assign in1505_1 = {pp88[57]};
    assign in1505_2 = {pp89[56]};
    Full_Adder FA_1505(s1505, c1505, in1505_1, in1505_2, pp87[58]);
    wire[0:0] s1506, in1506_1, in1506_2;
    wire c1506;
    assign in1506_1 = {pp91[54]};
    assign in1506_2 = {pp92[53]};
    Full_Adder FA_1506(s1506, c1506, in1506_1, in1506_2, pp90[55]);
    wire[0:0] s1507, in1507_1, in1507_2;
    wire c1507;
    assign in1507_1 = {pp20[126]};
    assign in1507_2 = {pp21[125]};
    Full_Adder FA_1507(s1507, c1507, in1507_1, in1507_2, pp19[127]);
    wire[0:0] s1508, in1508_1, in1508_2;
    wire c1508;
    assign in1508_1 = {pp23[123]};
    assign in1508_2 = {pp24[122]};
    Full_Adder FA_1508(s1508, c1508, in1508_1, in1508_2, pp22[124]);
    wire[0:0] s1509, in1509_1, in1509_2;
    wire c1509;
    assign in1509_1 = {pp26[120]};
    assign in1509_2 = {pp27[119]};
    Full_Adder FA_1509(s1509, c1509, in1509_1, in1509_2, pp25[121]);
    wire[0:0] s1510, in1510_1, in1510_2;
    wire c1510;
    assign in1510_1 = {pp29[117]};
    assign in1510_2 = {pp30[116]};
    Full_Adder FA_1510(s1510, c1510, in1510_1, in1510_2, pp28[118]);
    wire[0:0] s1511, in1511_1, in1511_2;
    wire c1511;
    assign in1511_1 = {pp32[114]};
    assign in1511_2 = {pp33[113]};
    Full_Adder FA_1511(s1511, c1511, in1511_1, in1511_2, pp31[115]);
    wire[0:0] s1512, in1512_1, in1512_2;
    wire c1512;
    assign in1512_1 = {pp35[111]};
    assign in1512_2 = {pp36[110]};
    Full_Adder FA_1512(s1512, c1512, in1512_1, in1512_2, pp34[112]);
    wire[0:0] s1513, in1513_1, in1513_2;
    wire c1513;
    assign in1513_1 = {pp38[108]};
    assign in1513_2 = {pp39[107]};
    Full_Adder FA_1513(s1513, c1513, in1513_1, in1513_2, pp37[109]);
    wire[0:0] s1514, in1514_1, in1514_2;
    wire c1514;
    assign in1514_1 = {pp41[105]};
    assign in1514_2 = {pp42[104]};
    Full_Adder FA_1514(s1514, c1514, in1514_1, in1514_2, pp40[106]);
    wire[0:0] s1515, in1515_1, in1515_2;
    wire c1515;
    assign in1515_1 = {pp44[102]};
    assign in1515_2 = {pp45[101]};
    Full_Adder FA_1515(s1515, c1515, in1515_1, in1515_2, pp43[103]);
    wire[0:0] s1516, in1516_1, in1516_2;
    wire c1516;
    assign in1516_1 = {pp47[99]};
    assign in1516_2 = {pp48[98]};
    Full_Adder FA_1516(s1516, c1516, in1516_1, in1516_2, pp46[100]);
    wire[0:0] s1517, in1517_1, in1517_2;
    wire c1517;
    assign in1517_1 = {pp50[96]};
    assign in1517_2 = {pp51[95]};
    Full_Adder FA_1517(s1517, c1517, in1517_1, in1517_2, pp49[97]);
    wire[0:0] s1518, in1518_1, in1518_2;
    wire c1518;
    assign in1518_1 = {pp53[93]};
    assign in1518_2 = {pp54[92]};
    Full_Adder FA_1518(s1518, c1518, in1518_1, in1518_2, pp52[94]);
    wire[0:0] s1519, in1519_1, in1519_2;
    wire c1519;
    assign in1519_1 = {pp56[90]};
    assign in1519_2 = {pp57[89]};
    Full_Adder FA_1519(s1519, c1519, in1519_1, in1519_2, pp55[91]);
    wire[0:0] s1520, in1520_1, in1520_2;
    wire c1520;
    assign in1520_1 = {pp59[87]};
    assign in1520_2 = {pp60[86]};
    Full_Adder FA_1520(s1520, c1520, in1520_1, in1520_2, pp58[88]);
    wire[0:0] s1521, in1521_1, in1521_2;
    wire c1521;
    assign in1521_1 = {pp62[84]};
    assign in1521_2 = {pp63[83]};
    Full_Adder FA_1521(s1521, c1521, in1521_1, in1521_2, pp61[85]);
    wire[0:0] s1522, in1522_1, in1522_2;
    wire c1522;
    assign in1522_1 = {pp65[81]};
    assign in1522_2 = {pp66[80]};
    Full_Adder FA_1522(s1522, c1522, in1522_1, in1522_2, pp64[82]);
    wire[0:0] s1523, in1523_1, in1523_2;
    wire c1523;
    assign in1523_1 = {pp68[78]};
    assign in1523_2 = {pp69[77]};
    Full_Adder FA_1523(s1523, c1523, in1523_1, in1523_2, pp67[79]);
    wire[0:0] s1524, in1524_1, in1524_2;
    wire c1524;
    assign in1524_1 = {pp71[75]};
    assign in1524_2 = {pp72[74]};
    Full_Adder FA_1524(s1524, c1524, in1524_1, in1524_2, pp70[76]);
    wire[0:0] s1525, in1525_1, in1525_2;
    wire c1525;
    assign in1525_1 = {pp74[72]};
    assign in1525_2 = {pp75[71]};
    Full_Adder FA_1525(s1525, c1525, in1525_1, in1525_2, pp73[73]);
    wire[0:0] s1526, in1526_1, in1526_2;
    wire c1526;
    assign in1526_1 = {pp77[69]};
    assign in1526_2 = {pp78[68]};
    Full_Adder FA_1526(s1526, c1526, in1526_1, in1526_2, pp76[70]);
    wire[0:0] s1527, in1527_1, in1527_2;
    wire c1527;
    assign in1527_1 = {pp80[66]};
    assign in1527_2 = {pp81[65]};
    Full_Adder FA_1527(s1527, c1527, in1527_1, in1527_2, pp79[67]);
    wire[0:0] s1528, in1528_1, in1528_2;
    wire c1528;
    assign in1528_1 = {pp83[63]};
    assign in1528_2 = {pp84[62]};
    Full_Adder FA_1528(s1528, c1528, in1528_1, in1528_2, pp82[64]);
    wire[0:0] s1529, in1529_1, in1529_2;
    wire c1529;
    assign in1529_1 = {pp86[60]};
    assign in1529_2 = {pp87[59]};
    Full_Adder FA_1529(s1529, c1529, in1529_1, in1529_2, pp85[61]);
    wire[0:0] s1530, in1530_1, in1530_2;
    wire c1530;
    assign in1530_1 = {pp89[57]};
    assign in1530_2 = {pp90[56]};
    Full_Adder FA_1530(s1530, c1530, in1530_1, in1530_2, pp88[58]);
    wire[0:0] s1531, in1531_1, in1531_2;
    wire c1531;
    assign in1531_1 = {pp21[126]};
    assign in1531_2 = {pp22[125]};
    Full_Adder FA_1531(s1531, c1531, in1531_1, in1531_2, pp20[127]);
    wire[0:0] s1532, in1532_1, in1532_2;
    wire c1532;
    assign in1532_1 = {pp24[123]};
    assign in1532_2 = {pp25[122]};
    Full_Adder FA_1532(s1532, c1532, in1532_1, in1532_2, pp23[124]);
    wire[0:0] s1533, in1533_1, in1533_2;
    wire c1533;
    assign in1533_1 = {pp27[120]};
    assign in1533_2 = {pp28[119]};
    Full_Adder FA_1533(s1533, c1533, in1533_1, in1533_2, pp26[121]);
    wire[0:0] s1534, in1534_1, in1534_2;
    wire c1534;
    assign in1534_1 = {pp30[117]};
    assign in1534_2 = {pp31[116]};
    Full_Adder FA_1534(s1534, c1534, in1534_1, in1534_2, pp29[118]);
    wire[0:0] s1535, in1535_1, in1535_2;
    wire c1535;
    assign in1535_1 = {pp33[114]};
    assign in1535_2 = {pp34[113]};
    Full_Adder FA_1535(s1535, c1535, in1535_1, in1535_2, pp32[115]);
    wire[0:0] s1536, in1536_1, in1536_2;
    wire c1536;
    assign in1536_1 = {pp36[111]};
    assign in1536_2 = {pp37[110]};
    Full_Adder FA_1536(s1536, c1536, in1536_1, in1536_2, pp35[112]);
    wire[0:0] s1537, in1537_1, in1537_2;
    wire c1537;
    assign in1537_1 = {pp39[108]};
    assign in1537_2 = {pp40[107]};
    Full_Adder FA_1537(s1537, c1537, in1537_1, in1537_2, pp38[109]);
    wire[0:0] s1538, in1538_1, in1538_2;
    wire c1538;
    assign in1538_1 = {pp42[105]};
    assign in1538_2 = {pp43[104]};
    Full_Adder FA_1538(s1538, c1538, in1538_1, in1538_2, pp41[106]);
    wire[0:0] s1539, in1539_1, in1539_2;
    wire c1539;
    assign in1539_1 = {pp45[102]};
    assign in1539_2 = {pp46[101]};
    Full_Adder FA_1539(s1539, c1539, in1539_1, in1539_2, pp44[103]);
    wire[0:0] s1540, in1540_1, in1540_2;
    wire c1540;
    assign in1540_1 = {pp48[99]};
    assign in1540_2 = {pp49[98]};
    Full_Adder FA_1540(s1540, c1540, in1540_1, in1540_2, pp47[100]);
    wire[0:0] s1541, in1541_1, in1541_2;
    wire c1541;
    assign in1541_1 = {pp51[96]};
    assign in1541_2 = {pp52[95]};
    Full_Adder FA_1541(s1541, c1541, in1541_1, in1541_2, pp50[97]);
    wire[0:0] s1542, in1542_1, in1542_2;
    wire c1542;
    assign in1542_1 = {pp54[93]};
    assign in1542_2 = {pp55[92]};
    Full_Adder FA_1542(s1542, c1542, in1542_1, in1542_2, pp53[94]);
    wire[0:0] s1543, in1543_1, in1543_2;
    wire c1543;
    assign in1543_1 = {pp57[90]};
    assign in1543_2 = {pp58[89]};
    Full_Adder FA_1543(s1543, c1543, in1543_1, in1543_2, pp56[91]);
    wire[0:0] s1544, in1544_1, in1544_2;
    wire c1544;
    assign in1544_1 = {pp60[87]};
    assign in1544_2 = {pp61[86]};
    Full_Adder FA_1544(s1544, c1544, in1544_1, in1544_2, pp59[88]);
    wire[0:0] s1545, in1545_1, in1545_2;
    wire c1545;
    assign in1545_1 = {pp63[84]};
    assign in1545_2 = {pp64[83]};
    Full_Adder FA_1545(s1545, c1545, in1545_1, in1545_2, pp62[85]);
    wire[0:0] s1546, in1546_1, in1546_2;
    wire c1546;
    assign in1546_1 = {pp66[81]};
    assign in1546_2 = {pp67[80]};
    Full_Adder FA_1546(s1546, c1546, in1546_1, in1546_2, pp65[82]);
    wire[0:0] s1547, in1547_1, in1547_2;
    wire c1547;
    assign in1547_1 = {pp69[78]};
    assign in1547_2 = {pp70[77]};
    Full_Adder FA_1547(s1547, c1547, in1547_1, in1547_2, pp68[79]);
    wire[0:0] s1548, in1548_1, in1548_2;
    wire c1548;
    assign in1548_1 = {pp72[75]};
    assign in1548_2 = {pp73[74]};
    Full_Adder FA_1548(s1548, c1548, in1548_1, in1548_2, pp71[76]);
    wire[0:0] s1549, in1549_1, in1549_2;
    wire c1549;
    assign in1549_1 = {pp75[72]};
    assign in1549_2 = {pp76[71]};
    Full_Adder FA_1549(s1549, c1549, in1549_1, in1549_2, pp74[73]);
    wire[0:0] s1550, in1550_1, in1550_2;
    wire c1550;
    assign in1550_1 = {pp78[69]};
    assign in1550_2 = {pp79[68]};
    Full_Adder FA_1550(s1550, c1550, in1550_1, in1550_2, pp77[70]);
    wire[0:0] s1551, in1551_1, in1551_2;
    wire c1551;
    assign in1551_1 = {pp81[66]};
    assign in1551_2 = {pp82[65]};
    Full_Adder FA_1551(s1551, c1551, in1551_1, in1551_2, pp80[67]);
    wire[0:0] s1552, in1552_1, in1552_2;
    wire c1552;
    assign in1552_1 = {pp84[63]};
    assign in1552_2 = {pp85[62]};
    Full_Adder FA_1552(s1552, c1552, in1552_1, in1552_2, pp83[64]);
    wire[0:0] s1553, in1553_1, in1553_2;
    wire c1553;
    assign in1553_1 = {pp87[60]};
    assign in1553_2 = {pp88[59]};
    Full_Adder FA_1553(s1553, c1553, in1553_1, in1553_2, pp86[61]);
    wire[0:0] s1554, in1554_1, in1554_2;
    wire c1554;
    assign in1554_1 = {pp22[126]};
    assign in1554_2 = {pp23[125]};
    Full_Adder FA_1554(s1554, c1554, in1554_1, in1554_2, pp21[127]);
    wire[0:0] s1555, in1555_1, in1555_2;
    wire c1555;
    assign in1555_1 = {pp25[123]};
    assign in1555_2 = {pp26[122]};
    Full_Adder FA_1555(s1555, c1555, in1555_1, in1555_2, pp24[124]);
    wire[0:0] s1556, in1556_1, in1556_2;
    wire c1556;
    assign in1556_1 = {pp28[120]};
    assign in1556_2 = {pp29[119]};
    Full_Adder FA_1556(s1556, c1556, in1556_1, in1556_2, pp27[121]);
    wire[0:0] s1557, in1557_1, in1557_2;
    wire c1557;
    assign in1557_1 = {pp31[117]};
    assign in1557_2 = {pp32[116]};
    Full_Adder FA_1557(s1557, c1557, in1557_1, in1557_2, pp30[118]);
    wire[0:0] s1558, in1558_1, in1558_2;
    wire c1558;
    assign in1558_1 = {pp34[114]};
    assign in1558_2 = {pp35[113]};
    Full_Adder FA_1558(s1558, c1558, in1558_1, in1558_2, pp33[115]);
    wire[0:0] s1559, in1559_1, in1559_2;
    wire c1559;
    assign in1559_1 = {pp37[111]};
    assign in1559_2 = {pp38[110]};
    Full_Adder FA_1559(s1559, c1559, in1559_1, in1559_2, pp36[112]);
    wire[0:0] s1560, in1560_1, in1560_2;
    wire c1560;
    assign in1560_1 = {pp40[108]};
    assign in1560_2 = {pp41[107]};
    Full_Adder FA_1560(s1560, c1560, in1560_1, in1560_2, pp39[109]);
    wire[0:0] s1561, in1561_1, in1561_2;
    wire c1561;
    assign in1561_1 = {pp43[105]};
    assign in1561_2 = {pp44[104]};
    Full_Adder FA_1561(s1561, c1561, in1561_1, in1561_2, pp42[106]);
    wire[0:0] s1562, in1562_1, in1562_2;
    wire c1562;
    assign in1562_1 = {pp46[102]};
    assign in1562_2 = {pp47[101]};
    Full_Adder FA_1562(s1562, c1562, in1562_1, in1562_2, pp45[103]);
    wire[0:0] s1563, in1563_1, in1563_2;
    wire c1563;
    assign in1563_1 = {pp49[99]};
    assign in1563_2 = {pp50[98]};
    Full_Adder FA_1563(s1563, c1563, in1563_1, in1563_2, pp48[100]);
    wire[0:0] s1564, in1564_1, in1564_2;
    wire c1564;
    assign in1564_1 = {pp52[96]};
    assign in1564_2 = {pp53[95]};
    Full_Adder FA_1564(s1564, c1564, in1564_1, in1564_2, pp51[97]);
    wire[0:0] s1565, in1565_1, in1565_2;
    wire c1565;
    assign in1565_1 = {pp55[93]};
    assign in1565_2 = {pp56[92]};
    Full_Adder FA_1565(s1565, c1565, in1565_1, in1565_2, pp54[94]);
    wire[0:0] s1566, in1566_1, in1566_2;
    wire c1566;
    assign in1566_1 = {pp58[90]};
    assign in1566_2 = {pp59[89]};
    Full_Adder FA_1566(s1566, c1566, in1566_1, in1566_2, pp57[91]);
    wire[0:0] s1567, in1567_1, in1567_2;
    wire c1567;
    assign in1567_1 = {pp61[87]};
    assign in1567_2 = {pp62[86]};
    Full_Adder FA_1567(s1567, c1567, in1567_1, in1567_2, pp60[88]);
    wire[0:0] s1568, in1568_1, in1568_2;
    wire c1568;
    assign in1568_1 = {pp64[84]};
    assign in1568_2 = {pp65[83]};
    Full_Adder FA_1568(s1568, c1568, in1568_1, in1568_2, pp63[85]);
    wire[0:0] s1569, in1569_1, in1569_2;
    wire c1569;
    assign in1569_1 = {pp67[81]};
    assign in1569_2 = {pp68[80]};
    Full_Adder FA_1569(s1569, c1569, in1569_1, in1569_2, pp66[82]);
    wire[0:0] s1570, in1570_1, in1570_2;
    wire c1570;
    assign in1570_1 = {pp70[78]};
    assign in1570_2 = {pp71[77]};
    Full_Adder FA_1570(s1570, c1570, in1570_1, in1570_2, pp69[79]);
    wire[0:0] s1571, in1571_1, in1571_2;
    wire c1571;
    assign in1571_1 = {pp73[75]};
    assign in1571_2 = {pp74[74]};
    Full_Adder FA_1571(s1571, c1571, in1571_1, in1571_2, pp72[76]);
    wire[0:0] s1572, in1572_1, in1572_2;
    wire c1572;
    assign in1572_1 = {pp76[72]};
    assign in1572_2 = {pp77[71]};
    Full_Adder FA_1572(s1572, c1572, in1572_1, in1572_2, pp75[73]);
    wire[0:0] s1573, in1573_1, in1573_2;
    wire c1573;
    assign in1573_1 = {pp79[69]};
    assign in1573_2 = {pp80[68]};
    Full_Adder FA_1573(s1573, c1573, in1573_1, in1573_2, pp78[70]);
    wire[0:0] s1574, in1574_1, in1574_2;
    wire c1574;
    assign in1574_1 = {pp82[66]};
    assign in1574_2 = {pp83[65]};
    Full_Adder FA_1574(s1574, c1574, in1574_1, in1574_2, pp81[67]);
    wire[0:0] s1575, in1575_1, in1575_2;
    wire c1575;
    assign in1575_1 = {pp85[63]};
    assign in1575_2 = {pp86[62]};
    Full_Adder FA_1575(s1575, c1575, in1575_1, in1575_2, pp84[64]);
    wire[0:0] s1576, in1576_1, in1576_2;
    wire c1576;
    assign in1576_1 = {pp23[126]};
    assign in1576_2 = {pp24[125]};
    Full_Adder FA_1576(s1576, c1576, in1576_1, in1576_2, pp22[127]);
    wire[0:0] s1577, in1577_1, in1577_2;
    wire c1577;
    assign in1577_1 = {pp26[123]};
    assign in1577_2 = {pp27[122]};
    Full_Adder FA_1577(s1577, c1577, in1577_1, in1577_2, pp25[124]);
    wire[0:0] s1578, in1578_1, in1578_2;
    wire c1578;
    assign in1578_1 = {pp29[120]};
    assign in1578_2 = {pp30[119]};
    Full_Adder FA_1578(s1578, c1578, in1578_1, in1578_2, pp28[121]);
    wire[0:0] s1579, in1579_1, in1579_2;
    wire c1579;
    assign in1579_1 = {pp32[117]};
    assign in1579_2 = {pp33[116]};
    Full_Adder FA_1579(s1579, c1579, in1579_1, in1579_2, pp31[118]);
    wire[0:0] s1580, in1580_1, in1580_2;
    wire c1580;
    assign in1580_1 = {pp35[114]};
    assign in1580_2 = {pp36[113]};
    Full_Adder FA_1580(s1580, c1580, in1580_1, in1580_2, pp34[115]);
    wire[0:0] s1581, in1581_1, in1581_2;
    wire c1581;
    assign in1581_1 = {pp38[111]};
    assign in1581_2 = {pp39[110]};
    Full_Adder FA_1581(s1581, c1581, in1581_1, in1581_2, pp37[112]);
    wire[0:0] s1582, in1582_1, in1582_2;
    wire c1582;
    assign in1582_1 = {pp41[108]};
    assign in1582_2 = {pp42[107]};
    Full_Adder FA_1582(s1582, c1582, in1582_1, in1582_2, pp40[109]);
    wire[0:0] s1583, in1583_1, in1583_2;
    wire c1583;
    assign in1583_1 = {pp44[105]};
    assign in1583_2 = {pp45[104]};
    Full_Adder FA_1583(s1583, c1583, in1583_1, in1583_2, pp43[106]);
    wire[0:0] s1584, in1584_1, in1584_2;
    wire c1584;
    assign in1584_1 = {pp47[102]};
    assign in1584_2 = {pp48[101]};
    Full_Adder FA_1584(s1584, c1584, in1584_1, in1584_2, pp46[103]);
    wire[0:0] s1585, in1585_1, in1585_2;
    wire c1585;
    assign in1585_1 = {pp50[99]};
    assign in1585_2 = {pp51[98]};
    Full_Adder FA_1585(s1585, c1585, in1585_1, in1585_2, pp49[100]);
    wire[0:0] s1586, in1586_1, in1586_2;
    wire c1586;
    assign in1586_1 = {pp53[96]};
    assign in1586_2 = {pp54[95]};
    Full_Adder FA_1586(s1586, c1586, in1586_1, in1586_2, pp52[97]);
    wire[0:0] s1587, in1587_1, in1587_2;
    wire c1587;
    assign in1587_1 = {pp56[93]};
    assign in1587_2 = {pp57[92]};
    Full_Adder FA_1587(s1587, c1587, in1587_1, in1587_2, pp55[94]);
    wire[0:0] s1588, in1588_1, in1588_2;
    wire c1588;
    assign in1588_1 = {pp59[90]};
    assign in1588_2 = {pp60[89]};
    Full_Adder FA_1588(s1588, c1588, in1588_1, in1588_2, pp58[91]);
    wire[0:0] s1589, in1589_1, in1589_2;
    wire c1589;
    assign in1589_1 = {pp62[87]};
    assign in1589_2 = {pp63[86]};
    Full_Adder FA_1589(s1589, c1589, in1589_1, in1589_2, pp61[88]);
    wire[0:0] s1590, in1590_1, in1590_2;
    wire c1590;
    assign in1590_1 = {pp65[84]};
    assign in1590_2 = {pp66[83]};
    Full_Adder FA_1590(s1590, c1590, in1590_1, in1590_2, pp64[85]);
    wire[0:0] s1591, in1591_1, in1591_2;
    wire c1591;
    assign in1591_1 = {pp68[81]};
    assign in1591_2 = {pp69[80]};
    Full_Adder FA_1591(s1591, c1591, in1591_1, in1591_2, pp67[82]);
    wire[0:0] s1592, in1592_1, in1592_2;
    wire c1592;
    assign in1592_1 = {pp71[78]};
    assign in1592_2 = {pp72[77]};
    Full_Adder FA_1592(s1592, c1592, in1592_1, in1592_2, pp70[79]);
    wire[0:0] s1593, in1593_1, in1593_2;
    wire c1593;
    assign in1593_1 = {pp74[75]};
    assign in1593_2 = {pp75[74]};
    Full_Adder FA_1593(s1593, c1593, in1593_1, in1593_2, pp73[76]);
    wire[0:0] s1594, in1594_1, in1594_2;
    wire c1594;
    assign in1594_1 = {pp77[72]};
    assign in1594_2 = {pp78[71]};
    Full_Adder FA_1594(s1594, c1594, in1594_1, in1594_2, pp76[73]);
    wire[0:0] s1595, in1595_1, in1595_2;
    wire c1595;
    assign in1595_1 = {pp80[69]};
    assign in1595_2 = {pp81[68]};
    Full_Adder FA_1595(s1595, c1595, in1595_1, in1595_2, pp79[70]);
    wire[0:0] s1596, in1596_1, in1596_2;
    wire c1596;
    assign in1596_1 = {pp83[66]};
    assign in1596_2 = {pp84[65]};
    Full_Adder FA_1596(s1596, c1596, in1596_1, in1596_2, pp82[67]);
    wire[0:0] s1597, in1597_1, in1597_2;
    wire c1597;
    assign in1597_1 = {pp24[126]};
    assign in1597_2 = {pp25[125]};
    Full_Adder FA_1597(s1597, c1597, in1597_1, in1597_2, pp23[127]);
    wire[0:0] s1598, in1598_1, in1598_2;
    wire c1598;
    assign in1598_1 = {pp27[123]};
    assign in1598_2 = {pp28[122]};
    Full_Adder FA_1598(s1598, c1598, in1598_1, in1598_2, pp26[124]);
    wire[0:0] s1599, in1599_1, in1599_2;
    wire c1599;
    assign in1599_1 = {pp30[120]};
    assign in1599_2 = {pp31[119]};
    Full_Adder FA_1599(s1599, c1599, in1599_1, in1599_2, pp29[121]);
    wire[0:0] s1600, in1600_1, in1600_2;
    wire c1600;
    assign in1600_1 = {pp33[117]};
    assign in1600_2 = {pp34[116]};
    Full_Adder FA_1600(s1600, c1600, in1600_1, in1600_2, pp32[118]);
    wire[0:0] s1601, in1601_1, in1601_2;
    wire c1601;
    assign in1601_1 = {pp36[114]};
    assign in1601_2 = {pp37[113]};
    Full_Adder FA_1601(s1601, c1601, in1601_1, in1601_2, pp35[115]);
    wire[0:0] s1602, in1602_1, in1602_2;
    wire c1602;
    assign in1602_1 = {pp39[111]};
    assign in1602_2 = {pp40[110]};
    Full_Adder FA_1602(s1602, c1602, in1602_1, in1602_2, pp38[112]);
    wire[0:0] s1603, in1603_1, in1603_2;
    wire c1603;
    assign in1603_1 = {pp42[108]};
    assign in1603_2 = {pp43[107]};
    Full_Adder FA_1603(s1603, c1603, in1603_1, in1603_2, pp41[109]);
    wire[0:0] s1604, in1604_1, in1604_2;
    wire c1604;
    assign in1604_1 = {pp45[105]};
    assign in1604_2 = {pp46[104]};
    Full_Adder FA_1604(s1604, c1604, in1604_1, in1604_2, pp44[106]);
    wire[0:0] s1605, in1605_1, in1605_2;
    wire c1605;
    assign in1605_1 = {pp48[102]};
    assign in1605_2 = {pp49[101]};
    Full_Adder FA_1605(s1605, c1605, in1605_1, in1605_2, pp47[103]);
    wire[0:0] s1606, in1606_1, in1606_2;
    wire c1606;
    assign in1606_1 = {pp51[99]};
    assign in1606_2 = {pp52[98]};
    Full_Adder FA_1606(s1606, c1606, in1606_1, in1606_2, pp50[100]);
    wire[0:0] s1607, in1607_1, in1607_2;
    wire c1607;
    assign in1607_1 = {pp54[96]};
    assign in1607_2 = {pp55[95]};
    Full_Adder FA_1607(s1607, c1607, in1607_1, in1607_2, pp53[97]);
    wire[0:0] s1608, in1608_1, in1608_2;
    wire c1608;
    assign in1608_1 = {pp57[93]};
    assign in1608_2 = {pp58[92]};
    Full_Adder FA_1608(s1608, c1608, in1608_1, in1608_2, pp56[94]);
    wire[0:0] s1609, in1609_1, in1609_2;
    wire c1609;
    assign in1609_1 = {pp60[90]};
    assign in1609_2 = {pp61[89]};
    Full_Adder FA_1609(s1609, c1609, in1609_1, in1609_2, pp59[91]);
    wire[0:0] s1610, in1610_1, in1610_2;
    wire c1610;
    assign in1610_1 = {pp63[87]};
    assign in1610_2 = {pp64[86]};
    Full_Adder FA_1610(s1610, c1610, in1610_1, in1610_2, pp62[88]);
    wire[0:0] s1611, in1611_1, in1611_2;
    wire c1611;
    assign in1611_1 = {pp66[84]};
    assign in1611_2 = {pp67[83]};
    Full_Adder FA_1611(s1611, c1611, in1611_1, in1611_2, pp65[85]);
    wire[0:0] s1612, in1612_1, in1612_2;
    wire c1612;
    assign in1612_1 = {pp69[81]};
    assign in1612_2 = {pp70[80]};
    Full_Adder FA_1612(s1612, c1612, in1612_1, in1612_2, pp68[82]);
    wire[0:0] s1613, in1613_1, in1613_2;
    wire c1613;
    assign in1613_1 = {pp72[78]};
    assign in1613_2 = {pp73[77]};
    Full_Adder FA_1613(s1613, c1613, in1613_1, in1613_2, pp71[79]);
    wire[0:0] s1614, in1614_1, in1614_2;
    wire c1614;
    assign in1614_1 = {pp75[75]};
    assign in1614_2 = {pp76[74]};
    Full_Adder FA_1614(s1614, c1614, in1614_1, in1614_2, pp74[76]);
    wire[0:0] s1615, in1615_1, in1615_2;
    wire c1615;
    assign in1615_1 = {pp78[72]};
    assign in1615_2 = {pp79[71]};
    Full_Adder FA_1615(s1615, c1615, in1615_1, in1615_2, pp77[73]);
    wire[0:0] s1616, in1616_1, in1616_2;
    wire c1616;
    assign in1616_1 = {pp81[69]};
    assign in1616_2 = {pp82[68]};
    Full_Adder FA_1616(s1616, c1616, in1616_1, in1616_2, pp80[70]);
    wire[0:0] s1617, in1617_1, in1617_2;
    wire c1617;
    assign in1617_1 = {pp25[126]};
    assign in1617_2 = {pp26[125]};
    Full_Adder FA_1617(s1617, c1617, in1617_1, in1617_2, pp24[127]);
    wire[0:0] s1618, in1618_1, in1618_2;
    wire c1618;
    assign in1618_1 = {pp28[123]};
    assign in1618_2 = {pp29[122]};
    Full_Adder FA_1618(s1618, c1618, in1618_1, in1618_2, pp27[124]);
    wire[0:0] s1619, in1619_1, in1619_2;
    wire c1619;
    assign in1619_1 = {pp31[120]};
    assign in1619_2 = {pp32[119]};
    Full_Adder FA_1619(s1619, c1619, in1619_1, in1619_2, pp30[121]);
    wire[0:0] s1620, in1620_1, in1620_2;
    wire c1620;
    assign in1620_1 = {pp34[117]};
    assign in1620_2 = {pp35[116]};
    Full_Adder FA_1620(s1620, c1620, in1620_1, in1620_2, pp33[118]);
    wire[0:0] s1621, in1621_1, in1621_2;
    wire c1621;
    assign in1621_1 = {pp37[114]};
    assign in1621_2 = {pp38[113]};
    Full_Adder FA_1621(s1621, c1621, in1621_1, in1621_2, pp36[115]);
    wire[0:0] s1622, in1622_1, in1622_2;
    wire c1622;
    assign in1622_1 = {pp40[111]};
    assign in1622_2 = {pp41[110]};
    Full_Adder FA_1622(s1622, c1622, in1622_1, in1622_2, pp39[112]);
    wire[0:0] s1623, in1623_1, in1623_2;
    wire c1623;
    assign in1623_1 = {pp43[108]};
    assign in1623_2 = {pp44[107]};
    Full_Adder FA_1623(s1623, c1623, in1623_1, in1623_2, pp42[109]);
    wire[0:0] s1624, in1624_1, in1624_2;
    wire c1624;
    assign in1624_1 = {pp46[105]};
    assign in1624_2 = {pp47[104]};
    Full_Adder FA_1624(s1624, c1624, in1624_1, in1624_2, pp45[106]);
    wire[0:0] s1625, in1625_1, in1625_2;
    wire c1625;
    assign in1625_1 = {pp49[102]};
    assign in1625_2 = {pp50[101]};
    Full_Adder FA_1625(s1625, c1625, in1625_1, in1625_2, pp48[103]);
    wire[0:0] s1626, in1626_1, in1626_2;
    wire c1626;
    assign in1626_1 = {pp52[99]};
    assign in1626_2 = {pp53[98]};
    Full_Adder FA_1626(s1626, c1626, in1626_1, in1626_2, pp51[100]);
    wire[0:0] s1627, in1627_1, in1627_2;
    wire c1627;
    assign in1627_1 = {pp55[96]};
    assign in1627_2 = {pp56[95]};
    Full_Adder FA_1627(s1627, c1627, in1627_1, in1627_2, pp54[97]);
    wire[0:0] s1628, in1628_1, in1628_2;
    wire c1628;
    assign in1628_1 = {pp58[93]};
    assign in1628_2 = {pp59[92]};
    Full_Adder FA_1628(s1628, c1628, in1628_1, in1628_2, pp57[94]);
    wire[0:0] s1629, in1629_1, in1629_2;
    wire c1629;
    assign in1629_1 = {pp61[90]};
    assign in1629_2 = {pp62[89]};
    Full_Adder FA_1629(s1629, c1629, in1629_1, in1629_2, pp60[91]);
    wire[0:0] s1630, in1630_1, in1630_2;
    wire c1630;
    assign in1630_1 = {pp64[87]};
    assign in1630_2 = {pp65[86]};
    Full_Adder FA_1630(s1630, c1630, in1630_1, in1630_2, pp63[88]);
    wire[0:0] s1631, in1631_1, in1631_2;
    wire c1631;
    assign in1631_1 = {pp67[84]};
    assign in1631_2 = {pp68[83]};
    Full_Adder FA_1631(s1631, c1631, in1631_1, in1631_2, pp66[85]);
    wire[0:0] s1632, in1632_1, in1632_2;
    wire c1632;
    assign in1632_1 = {pp70[81]};
    assign in1632_2 = {pp71[80]};
    Full_Adder FA_1632(s1632, c1632, in1632_1, in1632_2, pp69[82]);
    wire[0:0] s1633, in1633_1, in1633_2;
    wire c1633;
    assign in1633_1 = {pp73[78]};
    assign in1633_2 = {pp74[77]};
    Full_Adder FA_1633(s1633, c1633, in1633_1, in1633_2, pp72[79]);
    wire[0:0] s1634, in1634_1, in1634_2;
    wire c1634;
    assign in1634_1 = {pp76[75]};
    assign in1634_2 = {pp77[74]};
    Full_Adder FA_1634(s1634, c1634, in1634_1, in1634_2, pp75[76]);
    wire[0:0] s1635, in1635_1, in1635_2;
    wire c1635;
    assign in1635_1 = {pp79[72]};
    assign in1635_2 = {pp80[71]};
    Full_Adder FA_1635(s1635, c1635, in1635_1, in1635_2, pp78[73]);
    wire[0:0] s1636, in1636_1, in1636_2;
    wire c1636;
    assign in1636_1 = {pp26[126]};
    assign in1636_2 = {pp27[125]};
    Full_Adder FA_1636(s1636, c1636, in1636_1, in1636_2, pp25[127]);
    wire[0:0] s1637, in1637_1, in1637_2;
    wire c1637;
    assign in1637_1 = {pp29[123]};
    assign in1637_2 = {pp30[122]};
    Full_Adder FA_1637(s1637, c1637, in1637_1, in1637_2, pp28[124]);
    wire[0:0] s1638, in1638_1, in1638_2;
    wire c1638;
    assign in1638_1 = {pp32[120]};
    assign in1638_2 = {pp33[119]};
    Full_Adder FA_1638(s1638, c1638, in1638_1, in1638_2, pp31[121]);
    wire[0:0] s1639, in1639_1, in1639_2;
    wire c1639;
    assign in1639_1 = {pp35[117]};
    assign in1639_2 = {pp36[116]};
    Full_Adder FA_1639(s1639, c1639, in1639_1, in1639_2, pp34[118]);
    wire[0:0] s1640, in1640_1, in1640_2;
    wire c1640;
    assign in1640_1 = {pp38[114]};
    assign in1640_2 = {pp39[113]};
    Full_Adder FA_1640(s1640, c1640, in1640_1, in1640_2, pp37[115]);
    wire[0:0] s1641, in1641_1, in1641_2;
    wire c1641;
    assign in1641_1 = {pp41[111]};
    assign in1641_2 = {pp42[110]};
    Full_Adder FA_1641(s1641, c1641, in1641_1, in1641_2, pp40[112]);
    wire[0:0] s1642, in1642_1, in1642_2;
    wire c1642;
    assign in1642_1 = {pp44[108]};
    assign in1642_2 = {pp45[107]};
    Full_Adder FA_1642(s1642, c1642, in1642_1, in1642_2, pp43[109]);
    wire[0:0] s1643, in1643_1, in1643_2;
    wire c1643;
    assign in1643_1 = {pp47[105]};
    assign in1643_2 = {pp48[104]};
    Full_Adder FA_1643(s1643, c1643, in1643_1, in1643_2, pp46[106]);
    wire[0:0] s1644, in1644_1, in1644_2;
    wire c1644;
    assign in1644_1 = {pp50[102]};
    assign in1644_2 = {pp51[101]};
    Full_Adder FA_1644(s1644, c1644, in1644_1, in1644_2, pp49[103]);
    wire[0:0] s1645, in1645_1, in1645_2;
    wire c1645;
    assign in1645_1 = {pp53[99]};
    assign in1645_2 = {pp54[98]};
    Full_Adder FA_1645(s1645, c1645, in1645_1, in1645_2, pp52[100]);
    wire[0:0] s1646, in1646_1, in1646_2;
    wire c1646;
    assign in1646_1 = {pp56[96]};
    assign in1646_2 = {pp57[95]};
    Full_Adder FA_1646(s1646, c1646, in1646_1, in1646_2, pp55[97]);
    wire[0:0] s1647, in1647_1, in1647_2;
    wire c1647;
    assign in1647_1 = {pp59[93]};
    assign in1647_2 = {pp60[92]};
    Full_Adder FA_1647(s1647, c1647, in1647_1, in1647_2, pp58[94]);
    wire[0:0] s1648, in1648_1, in1648_2;
    wire c1648;
    assign in1648_1 = {pp62[90]};
    assign in1648_2 = {pp63[89]};
    Full_Adder FA_1648(s1648, c1648, in1648_1, in1648_2, pp61[91]);
    wire[0:0] s1649, in1649_1, in1649_2;
    wire c1649;
    assign in1649_1 = {pp65[87]};
    assign in1649_2 = {pp66[86]};
    Full_Adder FA_1649(s1649, c1649, in1649_1, in1649_2, pp64[88]);
    wire[0:0] s1650, in1650_1, in1650_2;
    wire c1650;
    assign in1650_1 = {pp68[84]};
    assign in1650_2 = {pp69[83]};
    Full_Adder FA_1650(s1650, c1650, in1650_1, in1650_2, pp67[85]);
    wire[0:0] s1651, in1651_1, in1651_2;
    wire c1651;
    assign in1651_1 = {pp71[81]};
    assign in1651_2 = {pp72[80]};
    Full_Adder FA_1651(s1651, c1651, in1651_1, in1651_2, pp70[82]);
    wire[0:0] s1652, in1652_1, in1652_2;
    wire c1652;
    assign in1652_1 = {pp74[78]};
    assign in1652_2 = {pp75[77]};
    Full_Adder FA_1652(s1652, c1652, in1652_1, in1652_2, pp73[79]);
    wire[0:0] s1653, in1653_1, in1653_2;
    wire c1653;
    assign in1653_1 = {pp77[75]};
    assign in1653_2 = {pp78[74]};
    Full_Adder FA_1653(s1653, c1653, in1653_1, in1653_2, pp76[76]);
    wire[0:0] s1654, in1654_1, in1654_2;
    wire c1654;
    assign in1654_1 = {pp27[126]};
    assign in1654_2 = {pp28[125]};
    Full_Adder FA_1654(s1654, c1654, in1654_1, in1654_2, pp26[127]);
    wire[0:0] s1655, in1655_1, in1655_2;
    wire c1655;
    assign in1655_1 = {pp30[123]};
    assign in1655_2 = {pp31[122]};
    Full_Adder FA_1655(s1655, c1655, in1655_1, in1655_2, pp29[124]);
    wire[0:0] s1656, in1656_1, in1656_2;
    wire c1656;
    assign in1656_1 = {pp33[120]};
    assign in1656_2 = {pp34[119]};
    Full_Adder FA_1656(s1656, c1656, in1656_1, in1656_2, pp32[121]);
    wire[0:0] s1657, in1657_1, in1657_2;
    wire c1657;
    assign in1657_1 = {pp36[117]};
    assign in1657_2 = {pp37[116]};
    Full_Adder FA_1657(s1657, c1657, in1657_1, in1657_2, pp35[118]);
    wire[0:0] s1658, in1658_1, in1658_2;
    wire c1658;
    assign in1658_1 = {pp39[114]};
    assign in1658_2 = {pp40[113]};
    Full_Adder FA_1658(s1658, c1658, in1658_1, in1658_2, pp38[115]);
    wire[0:0] s1659, in1659_1, in1659_2;
    wire c1659;
    assign in1659_1 = {pp42[111]};
    assign in1659_2 = {pp43[110]};
    Full_Adder FA_1659(s1659, c1659, in1659_1, in1659_2, pp41[112]);
    wire[0:0] s1660, in1660_1, in1660_2;
    wire c1660;
    assign in1660_1 = {pp45[108]};
    assign in1660_2 = {pp46[107]};
    Full_Adder FA_1660(s1660, c1660, in1660_1, in1660_2, pp44[109]);
    wire[0:0] s1661, in1661_1, in1661_2;
    wire c1661;
    assign in1661_1 = {pp48[105]};
    assign in1661_2 = {pp49[104]};
    Full_Adder FA_1661(s1661, c1661, in1661_1, in1661_2, pp47[106]);
    wire[0:0] s1662, in1662_1, in1662_2;
    wire c1662;
    assign in1662_1 = {pp51[102]};
    assign in1662_2 = {pp52[101]};
    Full_Adder FA_1662(s1662, c1662, in1662_1, in1662_2, pp50[103]);
    wire[0:0] s1663, in1663_1, in1663_2;
    wire c1663;
    assign in1663_1 = {pp54[99]};
    assign in1663_2 = {pp55[98]};
    Full_Adder FA_1663(s1663, c1663, in1663_1, in1663_2, pp53[100]);
    wire[0:0] s1664, in1664_1, in1664_2;
    wire c1664;
    assign in1664_1 = {pp57[96]};
    assign in1664_2 = {pp58[95]};
    Full_Adder FA_1664(s1664, c1664, in1664_1, in1664_2, pp56[97]);
    wire[0:0] s1665, in1665_1, in1665_2;
    wire c1665;
    assign in1665_1 = {pp60[93]};
    assign in1665_2 = {pp61[92]};
    Full_Adder FA_1665(s1665, c1665, in1665_1, in1665_2, pp59[94]);
    wire[0:0] s1666, in1666_1, in1666_2;
    wire c1666;
    assign in1666_1 = {pp63[90]};
    assign in1666_2 = {pp64[89]};
    Full_Adder FA_1666(s1666, c1666, in1666_1, in1666_2, pp62[91]);
    wire[0:0] s1667, in1667_1, in1667_2;
    wire c1667;
    assign in1667_1 = {pp66[87]};
    assign in1667_2 = {pp67[86]};
    Full_Adder FA_1667(s1667, c1667, in1667_1, in1667_2, pp65[88]);
    wire[0:0] s1668, in1668_1, in1668_2;
    wire c1668;
    assign in1668_1 = {pp69[84]};
    assign in1668_2 = {pp70[83]};
    Full_Adder FA_1668(s1668, c1668, in1668_1, in1668_2, pp68[85]);
    wire[0:0] s1669, in1669_1, in1669_2;
    wire c1669;
    assign in1669_1 = {pp72[81]};
    assign in1669_2 = {pp73[80]};
    Full_Adder FA_1669(s1669, c1669, in1669_1, in1669_2, pp71[82]);
    wire[0:0] s1670, in1670_1, in1670_2;
    wire c1670;
    assign in1670_1 = {pp75[78]};
    assign in1670_2 = {pp76[77]};
    Full_Adder FA_1670(s1670, c1670, in1670_1, in1670_2, pp74[79]);
    wire[0:0] s1671, in1671_1, in1671_2;
    wire c1671;
    assign in1671_1 = {pp28[126]};
    assign in1671_2 = {pp29[125]};
    Full_Adder FA_1671(s1671, c1671, in1671_1, in1671_2, pp27[127]);
    wire[0:0] s1672, in1672_1, in1672_2;
    wire c1672;
    assign in1672_1 = {pp31[123]};
    assign in1672_2 = {pp32[122]};
    Full_Adder FA_1672(s1672, c1672, in1672_1, in1672_2, pp30[124]);
    wire[0:0] s1673, in1673_1, in1673_2;
    wire c1673;
    assign in1673_1 = {pp34[120]};
    assign in1673_2 = {pp35[119]};
    Full_Adder FA_1673(s1673, c1673, in1673_1, in1673_2, pp33[121]);
    wire[0:0] s1674, in1674_1, in1674_2;
    wire c1674;
    assign in1674_1 = {pp37[117]};
    assign in1674_2 = {pp38[116]};
    Full_Adder FA_1674(s1674, c1674, in1674_1, in1674_2, pp36[118]);
    wire[0:0] s1675, in1675_1, in1675_2;
    wire c1675;
    assign in1675_1 = {pp40[114]};
    assign in1675_2 = {pp41[113]};
    Full_Adder FA_1675(s1675, c1675, in1675_1, in1675_2, pp39[115]);
    wire[0:0] s1676, in1676_1, in1676_2;
    wire c1676;
    assign in1676_1 = {pp43[111]};
    assign in1676_2 = {pp44[110]};
    Full_Adder FA_1676(s1676, c1676, in1676_1, in1676_2, pp42[112]);
    wire[0:0] s1677, in1677_1, in1677_2;
    wire c1677;
    assign in1677_1 = {pp46[108]};
    assign in1677_2 = {pp47[107]};
    Full_Adder FA_1677(s1677, c1677, in1677_1, in1677_2, pp45[109]);
    wire[0:0] s1678, in1678_1, in1678_2;
    wire c1678;
    assign in1678_1 = {pp49[105]};
    assign in1678_2 = {pp50[104]};
    Full_Adder FA_1678(s1678, c1678, in1678_1, in1678_2, pp48[106]);
    wire[0:0] s1679, in1679_1, in1679_2;
    wire c1679;
    assign in1679_1 = {pp52[102]};
    assign in1679_2 = {pp53[101]};
    Full_Adder FA_1679(s1679, c1679, in1679_1, in1679_2, pp51[103]);
    wire[0:0] s1680, in1680_1, in1680_2;
    wire c1680;
    assign in1680_1 = {pp55[99]};
    assign in1680_2 = {pp56[98]};
    Full_Adder FA_1680(s1680, c1680, in1680_1, in1680_2, pp54[100]);
    wire[0:0] s1681, in1681_1, in1681_2;
    wire c1681;
    assign in1681_1 = {pp58[96]};
    assign in1681_2 = {pp59[95]};
    Full_Adder FA_1681(s1681, c1681, in1681_1, in1681_2, pp57[97]);
    wire[0:0] s1682, in1682_1, in1682_2;
    wire c1682;
    assign in1682_1 = {pp61[93]};
    assign in1682_2 = {pp62[92]};
    Full_Adder FA_1682(s1682, c1682, in1682_1, in1682_2, pp60[94]);
    wire[0:0] s1683, in1683_1, in1683_2;
    wire c1683;
    assign in1683_1 = {pp64[90]};
    assign in1683_2 = {pp65[89]};
    Full_Adder FA_1683(s1683, c1683, in1683_1, in1683_2, pp63[91]);
    wire[0:0] s1684, in1684_1, in1684_2;
    wire c1684;
    assign in1684_1 = {pp67[87]};
    assign in1684_2 = {pp68[86]};
    Full_Adder FA_1684(s1684, c1684, in1684_1, in1684_2, pp66[88]);
    wire[0:0] s1685, in1685_1, in1685_2;
    wire c1685;
    assign in1685_1 = {pp70[84]};
    assign in1685_2 = {pp71[83]};
    Full_Adder FA_1685(s1685, c1685, in1685_1, in1685_2, pp69[85]);
    wire[0:0] s1686, in1686_1, in1686_2;
    wire c1686;
    assign in1686_1 = {pp73[81]};
    assign in1686_2 = {pp74[80]};
    Full_Adder FA_1686(s1686, c1686, in1686_1, in1686_2, pp72[82]);
    wire[0:0] s1687, in1687_1, in1687_2;
    wire c1687;
    assign in1687_1 = {pp29[126]};
    assign in1687_2 = {pp30[125]};
    Full_Adder FA_1687(s1687, c1687, in1687_1, in1687_2, pp28[127]);
    wire[0:0] s1688, in1688_1, in1688_2;
    wire c1688;
    assign in1688_1 = {pp32[123]};
    assign in1688_2 = {pp33[122]};
    Full_Adder FA_1688(s1688, c1688, in1688_1, in1688_2, pp31[124]);
    wire[0:0] s1689, in1689_1, in1689_2;
    wire c1689;
    assign in1689_1 = {pp35[120]};
    assign in1689_2 = {pp36[119]};
    Full_Adder FA_1689(s1689, c1689, in1689_1, in1689_2, pp34[121]);
    wire[0:0] s1690, in1690_1, in1690_2;
    wire c1690;
    assign in1690_1 = {pp38[117]};
    assign in1690_2 = {pp39[116]};
    Full_Adder FA_1690(s1690, c1690, in1690_1, in1690_2, pp37[118]);
    wire[0:0] s1691, in1691_1, in1691_2;
    wire c1691;
    assign in1691_1 = {pp41[114]};
    assign in1691_2 = {pp42[113]};
    Full_Adder FA_1691(s1691, c1691, in1691_1, in1691_2, pp40[115]);
    wire[0:0] s1692, in1692_1, in1692_2;
    wire c1692;
    assign in1692_1 = {pp44[111]};
    assign in1692_2 = {pp45[110]};
    Full_Adder FA_1692(s1692, c1692, in1692_1, in1692_2, pp43[112]);
    wire[0:0] s1693, in1693_1, in1693_2;
    wire c1693;
    assign in1693_1 = {pp47[108]};
    assign in1693_2 = {pp48[107]};
    Full_Adder FA_1693(s1693, c1693, in1693_1, in1693_2, pp46[109]);
    wire[0:0] s1694, in1694_1, in1694_2;
    wire c1694;
    assign in1694_1 = {pp50[105]};
    assign in1694_2 = {pp51[104]};
    Full_Adder FA_1694(s1694, c1694, in1694_1, in1694_2, pp49[106]);
    wire[0:0] s1695, in1695_1, in1695_2;
    wire c1695;
    assign in1695_1 = {pp53[102]};
    assign in1695_2 = {pp54[101]};
    Full_Adder FA_1695(s1695, c1695, in1695_1, in1695_2, pp52[103]);
    wire[0:0] s1696, in1696_1, in1696_2;
    wire c1696;
    assign in1696_1 = {pp56[99]};
    assign in1696_2 = {pp57[98]};
    Full_Adder FA_1696(s1696, c1696, in1696_1, in1696_2, pp55[100]);
    wire[0:0] s1697, in1697_1, in1697_2;
    wire c1697;
    assign in1697_1 = {pp59[96]};
    assign in1697_2 = {pp60[95]};
    Full_Adder FA_1697(s1697, c1697, in1697_1, in1697_2, pp58[97]);
    wire[0:0] s1698, in1698_1, in1698_2;
    wire c1698;
    assign in1698_1 = {pp62[93]};
    assign in1698_2 = {pp63[92]};
    Full_Adder FA_1698(s1698, c1698, in1698_1, in1698_2, pp61[94]);
    wire[0:0] s1699, in1699_1, in1699_2;
    wire c1699;
    assign in1699_1 = {pp65[90]};
    assign in1699_2 = {pp66[89]};
    Full_Adder FA_1699(s1699, c1699, in1699_1, in1699_2, pp64[91]);
    wire[0:0] s1700, in1700_1, in1700_2;
    wire c1700;
    assign in1700_1 = {pp68[87]};
    assign in1700_2 = {pp69[86]};
    Full_Adder FA_1700(s1700, c1700, in1700_1, in1700_2, pp67[88]);
    wire[0:0] s1701, in1701_1, in1701_2;
    wire c1701;
    assign in1701_1 = {pp71[84]};
    assign in1701_2 = {pp72[83]};
    Full_Adder FA_1701(s1701, c1701, in1701_1, in1701_2, pp70[85]);
    wire[0:0] s1702, in1702_1, in1702_2;
    wire c1702;
    assign in1702_1 = {pp30[126]};
    assign in1702_2 = {pp31[125]};
    Full_Adder FA_1702(s1702, c1702, in1702_1, in1702_2, pp29[127]);
    wire[0:0] s1703, in1703_1, in1703_2;
    wire c1703;
    assign in1703_1 = {pp33[123]};
    assign in1703_2 = {pp34[122]};
    Full_Adder FA_1703(s1703, c1703, in1703_1, in1703_2, pp32[124]);
    wire[0:0] s1704, in1704_1, in1704_2;
    wire c1704;
    assign in1704_1 = {pp36[120]};
    assign in1704_2 = {pp37[119]};
    Full_Adder FA_1704(s1704, c1704, in1704_1, in1704_2, pp35[121]);
    wire[0:0] s1705, in1705_1, in1705_2;
    wire c1705;
    assign in1705_1 = {pp39[117]};
    assign in1705_2 = {pp40[116]};
    Full_Adder FA_1705(s1705, c1705, in1705_1, in1705_2, pp38[118]);
    wire[0:0] s1706, in1706_1, in1706_2;
    wire c1706;
    assign in1706_1 = {pp42[114]};
    assign in1706_2 = {pp43[113]};
    Full_Adder FA_1706(s1706, c1706, in1706_1, in1706_2, pp41[115]);
    wire[0:0] s1707, in1707_1, in1707_2;
    wire c1707;
    assign in1707_1 = {pp45[111]};
    assign in1707_2 = {pp46[110]};
    Full_Adder FA_1707(s1707, c1707, in1707_1, in1707_2, pp44[112]);
    wire[0:0] s1708, in1708_1, in1708_2;
    wire c1708;
    assign in1708_1 = {pp48[108]};
    assign in1708_2 = {pp49[107]};
    Full_Adder FA_1708(s1708, c1708, in1708_1, in1708_2, pp47[109]);
    wire[0:0] s1709, in1709_1, in1709_2;
    wire c1709;
    assign in1709_1 = {pp51[105]};
    assign in1709_2 = {pp52[104]};
    Full_Adder FA_1709(s1709, c1709, in1709_1, in1709_2, pp50[106]);
    wire[0:0] s1710, in1710_1, in1710_2;
    wire c1710;
    assign in1710_1 = {pp54[102]};
    assign in1710_2 = {pp55[101]};
    Full_Adder FA_1710(s1710, c1710, in1710_1, in1710_2, pp53[103]);
    wire[0:0] s1711, in1711_1, in1711_2;
    wire c1711;
    assign in1711_1 = {pp57[99]};
    assign in1711_2 = {pp58[98]};
    Full_Adder FA_1711(s1711, c1711, in1711_1, in1711_2, pp56[100]);
    wire[0:0] s1712, in1712_1, in1712_2;
    wire c1712;
    assign in1712_1 = {pp60[96]};
    assign in1712_2 = {pp61[95]};
    Full_Adder FA_1712(s1712, c1712, in1712_1, in1712_2, pp59[97]);
    wire[0:0] s1713, in1713_1, in1713_2;
    wire c1713;
    assign in1713_1 = {pp63[93]};
    assign in1713_2 = {pp64[92]};
    Full_Adder FA_1713(s1713, c1713, in1713_1, in1713_2, pp62[94]);
    wire[0:0] s1714, in1714_1, in1714_2;
    wire c1714;
    assign in1714_1 = {pp66[90]};
    assign in1714_2 = {pp67[89]};
    Full_Adder FA_1714(s1714, c1714, in1714_1, in1714_2, pp65[91]);
    wire[0:0] s1715, in1715_1, in1715_2;
    wire c1715;
    assign in1715_1 = {pp69[87]};
    assign in1715_2 = {pp70[86]};
    Full_Adder FA_1715(s1715, c1715, in1715_1, in1715_2, pp68[88]);
    wire[0:0] s1716, in1716_1, in1716_2;
    wire c1716;
    assign in1716_1 = {pp31[126]};
    assign in1716_2 = {pp32[125]};
    Full_Adder FA_1716(s1716, c1716, in1716_1, in1716_2, pp30[127]);
    wire[0:0] s1717, in1717_1, in1717_2;
    wire c1717;
    assign in1717_1 = {pp34[123]};
    assign in1717_2 = {pp35[122]};
    Full_Adder FA_1717(s1717, c1717, in1717_1, in1717_2, pp33[124]);
    wire[0:0] s1718, in1718_1, in1718_2;
    wire c1718;
    assign in1718_1 = {pp37[120]};
    assign in1718_2 = {pp38[119]};
    Full_Adder FA_1718(s1718, c1718, in1718_1, in1718_2, pp36[121]);
    wire[0:0] s1719, in1719_1, in1719_2;
    wire c1719;
    assign in1719_1 = {pp40[117]};
    assign in1719_2 = {pp41[116]};
    Full_Adder FA_1719(s1719, c1719, in1719_1, in1719_2, pp39[118]);
    wire[0:0] s1720, in1720_1, in1720_2;
    wire c1720;
    assign in1720_1 = {pp43[114]};
    assign in1720_2 = {pp44[113]};
    Full_Adder FA_1720(s1720, c1720, in1720_1, in1720_2, pp42[115]);
    wire[0:0] s1721, in1721_1, in1721_2;
    wire c1721;
    assign in1721_1 = {pp46[111]};
    assign in1721_2 = {pp47[110]};
    Full_Adder FA_1721(s1721, c1721, in1721_1, in1721_2, pp45[112]);
    wire[0:0] s1722, in1722_1, in1722_2;
    wire c1722;
    assign in1722_1 = {pp49[108]};
    assign in1722_2 = {pp50[107]};
    Full_Adder FA_1722(s1722, c1722, in1722_1, in1722_2, pp48[109]);
    wire[0:0] s1723, in1723_1, in1723_2;
    wire c1723;
    assign in1723_1 = {pp52[105]};
    assign in1723_2 = {pp53[104]};
    Full_Adder FA_1723(s1723, c1723, in1723_1, in1723_2, pp51[106]);
    wire[0:0] s1724, in1724_1, in1724_2;
    wire c1724;
    assign in1724_1 = {pp55[102]};
    assign in1724_2 = {pp56[101]};
    Full_Adder FA_1724(s1724, c1724, in1724_1, in1724_2, pp54[103]);
    wire[0:0] s1725, in1725_1, in1725_2;
    wire c1725;
    assign in1725_1 = {pp58[99]};
    assign in1725_2 = {pp59[98]};
    Full_Adder FA_1725(s1725, c1725, in1725_1, in1725_2, pp57[100]);
    wire[0:0] s1726, in1726_1, in1726_2;
    wire c1726;
    assign in1726_1 = {pp61[96]};
    assign in1726_2 = {pp62[95]};
    Full_Adder FA_1726(s1726, c1726, in1726_1, in1726_2, pp60[97]);
    wire[0:0] s1727, in1727_1, in1727_2;
    wire c1727;
    assign in1727_1 = {pp64[93]};
    assign in1727_2 = {pp65[92]};
    Full_Adder FA_1727(s1727, c1727, in1727_1, in1727_2, pp63[94]);
    wire[0:0] s1728, in1728_1, in1728_2;
    wire c1728;
    assign in1728_1 = {pp67[90]};
    assign in1728_2 = {pp68[89]};
    Full_Adder FA_1728(s1728, c1728, in1728_1, in1728_2, pp66[91]);
    wire[0:0] s1729, in1729_1, in1729_2;
    wire c1729;
    assign in1729_1 = {pp32[126]};
    assign in1729_2 = {pp33[125]};
    Full_Adder FA_1729(s1729, c1729, in1729_1, in1729_2, pp31[127]);
    wire[0:0] s1730, in1730_1, in1730_2;
    wire c1730;
    assign in1730_1 = {pp35[123]};
    assign in1730_2 = {pp36[122]};
    Full_Adder FA_1730(s1730, c1730, in1730_1, in1730_2, pp34[124]);
    wire[0:0] s1731, in1731_1, in1731_2;
    wire c1731;
    assign in1731_1 = {pp38[120]};
    assign in1731_2 = {pp39[119]};
    Full_Adder FA_1731(s1731, c1731, in1731_1, in1731_2, pp37[121]);
    wire[0:0] s1732, in1732_1, in1732_2;
    wire c1732;
    assign in1732_1 = {pp41[117]};
    assign in1732_2 = {pp42[116]};
    Full_Adder FA_1732(s1732, c1732, in1732_1, in1732_2, pp40[118]);
    wire[0:0] s1733, in1733_1, in1733_2;
    wire c1733;
    assign in1733_1 = {pp44[114]};
    assign in1733_2 = {pp45[113]};
    Full_Adder FA_1733(s1733, c1733, in1733_1, in1733_2, pp43[115]);
    wire[0:0] s1734, in1734_1, in1734_2;
    wire c1734;
    assign in1734_1 = {pp47[111]};
    assign in1734_2 = {pp48[110]};
    Full_Adder FA_1734(s1734, c1734, in1734_1, in1734_2, pp46[112]);
    wire[0:0] s1735, in1735_1, in1735_2;
    wire c1735;
    assign in1735_1 = {pp50[108]};
    assign in1735_2 = {pp51[107]};
    Full_Adder FA_1735(s1735, c1735, in1735_1, in1735_2, pp49[109]);
    wire[0:0] s1736, in1736_1, in1736_2;
    wire c1736;
    assign in1736_1 = {pp53[105]};
    assign in1736_2 = {pp54[104]};
    Full_Adder FA_1736(s1736, c1736, in1736_1, in1736_2, pp52[106]);
    wire[0:0] s1737, in1737_1, in1737_2;
    wire c1737;
    assign in1737_1 = {pp56[102]};
    assign in1737_2 = {pp57[101]};
    Full_Adder FA_1737(s1737, c1737, in1737_1, in1737_2, pp55[103]);
    wire[0:0] s1738, in1738_1, in1738_2;
    wire c1738;
    assign in1738_1 = {pp59[99]};
    assign in1738_2 = {pp60[98]};
    Full_Adder FA_1738(s1738, c1738, in1738_1, in1738_2, pp58[100]);
    wire[0:0] s1739, in1739_1, in1739_2;
    wire c1739;
    assign in1739_1 = {pp62[96]};
    assign in1739_2 = {pp63[95]};
    Full_Adder FA_1739(s1739, c1739, in1739_1, in1739_2, pp61[97]);
    wire[0:0] s1740, in1740_1, in1740_2;
    wire c1740;
    assign in1740_1 = {pp65[93]};
    assign in1740_2 = {pp66[92]};
    Full_Adder FA_1740(s1740, c1740, in1740_1, in1740_2, pp64[94]);
    wire[0:0] s1741, in1741_1, in1741_2;
    wire c1741;
    assign in1741_1 = {pp33[126]};
    assign in1741_2 = {pp34[125]};
    Full_Adder FA_1741(s1741, c1741, in1741_1, in1741_2, pp32[127]);
    wire[0:0] s1742, in1742_1, in1742_2;
    wire c1742;
    assign in1742_1 = {pp36[123]};
    assign in1742_2 = {pp37[122]};
    Full_Adder FA_1742(s1742, c1742, in1742_1, in1742_2, pp35[124]);
    wire[0:0] s1743, in1743_1, in1743_2;
    wire c1743;
    assign in1743_1 = {pp39[120]};
    assign in1743_2 = {pp40[119]};
    Full_Adder FA_1743(s1743, c1743, in1743_1, in1743_2, pp38[121]);
    wire[0:0] s1744, in1744_1, in1744_2;
    wire c1744;
    assign in1744_1 = {pp42[117]};
    assign in1744_2 = {pp43[116]};
    Full_Adder FA_1744(s1744, c1744, in1744_1, in1744_2, pp41[118]);
    wire[0:0] s1745, in1745_1, in1745_2;
    wire c1745;
    assign in1745_1 = {pp45[114]};
    assign in1745_2 = {pp46[113]};
    Full_Adder FA_1745(s1745, c1745, in1745_1, in1745_2, pp44[115]);
    wire[0:0] s1746, in1746_1, in1746_2;
    wire c1746;
    assign in1746_1 = {pp48[111]};
    assign in1746_2 = {pp49[110]};
    Full_Adder FA_1746(s1746, c1746, in1746_1, in1746_2, pp47[112]);
    wire[0:0] s1747, in1747_1, in1747_2;
    wire c1747;
    assign in1747_1 = {pp51[108]};
    assign in1747_2 = {pp52[107]};
    Full_Adder FA_1747(s1747, c1747, in1747_1, in1747_2, pp50[109]);
    wire[0:0] s1748, in1748_1, in1748_2;
    wire c1748;
    assign in1748_1 = {pp54[105]};
    assign in1748_2 = {pp55[104]};
    Full_Adder FA_1748(s1748, c1748, in1748_1, in1748_2, pp53[106]);
    wire[0:0] s1749, in1749_1, in1749_2;
    wire c1749;
    assign in1749_1 = {pp57[102]};
    assign in1749_2 = {pp58[101]};
    Full_Adder FA_1749(s1749, c1749, in1749_1, in1749_2, pp56[103]);
    wire[0:0] s1750, in1750_1, in1750_2;
    wire c1750;
    assign in1750_1 = {pp60[99]};
    assign in1750_2 = {pp61[98]};
    Full_Adder FA_1750(s1750, c1750, in1750_1, in1750_2, pp59[100]);
    wire[0:0] s1751, in1751_1, in1751_2;
    wire c1751;
    assign in1751_1 = {pp63[96]};
    assign in1751_2 = {pp64[95]};
    Full_Adder FA_1751(s1751, c1751, in1751_1, in1751_2, pp62[97]);
    wire[0:0] s1752, in1752_1, in1752_2;
    wire c1752;
    assign in1752_1 = {pp34[126]};
    assign in1752_2 = {pp35[125]};
    Full_Adder FA_1752(s1752, c1752, in1752_1, in1752_2, pp33[127]);
    wire[0:0] s1753, in1753_1, in1753_2;
    wire c1753;
    assign in1753_1 = {pp37[123]};
    assign in1753_2 = {pp38[122]};
    Full_Adder FA_1753(s1753, c1753, in1753_1, in1753_2, pp36[124]);
    wire[0:0] s1754, in1754_1, in1754_2;
    wire c1754;
    assign in1754_1 = {pp40[120]};
    assign in1754_2 = {pp41[119]};
    Full_Adder FA_1754(s1754, c1754, in1754_1, in1754_2, pp39[121]);
    wire[0:0] s1755, in1755_1, in1755_2;
    wire c1755;
    assign in1755_1 = {pp43[117]};
    assign in1755_2 = {pp44[116]};
    Full_Adder FA_1755(s1755, c1755, in1755_1, in1755_2, pp42[118]);
    wire[0:0] s1756, in1756_1, in1756_2;
    wire c1756;
    assign in1756_1 = {pp46[114]};
    assign in1756_2 = {pp47[113]};
    Full_Adder FA_1756(s1756, c1756, in1756_1, in1756_2, pp45[115]);
    wire[0:0] s1757, in1757_1, in1757_2;
    wire c1757;
    assign in1757_1 = {pp49[111]};
    assign in1757_2 = {pp50[110]};
    Full_Adder FA_1757(s1757, c1757, in1757_1, in1757_2, pp48[112]);
    wire[0:0] s1758, in1758_1, in1758_2;
    wire c1758;
    assign in1758_1 = {pp52[108]};
    assign in1758_2 = {pp53[107]};
    Full_Adder FA_1758(s1758, c1758, in1758_1, in1758_2, pp51[109]);
    wire[0:0] s1759, in1759_1, in1759_2;
    wire c1759;
    assign in1759_1 = {pp55[105]};
    assign in1759_2 = {pp56[104]};
    Full_Adder FA_1759(s1759, c1759, in1759_1, in1759_2, pp54[106]);
    wire[0:0] s1760, in1760_1, in1760_2;
    wire c1760;
    assign in1760_1 = {pp58[102]};
    assign in1760_2 = {pp59[101]};
    Full_Adder FA_1760(s1760, c1760, in1760_1, in1760_2, pp57[103]);
    wire[0:0] s1761, in1761_1, in1761_2;
    wire c1761;
    assign in1761_1 = {pp61[99]};
    assign in1761_2 = {pp62[98]};
    Full_Adder FA_1761(s1761, c1761, in1761_1, in1761_2, pp60[100]);
    wire[0:0] s1762, in1762_1, in1762_2;
    wire c1762;
    assign in1762_1 = {pp35[126]};
    assign in1762_2 = {pp36[125]};
    Full_Adder FA_1762(s1762, c1762, in1762_1, in1762_2, pp34[127]);
    wire[0:0] s1763, in1763_1, in1763_2;
    wire c1763;
    assign in1763_1 = {pp38[123]};
    assign in1763_2 = {pp39[122]};
    Full_Adder FA_1763(s1763, c1763, in1763_1, in1763_2, pp37[124]);
    wire[0:0] s1764, in1764_1, in1764_2;
    wire c1764;
    assign in1764_1 = {pp41[120]};
    assign in1764_2 = {pp42[119]};
    Full_Adder FA_1764(s1764, c1764, in1764_1, in1764_2, pp40[121]);
    wire[0:0] s1765, in1765_1, in1765_2;
    wire c1765;
    assign in1765_1 = {pp44[117]};
    assign in1765_2 = {pp45[116]};
    Full_Adder FA_1765(s1765, c1765, in1765_1, in1765_2, pp43[118]);
    wire[0:0] s1766, in1766_1, in1766_2;
    wire c1766;
    assign in1766_1 = {pp47[114]};
    assign in1766_2 = {pp48[113]};
    Full_Adder FA_1766(s1766, c1766, in1766_1, in1766_2, pp46[115]);
    wire[0:0] s1767, in1767_1, in1767_2;
    wire c1767;
    assign in1767_1 = {pp50[111]};
    assign in1767_2 = {pp51[110]};
    Full_Adder FA_1767(s1767, c1767, in1767_1, in1767_2, pp49[112]);
    wire[0:0] s1768, in1768_1, in1768_2;
    wire c1768;
    assign in1768_1 = {pp53[108]};
    assign in1768_2 = {pp54[107]};
    Full_Adder FA_1768(s1768, c1768, in1768_1, in1768_2, pp52[109]);
    wire[0:0] s1769, in1769_1, in1769_2;
    wire c1769;
    assign in1769_1 = {pp56[105]};
    assign in1769_2 = {pp57[104]};
    Full_Adder FA_1769(s1769, c1769, in1769_1, in1769_2, pp55[106]);
    wire[0:0] s1770, in1770_1, in1770_2;
    wire c1770;
    assign in1770_1 = {pp59[102]};
    assign in1770_2 = {pp60[101]};
    Full_Adder FA_1770(s1770, c1770, in1770_1, in1770_2, pp58[103]);
    wire[0:0] s1771, in1771_1, in1771_2;
    wire c1771;
    assign in1771_1 = {pp36[126]};
    assign in1771_2 = {pp37[125]};
    Full_Adder FA_1771(s1771, c1771, in1771_1, in1771_2, pp35[127]);
    wire[0:0] s1772, in1772_1, in1772_2;
    wire c1772;
    assign in1772_1 = {pp39[123]};
    assign in1772_2 = {pp40[122]};
    Full_Adder FA_1772(s1772, c1772, in1772_1, in1772_2, pp38[124]);
    wire[0:0] s1773, in1773_1, in1773_2;
    wire c1773;
    assign in1773_1 = {pp42[120]};
    assign in1773_2 = {pp43[119]};
    Full_Adder FA_1773(s1773, c1773, in1773_1, in1773_2, pp41[121]);
    wire[0:0] s1774, in1774_1, in1774_2;
    wire c1774;
    assign in1774_1 = {pp45[117]};
    assign in1774_2 = {pp46[116]};
    Full_Adder FA_1774(s1774, c1774, in1774_1, in1774_2, pp44[118]);
    wire[0:0] s1775, in1775_1, in1775_2;
    wire c1775;
    assign in1775_1 = {pp48[114]};
    assign in1775_2 = {pp49[113]};
    Full_Adder FA_1775(s1775, c1775, in1775_1, in1775_2, pp47[115]);
    wire[0:0] s1776, in1776_1, in1776_2;
    wire c1776;
    assign in1776_1 = {pp51[111]};
    assign in1776_2 = {pp52[110]};
    Full_Adder FA_1776(s1776, c1776, in1776_1, in1776_2, pp50[112]);
    wire[0:0] s1777, in1777_1, in1777_2;
    wire c1777;
    assign in1777_1 = {pp54[108]};
    assign in1777_2 = {pp55[107]};
    Full_Adder FA_1777(s1777, c1777, in1777_1, in1777_2, pp53[109]);
    wire[0:0] s1778, in1778_1, in1778_2;
    wire c1778;
    assign in1778_1 = {pp57[105]};
    assign in1778_2 = {pp58[104]};
    Full_Adder FA_1778(s1778, c1778, in1778_1, in1778_2, pp56[106]);
    wire[0:0] s1779, in1779_1, in1779_2;
    wire c1779;
    assign in1779_1 = {pp37[126]};
    assign in1779_2 = {pp38[125]};
    Full_Adder FA_1779(s1779, c1779, in1779_1, in1779_2, pp36[127]);
    wire[0:0] s1780, in1780_1, in1780_2;
    wire c1780;
    assign in1780_1 = {pp40[123]};
    assign in1780_2 = {pp41[122]};
    Full_Adder FA_1780(s1780, c1780, in1780_1, in1780_2, pp39[124]);
    wire[0:0] s1781, in1781_1, in1781_2;
    wire c1781;
    assign in1781_1 = {pp43[120]};
    assign in1781_2 = {pp44[119]};
    Full_Adder FA_1781(s1781, c1781, in1781_1, in1781_2, pp42[121]);
    wire[0:0] s1782, in1782_1, in1782_2;
    wire c1782;
    assign in1782_1 = {pp46[117]};
    assign in1782_2 = {pp47[116]};
    Full_Adder FA_1782(s1782, c1782, in1782_1, in1782_2, pp45[118]);
    wire[0:0] s1783, in1783_1, in1783_2;
    wire c1783;
    assign in1783_1 = {pp49[114]};
    assign in1783_2 = {pp50[113]};
    Full_Adder FA_1783(s1783, c1783, in1783_1, in1783_2, pp48[115]);
    wire[0:0] s1784, in1784_1, in1784_2;
    wire c1784;
    assign in1784_1 = {pp52[111]};
    assign in1784_2 = {pp53[110]};
    Full_Adder FA_1784(s1784, c1784, in1784_1, in1784_2, pp51[112]);
    wire[0:0] s1785, in1785_1, in1785_2;
    wire c1785;
    assign in1785_1 = {pp55[108]};
    assign in1785_2 = {pp56[107]};
    Full_Adder FA_1785(s1785, c1785, in1785_1, in1785_2, pp54[109]);
    wire[0:0] s1786, in1786_1, in1786_2;
    wire c1786;
    assign in1786_1 = {pp38[126]};
    assign in1786_2 = {pp39[125]};
    Full_Adder FA_1786(s1786, c1786, in1786_1, in1786_2, pp37[127]);
    wire[0:0] s1787, in1787_1, in1787_2;
    wire c1787;
    assign in1787_1 = {pp41[123]};
    assign in1787_2 = {pp42[122]};
    Full_Adder FA_1787(s1787, c1787, in1787_1, in1787_2, pp40[124]);
    wire[0:0] s1788, in1788_1, in1788_2;
    wire c1788;
    assign in1788_1 = {pp44[120]};
    assign in1788_2 = {pp45[119]};
    Full_Adder FA_1788(s1788, c1788, in1788_1, in1788_2, pp43[121]);
    wire[0:0] s1789, in1789_1, in1789_2;
    wire c1789;
    assign in1789_1 = {pp47[117]};
    assign in1789_2 = {pp48[116]};
    Full_Adder FA_1789(s1789, c1789, in1789_1, in1789_2, pp46[118]);
    wire[0:0] s1790, in1790_1, in1790_2;
    wire c1790;
    assign in1790_1 = {pp50[114]};
    assign in1790_2 = {pp51[113]};
    Full_Adder FA_1790(s1790, c1790, in1790_1, in1790_2, pp49[115]);
    wire[0:0] s1791, in1791_1, in1791_2;
    wire c1791;
    assign in1791_1 = {pp53[111]};
    assign in1791_2 = {pp54[110]};
    Full_Adder FA_1791(s1791, c1791, in1791_1, in1791_2, pp52[112]);
    wire[0:0] s1792, in1792_1, in1792_2;
    wire c1792;
    assign in1792_1 = {pp39[126]};
    assign in1792_2 = {pp40[125]};
    Full_Adder FA_1792(s1792, c1792, in1792_1, in1792_2, pp38[127]);
    wire[0:0] s1793, in1793_1, in1793_2;
    wire c1793;
    assign in1793_1 = {pp42[123]};
    assign in1793_2 = {pp43[122]};
    Full_Adder FA_1793(s1793, c1793, in1793_1, in1793_2, pp41[124]);
    wire[0:0] s1794, in1794_1, in1794_2;
    wire c1794;
    assign in1794_1 = {pp45[120]};
    assign in1794_2 = {pp46[119]};
    Full_Adder FA_1794(s1794, c1794, in1794_1, in1794_2, pp44[121]);
    wire[0:0] s1795, in1795_1, in1795_2;
    wire c1795;
    assign in1795_1 = {pp48[117]};
    assign in1795_2 = {pp49[116]};
    Full_Adder FA_1795(s1795, c1795, in1795_1, in1795_2, pp47[118]);
    wire[0:0] s1796, in1796_1, in1796_2;
    wire c1796;
    assign in1796_1 = {pp51[114]};
    assign in1796_2 = {pp52[113]};
    Full_Adder FA_1796(s1796, c1796, in1796_1, in1796_2, pp50[115]);
    wire[0:0] s1797, in1797_1, in1797_2;
    wire c1797;
    assign in1797_1 = {pp40[126]};
    assign in1797_2 = {pp41[125]};
    Full_Adder FA_1797(s1797, c1797, in1797_1, in1797_2, pp39[127]);
    wire[0:0] s1798, in1798_1, in1798_2;
    wire c1798;
    assign in1798_1 = {pp43[123]};
    assign in1798_2 = {pp44[122]};
    Full_Adder FA_1798(s1798, c1798, in1798_1, in1798_2, pp42[124]);
    wire[0:0] s1799, in1799_1, in1799_2;
    wire c1799;
    assign in1799_1 = {pp46[120]};
    assign in1799_2 = {pp47[119]};
    Full_Adder FA_1799(s1799, c1799, in1799_1, in1799_2, pp45[121]);
    wire[0:0] s1800, in1800_1, in1800_2;
    wire c1800;
    assign in1800_1 = {pp49[117]};
    assign in1800_2 = {pp50[116]};
    Full_Adder FA_1800(s1800, c1800, in1800_1, in1800_2, pp48[118]);
    wire[0:0] s1801, in1801_1, in1801_2;
    wire c1801;
    assign in1801_1 = {pp41[126]};
    assign in1801_2 = {pp42[125]};
    Full_Adder FA_1801(s1801, c1801, in1801_1, in1801_2, pp40[127]);
    wire[0:0] s1802, in1802_1, in1802_2;
    wire c1802;
    assign in1802_1 = {pp44[123]};
    assign in1802_2 = {pp45[122]};
    Full_Adder FA_1802(s1802, c1802, in1802_1, in1802_2, pp43[124]);
    wire[0:0] s1803, in1803_1, in1803_2;
    wire c1803;
    assign in1803_1 = {pp47[120]};
    assign in1803_2 = {pp48[119]};
    Full_Adder FA_1803(s1803, c1803, in1803_1, in1803_2, pp46[121]);
    wire[0:0] s1804, in1804_1, in1804_2;
    wire c1804;
    assign in1804_1 = {pp42[126]};
    assign in1804_2 = {pp43[125]};
    Full_Adder FA_1804(s1804, c1804, in1804_1, in1804_2, pp41[127]);
    wire[0:0] s1805, in1805_1, in1805_2;
    wire c1805;
    assign in1805_1 = {pp45[123]};
    assign in1805_2 = {pp46[122]};
    Full_Adder FA_1805(s1805, c1805, in1805_1, in1805_2, pp44[124]);
    wire[0:0] s1806, in1806_1, in1806_2;
    wire c1806;
    assign in1806_1 = {pp43[126]};
    assign in1806_2 = {pp44[125]};
    Full_Adder FA_1806(s1806, c1806, in1806_1, in1806_2, pp42[127]);

    /*Stage 2*/
    wire[0:0] s1807, in1807_1, in1807_2;
    wire c1807;
    assign in1807_1 = {pp0[58]};
    assign in1807_2 = {pp1[57]};
    Half_Adder HA_1807(s1807, c1807, in1807_1, in1807_2);
    wire[0:0] s1808, in1808_1, in1808_2;
    wire c1808;
    assign in1808_1 = {pp1[58]};
    assign in1808_2 = {pp2[57]};
    Full_Adder FA_1808(s1808, c1808, in1808_1, in1808_2, pp0[59]);
    wire[0:0] s1809, in1809_1, in1809_2;
    wire c1809;
    assign in1809_1 = {pp3[56]};
    assign in1809_2 = {pp4[55]};
    Half_Adder HA_1809(s1809, c1809, in1809_1, in1809_2);
    wire[0:0] s1810, in1810_1, in1810_2;
    wire c1810;
    assign in1810_1 = {pp1[59]};
    assign in1810_2 = {pp2[58]};
    Full_Adder FA_1810(s1810, c1810, in1810_1, in1810_2, pp0[60]);
    wire[0:0] s1811, in1811_1, in1811_2;
    wire c1811;
    assign in1811_1 = {pp4[56]};
    assign in1811_2 = {pp5[55]};
    Full_Adder FA_1811(s1811, c1811, in1811_1, in1811_2, pp3[57]);
    wire[0:0] s1812, in1812_1, in1812_2;
    wire c1812;
    assign in1812_1 = {pp6[54]};
    assign in1812_2 = {pp7[53]};
    Half_Adder HA_1812(s1812, c1812, in1812_1, in1812_2);
    wire[0:0] s1813, in1813_1, in1813_2;
    wire c1813;
    assign in1813_1 = {pp1[60]};
    assign in1813_2 = {pp2[59]};
    Full_Adder FA_1813(s1813, c1813, in1813_1, in1813_2, pp0[61]);
    wire[0:0] s1814, in1814_1, in1814_2;
    wire c1814;
    assign in1814_1 = {pp4[57]};
    assign in1814_2 = {pp5[56]};
    Full_Adder FA_1814(s1814, c1814, in1814_1, in1814_2, pp3[58]);
    wire[0:0] s1815, in1815_1, in1815_2;
    wire c1815;
    assign in1815_1 = {pp7[54]};
    assign in1815_2 = {pp8[53]};
    Full_Adder FA_1815(s1815, c1815, in1815_1, in1815_2, pp6[55]);
    wire[0:0] s1816, in1816_1, in1816_2;
    wire c1816;
    assign in1816_1 = {pp9[52]};
    assign in1816_2 = {pp10[51]};
    Half_Adder HA_1816(s1816, c1816, in1816_1, in1816_2);
    wire[0:0] s1817, in1817_1, in1817_2;
    wire c1817;
    assign in1817_1 = {pp1[61]};
    assign in1817_2 = {pp2[60]};
    Full_Adder FA_1817(s1817, c1817, in1817_1, in1817_2, pp0[62]);
    wire[0:0] s1818, in1818_1, in1818_2;
    wire c1818;
    assign in1818_1 = {pp4[58]};
    assign in1818_2 = {pp5[57]};
    Full_Adder FA_1818(s1818, c1818, in1818_1, in1818_2, pp3[59]);
    wire[0:0] s1819, in1819_1, in1819_2;
    wire c1819;
    assign in1819_1 = {pp7[55]};
    assign in1819_2 = {pp8[54]};
    Full_Adder FA_1819(s1819, c1819, in1819_1, in1819_2, pp6[56]);
    wire[0:0] s1820, in1820_1, in1820_2;
    wire c1820;
    assign in1820_1 = {pp10[52]};
    assign in1820_2 = {pp11[51]};
    Full_Adder FA_1820(s1820, c1820, in1820_1, in1820_2, pp9[53]);
    wire[0:0] s1821, in1821_1, in1821_2;
    wire c1821;
    assign in1821_1 = {pp12[50]};
    assign in1821_2 = {pp13[49]};
    Half_Adder HA_1821(s1821, c1821, in1821_1, in1821_2);
    wire[0:0] s1822, in1822_1, in1822_2;
    wire c1822;
    assign in1822_1 = {pp1[62]};
    assign in1822_2 = {pp2[61]};
    Full_Adder FA_1822(s1822, c1822, in1822_1, in1822_2, pp0[63]);
    wire[0:0] s1823, in1823_1, in1823_2;
    wire c1823;
    assign in1823_1 = {pp4[59]};
    assign in1823_2 = {pp5[58]};
    Full_Adder FA_1823(s1823, c1823, in1823_1, in1823_2, pp3[60]);
    wire[0:0] s1824, in1824_1, in1824_2;
    wire c1824;
    assign in1824_1 = {pp7[56]};
    assign in1824_2 = {pp8[55]};
    Full_Adder FA_1824(s1824, c1824, in1824_1, in1824_2, pp6[57]);
    wire[0:0] s1825, in1825_1, in1825_2;
    wire c1825;
    assign in1825_1 = {pp10[53]};
    assign in1825_2 = {pp11[52]};
    Full_Adder FA_1825(s1825, c1825, in1825_1, in1825_2, pp9[54]);
    wire[0:0] s1826, in1826_1, in1826_2;
    wire c1826;
    assign in1826_1 = {pp13[50]};
    assign in1826_2 = {pp14[49]};
    Full_Adder FA_1826(s1826, c1826, in1826_1, in1826_2, pp12[51]);
    wire[0:0] s1827, in1827_1, in1827_2;
    wire c1827;
    assign in1827_1 = {pp15[48]};
    assign in1827_2 = {pp16[47]};
    Half_Adder HA_1827(s1827, c1827, in1827_1, in1827_2);
    wire[0:0] s1828, in1828_1, in1828_2;
    wire c1828;
    assign in1828_1 = {pp1[63]};
    assign in1828_2 = {pp2[62]};
    Full_Adder FA_1828(s1828, c1828, in1828_1, in1828_2, pp0[64]);
    wire[0:0] s1829, in1829_1, in1829_2;
    wire c1829;
    assign in1829_1 = {pp4[60]};
    assign in1829_2 = {pp5[59]};
    Full_Adder FA_1829(s1829, c1829, in1829_1, in1829_2, pp3[61]);
    wire[0:0] s1830, in1830_1, in1830_2;
    wire c1830;
    assign in1830_1 = {pp7[57]};
    assign in1830_2 = {pp8[56]};
    Full_Adder FA_1830(s1830, c1830, in1830_1, in1830_2, pp6[58]);
    wire[0:0] s1831, in1831_1, in1831_2;
    wire c1831;
    assign in1831_1 = {pp10[54]};
    assign in1831_2 = {pp11[53]};
    Full_Adder FA_1831(s1831, c1831, in1831_1, in1831_2, pp9[55]);
    wire[0:0] s1832, in1832_1, in1832_2;
    wire c1832;
    assign in1832_1 = {pp13[51]};
    assign in1832_2 = {pp14[50]};
    Full_Adder FA_1832(s1832, c1832, in1832_1, in1832_2, pp12[52]);
    wire[0:0] s1833, in1833_1, in1833_2;
    wire c1833;
    assign in1833_1 = {pp16[48]};
    assign in1833_2 = {pp17[47]};
    Full_Adder FA_1833(s1833, c1833, in1833_1, in1833_2, pp15[49]);
    wire[0:0] s1834, in1834_1, in1834_2;
    wire c1834;
    assign in1834_1 = {pp18[46]};
    assign in1834_2 = {pp19[45]};
    Half_Adder HA_1834(s1834, c1834, in1834_1, in1834_2);
    wire[0:0] s1835, in1835_1, in1835_2;
    wire c1835;
    assign in1835_1 = {pp1[64]};
    assign in1835_2 = {pp2[63]};
    Full_Adder FA_1835(s1835, c1835, in1835_1, in1835_2, pp0[65]);
    wire[0:0] s1836, in1836_1, in1836_2;
    wire c1836;
    assign in1836_1 = {pp4[61]};
    assign in1836_2 = {pp5[60]};
    Full_Adder FA_1836(s1836, c1836, in1836_1, in1836_2, pp3[62]);
    wire[0:0] s1837, in1837_1, in1837_2;
    wire c1837;
    assign in1837_1 = {pp7[58]};
    assign in1837_2 = {pp8[57]};
    Full_Adder FA_1837(s1837, c1837, in1837_1, in1837_2, pp6[59]);
    wire[0:0] s1838, in1838_1, in1838_2;
    wire c1838;
    assign in1838_1 = {pp10[55]};
    assign in1838_2 = {pp11[54]};
    Full_Adder FA_1838(s1838, c1838, in1838_1, in1838_2, pp9[56]);
    wire[0:0] s1839, in1839_1, in1839_2;
    wire c1839;
    assign in1839_1 = {pp13[52]};
    assign in1839_2 = {pp14[51]};
    Full_Adder FA_1839(s1839, c1839, in1839_1, in1839_2, pp12[53]);
    wire[0:0] s1840, in1840_1, in1840_2;
    wire c1840;
    assign in1840_1 = {pp16[49]};
    assign in1840_2 = {pp17[48]};
    Full_Adder FA_1840(s1840, c1840, in1840_1, in1840_2, pp15[50]);
    wire[0:0] s1841, in1841_1, in1841_2;
    wire c1841;
    assign in1841_1 = {pp19[46]};
    assign in1841_2 = {pp20[45]};
    Full_Adder FA_1841(s1841, c1841, in1841_1, in1841_2, pp18[47]);
    wire[0:0] s1842, in1842_1, in1842_2;
    wire c1842;
    assign in1842_1 = {pp21[44]};
    assign in1842_2 = {pp22[43]};
    Half_Adder HA_1842(s1842, c1842, in1842_1, in1842_2);
    wire[0:0] s1843, in1843_1, in1843_2;
    wire c1843;
    assign in1843_1 = {pp1[65]};
    assign in1843_2 = {pp2[64]};
    Full_Adder FA_1843(s1843, c1843, in1843_1, in1843_2, pp0[66]);
    wire[0:0] s1844, in1844_1, in1844_2;
    wire c1844;
    assign in1844_1 = {pp4[62]};
    assign in1844_2 = {pp5[61]};
    Full_Adder FA_1844(s1844, c1844, in1844_1, in1844_2, pp3[63]);
    wire[0:0] s1845, in1845_1, in1845_2;
    wire c1845;
    assign in1845_1 = {pp7[59]};
    assign in1845_2 = {pp8[58]};
    Full_Adder FA_1845(s1845, c1845, in1845_1, in1845_2, pp6[60]);
    wire[0:0] s1846, in1846_1, in1846_2;
    wire c1846;
    assign in1846_1 = {pp10[56]};
    assign in1846_2 = {pp11[55]};
    Full_Adder FA_1846(s1846, c1846, in1846_1, in1846_2, pp9[57]);
    wire[0:0] s1847, in1847_1, in1847_2;
    wire c1847;
    assign in1847_1 = {pp13[53]};
    assign in1847_2 = {pp14[52]};
    Full_Adder FA_1847(s1847, c1847, in1847_1, in1847_2, pp12[54]);
    wire[0:0] s1848, in1848_1, in1848_2;
    wire c1848;
    assign in1848_1 = {pp16[50]};
    assign in1848_2 = {pp17[49]};
    Full_Adder FA_1848(s1848, c1848, in1848_1, in1848_2, pp15[51]);
    wire[0:0] s1849, in1849_1, in1849_2;
    wire c1849;
    assign in1849_1 = {pp19[47]};
    assign in1849_2 = {pp20[46]};
    Full_Adder FA_1849(s1849, c1849, in1849_1, in1849_2, pp18[48]);
    wire[0:0] s1850, in1850_1, in1850_2;
    wire c1850;
    assign in1850_1 = {pp22[44]};
    assign in1850_2 = {pp23[43]};
    Full_Adder FA_1850(s1850, c1850, in1850_1, in1850_2, pp21[45]);
    wire[0:0] s1851, in1851_1, in1851_2;
    wire c1851;
    assign in1851_1 = {pp24[42]};
    assign in1851_2 = {pp25[41]};
    Half_Adder HA_1851(s1851, c1851, in1851_1, in1851_2);
    wire[0:0] s1852, in1852_1, in1852_2;
    wire c1852;
    assign in1852_1 = {pp1[66]};
    assign in1852_2 = {pp2[65]};
    Full_Adder FA_1852(s1852, c1852, in1852_1, in1852_2, pp0[67]);
    wire[0:0] s1853, in1853_1, in1853_2;
    wire c1853;
    assign in1853_1 = {pp4[63]};
    assign in1853_2 = {pp5[62]};
    Full_Adder FA_1853(s1853, c1853, in1853_1, in1853_2, pp3[64]);
    wire[0:0] s1854, in1854_1, in1854_2;
    wire c1854;
    assign in1854_1 = {pp7[60]};
    assign in1854_2 = {pp8[59]};
    Full_Adder FA_1854(s1854, c1854, in1854_1, in1854_2, pp6[61]);
    wire[0:0] s1855, in1855_1, in1855_2;
    wire c1855;
    assign in1855_1 = {pp10[57]};
    assign in1855_2 = {pp11[56]};
    Full_Adder FA_1855(s1855, c1855, in1855_1, in1855_2, pp9[58]);
    wire[0:0] s1856, in1856_1, in1856_2;
    wire c1856;
    assign in1856_1 = {pp13[54]};
    assign in1856_2 = {pp14[53]};
    Full_Adder FA_1856(s1856, c1856, in1856_1, in1856_2, pp12[55]);
    wire[0:0] s1857, in1857_1, in1857_2;
    wire c1857;
    assign in1857_1 = {pp16[51]};
    assign in1857_2 = {pp17[50]};
    Full_Adder FA_1857(s1857, c1857, in1857_1, in1857_2, pp15[52]);
    wire[0:0] s1858, in1858_1, in1858_2;
    wire c1858;
    assign in1858_1 = {pp19[48]};
    assign in1858_2 = {pp20[47]};
    Full_Adder FA_1858(s1858, c1858, in1858_1, in1858_2, pp18[49]);
    wire[0:0] s1859, in1859_1, in1859_2;
    wire c1859;
    assign in1859_1 = {pp22[45]};
    assign in1859_2 = {pp23[44]};
    Full_Adder FA_1859(s1859, c1859, in1859_1, in1859_2, pp21[46]);
    wire[0:0] s1860, in1860_1, in1860_2;
    wire c1860;
    assign in1860_1 = {pp25[42]};
    assign in1860_2 = {pp26[41]};
    Full_Adder FA_1860(s1860, c1860, in1860_1, in1860_2, pp24[43]);
    wire[0:0] s1861, in1861_1, in1861_2;
    wire c1861;
    assign in1861_1 = {pp27[40]};
    assign in1861_2 = {pp28[39]};
    Half_Adder HA_1861(s1861, c1861, in1861_1, in1861_2);
    wire[0:0] s1862, in1862_1, in1862_2;
    wire c1862;
    assign in1862_1 = {pp1[67]};
    assign in1862_2 = {pp2[66]};
    Full_Adder FA_1862(s1862, c1862, in1862_1, in1862_2, pp0[68]);
    wire[0:0] s1863, in1863_1, in1863_2;
    wire c1863;
    assign in1863_1 = {pp4[64]};
    assign in1863_2 = {pp5[63]};
    Full_Adder FA_1863(s1863, c1863, in1863_1, in1863_2, pp3[65]);
    wire[0:0] s1864, in1864_1, in1864_2;
    wire c1864;
    assign in1864_1 = {pp7[61]};
    assign in1864_2 = {pp8[60]};
    Full_Adder FA_1864(s1864, c1864, in1864_1, in1864_2, pp6[62]);
    wire[0:0] s1865, in1865_1, in1865_2;
    wire c1865;
    assign in1865_1 = {pp10[58]};
    assign in1865_2 = {pp11[57]};
    Full_Adder FA_1865(s1865, c1865, in1865_1, in1865_2, pp9[59]);
    wire[0:0] s1866, in1866_1, in1866_2;
    wire c1866;
    assign in1866_1 = {pp13[55]};
    assign in1866_2 = {pp14[54]};
    Full_Adder FA_1866(s1866, c1866, in1866_1, in1866_2, pp12[56]);
    wire[0:0] s1867, in1867_1, in1867_2;
    wire c1867;
    assign in1867_1 = {pp16[52]};
    assign in1867_2 = {pp17[51]};
    Full_Adder FA_1867(s1867, c1867, in1867_1, in1867_2, pp15[53]);
    wire[0:0] s1868, in1868_1, in1868_2;
    wire c1868;
    assign in1868_1 = {pp19[49]};
    assign in1868_2 = {pp20[48]};
    Full_Adder FA_1868(s1868, c1868, in1868_1, in1868_2, pp18[50]);
    wire[0:0] s1869, in1869_1, in1869_2;
    wire c1869;
    assign in1869_1 = {pp22[46]};
    assign in1869_2 = {pp23[45]};
    Full_Adder FA_1869(s1869, c1869, in1869_1, in1869_2, pp21[47]);
    wire[0:0] s1870, in1870_1, in1870_2;
    wire c1870;
    assign in1870_1 = {pp25[43]};
    assign in1870_2 = {pp26[42]};
    Full_Adder FA_1870(s1870, c1870, in1870_1, in1870_2, pp24[44]);
    wire[0:0] s1871, in1871_1, in1871_2;
    wire c1871;
    assign in1871_1 = {pp28[40]};
    assign in1871_2 = {pp29[39]};
    Full_Adder FA_1871(s1871, c1871, in1871_1, in1871_2, pp27[41]);
    wire[0:0] s1872, in1872_1, in1872_2;
    wire c1872;
    assign in1872_1 = {pp30[38]};
    assign in1872_2 = {pp31[37]};
    Half_Adder HA_1872(s1872, c1872, in1872_1, in1872_2);
    wire[0:0] s1873, in1873_1, in1873_2;
    wire c1873;
    assign in1873_1 = {pp1[68]};
    assign in1873_2 = {pp2[67]};
    Full_Adder FA_1873(s1873, c1873, in1873_1, in1873_2, pp0[69]);
    wire[0:0] s1874, in1874_1, in1874_2;
    wire c1874;
    assign in1874_1 = {pp4[65]};
    assign in1874_2 = {pp5[64]};
    Full_Adder FA_1874(s1874, c1874, in1874_1, in1874_2, pp3[66]);
    wire[0:0] s1875, in1875_1, in1875_2;
    wire c1875;
    assign in1875_1 = {pp7[62]};
    assign in1875_2 = {pp8[61]};
    Full_Adder FA_1875(s1875, c1875, in1875_1, in1875_2, pp6[63]);
    wire[0:0] s1876, in1876_1, in1876_2;
    wire c1876;
    assign in1876_1 = {pp10[59]};
    assign in1876_2 = {pp11[58]};
    Full_Adder FA_1876(s1876, c1876, in1876_1, in1876_2, pp9[60]);
    wire[0:0] s1877, in1877_1, in1877_2;
    wire c1877;
    assign in1877_1 = {pp13[56]};
    assign in1877_2 = {pp14[55]};
    Full_Adder FA_1877(s1877, c1877, in1877_1, in1877_2, pp12[57]);
    wire[0:0] s1878, in1878_1, in1878_2;
    wire c1878;
    assign in1878_1 = {pp16[53]};
    assign in1878_2 = {pp17[52]};
    Full_Adder FA_1878(s1878, c1878, in1878_1, in1878_2, pp15[54]);
    wire[0:0] s1879, in1879_1, in1879_2;
    wire c1879;
    assign in1879_1 = {pp19[50]};
    assign in1879_2 = {pp20[49]};
    Full_Adder FA_1879(s1879, c1879, in1879_1, in1879_2, pp18[51]);
    wire[0:0] s1880, in1880_1, in1880_2;
    wire c1880;
    assign in1880_1 = {pp22[47]};
    assign in1880_2 = {pp23[46]};
    Full_Adder FA_1880(s1880, c1880, in1880_1, in1880_2, pp21[48]);
    wire[0:0] s1881, in1881_1, in1881_2;
    wire c1881;
    assign in1881_1 = {pp25[44]};
    assign in1881_2 = {pp26[43]};
    Full_Adder FA_1881(s1881, c1881, in1881_1, in1881_2, pp24[45]);
    wire[0:0] s1882, in1882_1, in1882_2;
    wire c1882;
    assign in1882_1 = {pp28[41]};
    assign in1882_2 = {pp29[40]};
    Full_Adder FA_1882(s1882, c1882, in1882_1, in1882_2, pp27[42]);
    wire[0:0] s1883, in1883_1, in1883_2;
    wire c1883;
    assign in1883_1 = {pp31[38]};
    assign in1883_2 = {pp32[37]};
    Full_Adder FA_1883(s1883, c1883, in1883_1, in1883_2, pp30[39]);
    wire[0:0] s1884, in1884_1, in1884_2;
    wire c1884;
    assign in1884_1 = {pp33[36]};
    assign in1884_2 = {pp34[35]};
    Half_Adder HA_1884(s1884, c1884, in1884_1, in1884_2);
    wire[0:0] s1885, in1885_1, in1885_2;
    wire c1885;
    assign in1885_1 = {pp1[69]};
    assign in1885_2 = {pp2[68]};
    Full_Adder FA_1885(s1885, c1885, in1885_1, in1885_2, pp0[70]);
    wire[0:0] s1886, in1886_1, in1886_2;
    wire c1886;
    assign in1886_1 = {pp4[66]};
    assign in1886_2 = {pp5[65]};
    Full_Adder FA_1886(s1886, c1886, in1886_1, in1886_2, pp3[67]);
    wire[0:0] s1887, in1887_1, in1887_2;
    wire c1887;
    assign in1887_1 = {pp7[63]};
    assign in1887_2 = {pp8[62]};
    Full_Adder FA_1887(s1887, c1887, in1887_1, in1887_2, pp6[64]);
    wire[0:0] s1888, in1888_1, in1888_2;
    wire c1888;
    assign in1888_1 = {pp10[60]};
    assign in1888_2 = {pp11[59]};
    Full_Adder FA_1888(s1888, c1888, in1888_1, in1888_2, pp9[61]);
    wire[0:0] s1889, in1889_1, in1889_2;
    wire c1889;
    assign in1889_1 = {pp13[57]};
    assign in1889_2 = {pp14[56]};
    Full_Adder FA_1889(s1889, c1889, in1889_1, in1889_2, pp12[58]);
    wire[0:0] s1890, in1890_1, in1890_2;
    wire c1890;
    assign in1890_1 = {pp16[54]};
    assign in1890_2 = {pp17[53]};
    Full_Adder FA_1890(s1890, c1890, in1890_1, in1890_2, pp15[55]);
    wire[0:0] s1891, in1891_1, in1891_2;
    wire c1891;
    assign in1891_1 = {pp19[51]};
    assign in1891_2 = {pp20[50]};
    Full_Adder FA_1891(s1891, c1891, in1891_1, in1891_2, pp18[52]);
    wire[0:0] s1892, in1892_1, in1892_2;
    wire c1892;
    assign in1892_1 = {pp22[48]};
    assign in1892_2 = {pp23[47]};
    Full_Adder FA_1892(s1892, c1892, in1892_1, in1892_2, pp21[49]);
    wire[0:0] s1893, in1893_1, in1893_2;
    wire c1893;
    assign in1893_1 = {pp25[45]};
    assign in1893_2 = {pp26[44]};
    Full_Adder FA_1893(s1893, c1893, in1893_1, in1893_2, pp24[46]);
    wire[0:0] s1894, in1894_1, in1894_2;
    wire c1894;
    assign in1894_1 = {pp28[42]};
    assign in1894_2 = {pp29[41]};
    Full_Adder FA_1894(s1894, c1894, in1894_1, in1894_2, pp27[43]);
    wire[0:0] s1895, in1895_1, in1895_2;
    wire c1895;
    assign in1895_1 = {pp31[39]};
    assign in1895_2 = {pp32[38]};
    Full_Adder FA_1895(s1895, c1895, in1895_1, in1895_2, pp30[40]);
    wire[0:0] s1896, in1896_1, in1896_2;
    wire c1896;
    assign in1896_1 = {pp34[36]};
    assign in1896_2 = {pp35[35]};
    Full_Adder FA_1896(s1896, c1896, in1896_1, in1896_2, pp33[37]);
    wire[0:0] s1897, in1897_1, in1897_2;
    wire c1897;
    assign in1897_1 = {pp36[34]};
    assign in1897_2 = {pp37[33]};
    Half_Adder HA_1897(s1897, c1897, in1897_1, in1897_2);
    wire[0:0] s1898, in1898_1, in1898_2;
    wire c1898;
    assign in1898_1 = {pp1[70]};
    assign in1898_2 = {pp2[69]};
    Full_Adder FA_1898(s1898, c1898, in1898_1, in1898_2, pp0[71]);
    wire[0:0] s1899, in1899_1, in1899_2;
    wire c1899;
    assign in1899_1 = {pp4[67]};
    assign in1899_2 = {pp5[66]};
    Full_Adder FA_1899(s1899, c1899, in1899_1, in1899_2, pp3[68]);
    wire[0:0] s1900, in1900_1, in1900_2;
    wire c1900;
    assign in1900_1 = {pp7[64]};
    assign in1900_2 = {pp8[63]};
    Full_Adder FA_1900(s1900, c1900, in1900_1, in1900_2, pp6[65]);
    wire[0:0] s1901, in1901_1, in1901_2;
    wire c1901;
    assign in1901_1 = {pp10[61]};
    assign in1901_2 = {pp11[60]};
    Full_Adder FA_1901(s1901, c1901, in1901_1, in1901_2, pp9[62]);
    wire[0:0] s1902, in1902_1, in1902_2;
    wire c1902;
    assign in1902_1 = {pp13[58]};
    assign in1902_2 = {pp14[57]};
    Full_Adder FA_1902(s1902, c1902, in1902_1, in1902_2, pp12[59]);
    wire[0:0] s1903, in1903_1, in1903_2;
    wire c1903;
    assign in1903_1 = {pp16[55]};
    assign in1903_2 = {pp17[54]};
    Full_Adder FA_1903(s1903, c1903, in1903_1, in1903_2, pp15[56]);
    wire[0:0] s1904, in1904_1, in1904_2;
    wire c1904;
    assign in1904_1 = {pp19[52]};
    assign in1904_2 = {pp20[51]};
    Full_Adder FA_1904(s1904, c1904, in1904_1, in1904_2, pp18[53]);
    wire[0:0] s1905, in1905_1, in1905_2;
    wire c1905;
    assign in1905_1 = {pp22[49]};
    assign in1905_2 = {pp23[48]};
    Full_Adder FA_1905(s1905, c1905, in1905_1, in1905_2, pp21[50]);
    wire[0:0] s1906, in1906_1, in1906_2;
    wire c1906;
    assign in1906_1 = {pp25[46]};
    assign in1906_2 = {pp26[45]};
    Full_Adder FA_1906(s1906, c1906, in1906_1, in1906_2, pp24[47]);
    wire[0:0] s1907, in1907_1, in1907_2;
    wire c1907;
    assign in1907_1 = {pp28[43]};
    assign in1907_2 = {pp29[42]};
    Full_Adder FA_1907(s1907, c1907, in1907_1, in1907_2, pp27[44]);
    wire[0:0] s1908, in1908_1, in1908_2;
    wire c1908;
    assign in1908_1 = {pp31[40]};
    assign in1908_2 = {pp32[39]};
    Full_Adder FA_1908(s1908, c1908, in1908_1, in1908_2, pp30[41]);
    wire[0:0] s1909, in1909_1, in1909_2;
    wire c1909;
    assign in1909_1 = {pp34[37]};
    assign in1909_2 = {pp35[36]};
    Full_Adder FA_1909(s1909, c1909, in1909_1, in1909_2, pp33[38]);
    wire[0:0] s1910, in1910_1, in1910_2;
    wire c1910;
    assign in1910_1 = {pp37[34]};
    assign in1910_2 = {pp38[33]};
    Full_Adder FA_1910(s1910, c1910, in1910_1, in1910_2, pp36[35]);
    wire[0:0] s1911, in1911_1, in1911_2;
    wire c1911;
    assign in1911_1 = {pp39[32]};
    assign in1911_2 = {pp40[31]};
    Half_Adder HA_1911(s1911, c1911, in1911_1, in1911_2);
    wire[0:0] s1912, in1912_1, in1912_2;
    wire c1912;
    assign in1912_1 = {pp1[71]};
    assign in1912_2 = {pp2[70]};
    Full_Adder FA_1912(s1912, c1912, in1912_1, in1912_2, pp0[72]);
    wire[0:0] s1913, in1913_1, in1913_2;
    wire c1913;
    assign in1913_1 = {pp4[68]};
    assign in1913_2 = {pp5[67]};
    Full_Adder FA_1913(s1913, c1913, in1913_1, in1913_2, pp3[69]);
    wire[0:0] s1914, in1914_1, in1914_2;
    wire c1914;
    assign in1914_1 = {pp7[65]};
    assign in1914_2 = {pp8[64]};
    Full_Adder FA_1914(s1914, c1914, in1914_1, in1914_2, pp6[66]);
    wire[0:0] s1915, in1915_1, in1915_2;
    wire c1915;
    assign in1915_1 = {pp10[62]};
    assign in1915_2 = {pp11[61]};
    Full_Adder FA_1915(s1915, c1915, in1915_1, in1915_2, pp9[63]);
    wire[0:0] s1916, in1916_1, in1916_2;
    wire c1916;
    assign in1916_1 = {pp13[59]};
    assign in1916_2 = {pp14[58]};
    Full_Adder FA_1916(s1916, c1916, in1916_1, in1916_2, pp12[60]);
    wire[0:0] s1917, in1917_1, in1917_2;
    wire c1917;
    assign in1917_1 = {pp16[56]};
    assign in1917_2 = {pp17[55]};
    Full_Adder FA_1917(s1917, c1917, in1917_1, in1917_2, pp15[57]);
    wire[0:0] s1918, in1918_1, in1918_2;
    wire c1918;
    assign in1918_1 = {pp19[53]};
    assign in1918_2 = {pp20[52]};
    Full_Adder FA_1918(s1918, c1918, in1918_1, in1918_2, pp18[54]);
    wire[0:0] s1919, in1919_1, in1919_2;
    wire c1919;
    assign in1919_1 = {pp22[50]};
    assign in1919_2 = {pp23[49]};
    Full_Adder FA_1919(s1919, c1919, in1919_1, in1919_2, pp21[51]);
    wire[0:0] s1920, in1920_1, in1920_2;
    wire c1920;
    assign in1920_1 = {pp25[47]};
    assign in1920_2 = {pp26[46]};
    Full_Adder FA_1920(s1920, c1920, in1920_1, in1920_2, pp24[48]);
    wire[0:0] s1921, in1921_1, in1921_2;
    wire c1921;
    assign in1921_1 = {pp28[44]};
    assign in1921_2 = {pp29[43]};
    Full_Adder FA_1921(s1921, c1921, in1921_1, in1921_2, pp27[45]);
    wire[0:0] s1922, in1922_1, in1922_2;
    wire c1922;
    assign in1922_1 = {pp31[41]};
    assign in1922_2 = {pp32[40]};
    Full_Adder FA_1922(s1922, c1922, in1922_1, in1922_2, pp30[42]);
    wire[0:0] s1923, in1923_1, in1923_2;
    wire c1923;
    assign in1923_1 = {pp34[38]};
    assign in1923_2 = {pp35[37]};
    Full_Adder FA_1923(s1923, c1923, in1923_1, in1923_2, pp33[39]);
    wire[0:0] s1924, in1924_1, in1924_2;
    wire c1924;
    assign in1924_1 = {pp37[35]};
    assign in1924_2 = {pp38[34]};
    Full_Adder FA_1924(s1924, c1924, in1924_1, in1924_2, pp36[36]);
    wire[0:0] s1925, in1925_1, in1925_2;
    wire c1925;
    assign in1925_1 = {pp40[32]};
    assign in1925_2 = {pp41[31]};
    Full_Adder FA_1925(s1925, c1925, in1925_1, in1925_2, pp39[33]);
    wire[0:0] s1926, in1926_1, in1926_2;
    wire c1926;
    assign in1926_1 = {pp42[30]};
    assign in1926_2 = {pp43[29]};
    Half_Adder HA_1926(s1926, c1926, in1926_1, in1926_2);
    wire[0:0] s1927, in1927_1, in1927_2;
    wire c1927;
    assign in1927_1 = {pp1[72]};
    assign in1927_2 = {pp2[71]};
    Full_Adder FA_1927(s1927, c1927, in1927_1, in1927_2, pp0[73]);
    wire[0:0] s1928, in1928_1, in1928_2;
    wire c1928;
    assign in1928_1 = {pp4[69]};
    assign in1928_2 = {pp5[68]};
    Full_Adder FA_1928(s1928, c1928, in1928_1, in1928_2, pp3[70]);
    wire[0:0] s1929, in1929_1, in1929_2;
    wire c1929;
    assign in1929_1 = {pp7[66]};
    assign in1929_2 = {pp8[65]};
    Full_Adder FA_1929(s1929, c1929, in1929_1, in1929_2, pp6[67]);
    wire[0:0] s1930, in1930_1, in1930_2;
    wire c1930;
    assign in1930_1 = {pp10[63]};
    assign in1930_2 = {pp11[62]};
    Full_Adder FA_1930(s1930, c1930, in1930_1, in1930_2, pp9[64]);
    wire[0:0] s1931, in1931_1, in1931_2;
    wire c1931;
    assign in1931_1 = {pp13[60]};
    assign in1931_2 = {pp14[59]};
    Full_Adder FA_1931(s1931, c1931, in1931_1, in1931_2, pp12[61]);
    wire[0:0] s1932, in1932_1, in1932_2;
    wire c1932;
    assign in1932_1 = {pp16[57]};
    assign in1932_2 = {pp17[56]};
    Full_Adder FA_1932(s1932, c1932, in1932_1, in1932_2, pp15[58]);
    wire[0:0] s1933, in1933_1, in1933_2;
    wire c1933;
    assign in1933_1 = {pp19[54]};
    assign in1933_2 = {pp20[53]};
    Full_Adder FA_1933(s1933, c1933, in1933_1, in1933_2, pp18[55]);
    wire[0:0] s1934, in1934_1, in1934_2;
    wire c1934;
    assign in1934_1 = {pp22[51]};
    assign in1934_2 = {pp23[50]};
    Full_Adder FA_1934(s1934, c1934, in1934_1, in1934_2, pp21[52]);
    wire[0:0] s1935, in1935_1, in1935_2;
    wire c1935;
    assign in1935_1 = {pp25[48]};
    assign in1935_2 = {pp26[47]};
    Full_Adder FA_1935(s1935, c1935, in1935_1, in1935_2, pp24[49]);
    wire[0:0] s1936, in1936_1, in1936_2;
    wire c1936;
    assign in1936_1 = {pp28[45]};
    assign in1936_2 = {pp29[44]};
    Full_Adder FA_1936(s1936, c1936, in1936_1, in1936_2, pp27[46]);
    wire[0:0] s1937, in1937_1, in1937_2;
    wire c1937;
    assign in1937_1 = {pp31[42]};
    assign in1937_2 = {pp32[41]};
    Full_Adder FA_1937(s1937, c1937, in1937_1, in1937_2, pp30[43]);
    wire[0:0] s1938, in1938_1, in1938_2;
    wire c1938;
    assign in1938_1 = {pp34[39]};
    assign in1938_2 = {pp35[38]};
    Full_Adder FA_1938(s1938, c1938, in1938_1, in1938_2, pp33[40]);
    wire[0:0] s1939, in1939_1, in1939_2;
    wire c1939;
    assign in1939_1 = {pp37[36]};
    assign in1939_2 = {pp38[35]};
    Full_Adder FA_1939(s1939, c1939, in1939_1, in1939_2, pp36[37]);
    wire[0:0] s1940, in1940_1, in1940_2;
    wire c1940;
    assign in1940_1 = {pp40[33]};
    assign in1940_2 = {pp41[32]};
    Full_Adder FA_1940(s1940, c1940, in1940_1, in1940_2, pp39[34]);
    wire[0:0] s1941, in1941_1, in1941_2;
    wire c1941;
    assign in1941_1 = {pp43[30]};
    assign in1941_2 = {pp44[29]};
    Full_Adder FA_1941(s1941, c1941, in1941_1, in1941_2, pp42[31]);
    wire[0:0] s1942, in1942_1, in1942_2;
    wire c1942;
    assign in1942_1 = {pp45[28]};
    assign in1942_2 = {pp46[27]};
    Half_Adder HA_1942(s1942, c1942, in1942_1, in1942_2);
    wire[0:0] s1943, in1943_1, in1943_2;
    wire c1943;
    assign in1943_1 = {pp1[73]};
    assign in1943_2 = {pp2[72]};
    Full_Adder FA_1943(s1943, c1943, in1943_1, in1943_2, pp0[74]);
    wire[0:0] s1944, in1944_1, in1944_2;
    wire c1944;
    assign in1944_1 = {pp4[70]};
    assign in1944_2 = {pp5[69]};
    Full_Adder FA_1944(s1944, c1944, in1944_1, in1944_2, pp3[71]);
    wire[0:0] s1945, in1945_1, in1945_2;
    wire c1945;
    assign in1945_1 = {pp7[67]};
    assign in1945_2 = {pp8[66]};
    Full_Adder FA_1945(s1945, c1945, in1945_1, in1945_2, pp6[68]);
    wire[0:0] s1946, in1946_1, in1946_2;
    wire c1946;
    assign in1946_1 = {pp10[64]};
    assign in1946_2 = {pp11[63]};
    Full_Adder FA_1946(s1946, c1946, in1946_1, in1946_2, pp9[65]);
    wire[0:0] s1947, in1947_1, in1947_2;
    wire c1947;
    assign in1947_1 = {pp13[61]};
    assign in1947_2 = {pp14[60]};
    Full_Adder FA_1947(s1947, c1947, in1947_1, in1947_2, pp12[62]);
    wire[0:0] s1948, in1948_1, in1948_2;
    wire c1948;
    assign in1948_1 = {pp16[58]};
    assign in1948_2 = {pp17[57]};
    Full_Adder FA_1948(s1948, c1948, in1948_1, in1948_2, pp15[59]);
    wire[0:0] s1949, in1949_1, in1949_2;
    wire c1949;
    assign in1949_1 = {pp19[55]};
    assign in1949_2 = {pp20[54]};
    Full_Adder FA_1949(s1949, c1949, in1949_1, in1949_2, pp18[56]);
    wire[0:0] s1950, in1950_1, in1950_2;
    wire c1950;
    assign in1950_1 = {pp22[52]};
    assign in1950_2 = {pp23[51]};
    Full_Adder FA_1950(s1950, c1950, in1950_1, in1950_2, pp21[53]);
    wire[0:0] s1951, in1951_1, in1951_2;
    wire c1951;
    assign in1951_1 = {pp25[49]};
    assign in1951_2 = {pp26[48]};
    Full_Adder FA_1951(s1951, c1951, in1951_1, in1951_2, pp24[50]);
    wire[0:0] s1952, in1952_1, in1952_2;
    wire c1952;
    assign in1952_1 = {pp28[46]};
    assign in1952_2 = {pp29[45]};
    Full_Adder FA_1952(s1952, c1952, in1952_1, in1952_2, pp27[47]);
    wire[0:0] s1953, in1953_1, in1953_2;
    wire c1953;
    assign in1953_1 = {pp31[43]};
    assign in1953_2 = {pp32[42]};
    Full_Adder FA_1953(s1953, c1953, in1953_1, in1953_2, pp30[44]);
    wire[0:0] s1954, in1954_1, in1954_2;
    wire c1954;
    assign in1954_1 = {pp34[40]};
    assign in1954_2 = {pp35[39]};
    Full_Adder FA_1954(s1954, c1954, in1954_1, in1954_2, pp33[41]);
    wire[0:0] s1955, in1955_1, in1955_2;
    wire c1955;
    assign in1955_1 = {pp37[37]};
    assign in1955_2 = {pp38[36]};
    Full_Adder FA_1955(s1955, c1955, in1955_1, in1955_2, pp36[38]);
    wire[0:0] s1956, in1956_1, in1956_2;
    wire c1956;
    assign in1956_1 = {pp40[34]};
    assign in1956_2 = {pp41[33]};
    Full_Adder FA_1956(s1956, c1956, in1956_1, in1956_2, pp39[35]);
    wire[0:0] s1957, in1957_1, in1957_2;
    wire c1957;
    assign in1957_1 = {pp43[31]};
    assign in1957_2 = {pp44[30]};
    Full_Adder FA_1957(s1957, c1957, in1957_1, in1957_2, pp42[32]);
    wire[0:0] s1958, in1958_1, in1958_2;
    wire c1958;
    assign in1958_1 = {pp46[28]};
    assign in1958_2 = {pp47[27]};
    Full_Adder FA_1958(s1958, c1958, in1958_1, in1958_2, pp45[29]);
    wire[0:0] s1959, in1959_1, in1959_2;
    wire c1959;
    assign in1959_1 = {pp48[26]};
    assign in1959_2 = {pp49[25]};
    Half_Adder HA_1959(s1959, c1959, in1959_1, in1959_2);
    wire[0:0] s1960, in1960_1, in1960_2;
    wire c1960;
    assign in1960_1 = {pp1[74]};
    assign in1960_2 = {pp2[73]};
    Full_Adder FA_1960(s1960, c1960, in1960_1, in1960_2, pp0[75]);
    wire[0:0] s1961, in1961_1, in1961_2;
    wire c1961;
    assign in1961_1 = {pp4[71]};
    assign in1961_2 = {pp5[70]};
    Full_Adder FA_1961(s1961, c1961, in1961_1, in1961_2, pp3[72]);
    wire[0:0] s1962, in1962_1, in1962_2;
    wire c1962;
    assign in1962_1 = {pp7[68]};
    assign in1962_2 = {pp8[67]};
    Full_Adder FA_1962(s1962, c1962, in1962_1, in1962_2, pp6[69]);
    wire[0:0] s1963, in1963_1, in1963_2;
    wire c1963;
    assign in1963_1 = {pp10[65]};
    assign in1963_2 = {pp11[64]};
    Full_Adder FA_1963(s1963, c1963, in1963_1, in1963_2, pp9[66]);
    wire[0:0] s1964, in1964_1, in1964_2;
    wire c1964;
    assign in1964_1 = {pp13[62]};
    assign in1964_2 = {pp14[61]};
    Full_Adder FA_1964(s1964, c1964, in1964_1, in1964_2, pp12[63]);
    wire[0:0] s1965, in1965_1, in1965_2;
    wire c1965;
    assign in1965_1 = {pp16[59]};
    assign in1965_2 = {pp17[58]};
    Full_Adder FA_1965(s1965, c1965, in1965_1, in1965_2, pp15[60]);
    wire[0:0] s1966, in1966_1, in1966_2;
    wire c1966;
    assign in1966_1 = {pp19[56]};
    assign in1966_2 = {pp20[55]};
    Full_Adder FA_1966(s1966, c1966, in1966_1, in1966_2, pp18[57]);
    wire[0:0] s1967, in1967_1, in1967_2;
    wire c1967;
    assign in1967_1 = {pp22[53]};
    assign in1967_2 = {pp23[52]};
    Full_Adder FA_1967(s1967, c1967, in1967_1, in1967_2, pp21[54]);
    wire[0:0] s1968, in1968_1, in1968_2;
    wire c1968;
    assign in1968_1 = {pp25[50]};
    assign in1968_2 = {pp26[49]};
    Full_Adder FA_1968(s1968, c1968, in1968_1, in1968_2, pp24[51]);
    wire[0:0] s1969, in1969_1, in1969_2;
    wire c1969;
    assign in1969_1 = {pp28[47]};
    assign in1969_2 = {pp29[46]};
    Full_Adder FA_1969(s1969, c1969, in1969_1, in1969_2, pp27[48]);
    wire[0:0] s1970, in1970_1, in1970_2;
    wire c1970;
    assign in1970_1 = {pp31[44]};
    assign in1970_2 = {pp32[43]};
    Full_Adder FA_1970(s1970, c1970, in1970_1, in1970_2, pp30[45]);
    wire[0:0] s1971, in1971_1, in1971_2;
    wire c1971;
    assign in1971_1 = {pp34[41]};
    assign in1971_2 = {pp35[40]};
    Full_Adder FA_1971(s1971, c1971, in1971_1, in1971_2, pp33[42]);
    wire[0:0] s1972, in1972_1, in1972_2;
    wire c1972;
    assign in1972_1 = {pp37[38]};
    assign in1972_2 = {pp38[37]};
    Full_Adder FA_1972(s1972, c1972, in1972_1, in1972_2, pp36[39]);
    wire[0:0] s1973, in1973_1, in1973_2;
    wire c1973;
    assign in1973_1 = {pp40[35]};
    assign in1973_2 = {pp41[34]};
    Full_Adder FA_1973(s1973, c1973, in1973_1, in1973_2, pp39[36]);
    wire[0:0] s1974, in1974_1, in1974_2;
    wire c1974;
    assign in1974_1 = {pp43[32]};
    assign in1974_2 = {pp44[31]};
    Full_Adder FA_1974(s1974, c1974, in1974_1, in1974_2, pp42[33]);
    wire[0:0] s1975, in1975_1, in1975_2;
    wire c1975;
    assign in1975_1 = {pp46[29]};
    assign in1975_2 = {pp47[28]};
    Full_Adder FA_1975(s1975, c1975, in1975_1, in1975_2, pp45[30]);
    wire[0:0] s1976, in1976_1, in1976_2;
    wire c1976;
    assign in1976_1 = {pp49[26]};
    assign in1976_2 = {pp50[25]};
    Full_Adder FA_1976(s1976, c1976, in1976_1, in1976_2, pp48[27]);
    wire[0:0] s1977, in1977_1, in1977_2;
    wire c1977;
    assign in1977_1 = {pp51[24]};
    assign in1977_2 = {pp52[23]};
    Half_Adder HA_1977(s1977, c1977, in1977_1, in1977_2);
    wire[0:0] s1978, in1978_1, in1978_2;
    wire c1978;
    assign in1978_1 = {pp1[75]};
    assign in1978_2 = {pp2[74]};
    Full_Adder FA_1978(s1978, c1978, in1978_1, in1978_2, pp0[76]);
    wire[0:0] s1979, in1979_1, in1979_2;
    wire c1979;
    assign in1979_1 = {pp4[72]};
    assign in1979_2 = {pp5[71]};
    Full_Adder FA_1979(s1979, c1979, in1979_1, in1979_2, pp3[73]);
    wire[0:0] s1980, in1980_1, in1980_2;
    wire c1980;
    assign in1980_1 = {pp7[69]};
    assign in1980_2 = {pp8[68]};
    Full_Adder FA_1980(s1980, c1980, in1980_1, in1980_2, pp6[70]);
    wire[0:0] s1981, in1981_1, in1981_2;
    wire c1981;
    assign in1981_1 = {pp10[66]};
    assign in1981_2 = {pp11[65]};
    Full_Adder FA_1981(s1981, c1981, in1981_1, in1981_2, pp9[67]);
    wire[0:0] s1982, in1982_1, in1982_2;
    wire c1982;
    assign in1982_1 = {pp13[63]};
    assign in1982_2 = {pp14[62]};
    Full_Adder FA_1982(s1982, c1982, in1982_1, in1982_2, pp12[64]);
    wire[0:0] s1983, in1983_1, in1983_2;
    wire c1983;
    assign in1983_1 = {pp16[60]};
    assign in1983_2 = {pp17[59]};
    Full_Adder FA_1983(s1983, c1983, in1983_1, in1983_2, pp15[61]);
    wire[0:0] s1984, in1984_1, in1984_2;
    wire c1984;
    assign in1984_1 = {pp19[57]};
    assign in1984_2 = {pp20[56]};
    Full_Adder FA_1984(s1984, c1984, in1984_1, in1984_2, pp18[58]);
    wire[0:0] s1985, in1985_1, in1985_2;
    wire c1985;
    assign in1985_1 = {pp22[54]};
    assign in1985_2 = {pp23[53]};
    Full_Adder FA_1985(s1985, c1985, in1985_1, in1985_2, pp21[55]);
    wire[0:0] s1986, in1986_1, in1986_2;
    wire c1986;
    assign in1986_1 = {pp25[51]};
    assign in1986_2 = {pp26[50]};
    Full_Adder FA_1986(s1986, c1986, in1986_1, in1986_2, pp24[52]);
    wire[0:0] s1987, in1987_1, in1987_2;
    wire c1987;
    assign in1987_1 = {pp28[48]};
    assign in1987_2 = {pp29[47]};
    Full_Adder FA_1987(s1987, c1987, in1987_1, in1987_2, pp27[49]);
    wire[0:0] s1988, in1988_1, in1988_2;
    wire c1988;
    assign in1988_1 = {pp31[45]};
    assign in1988_2 = {pp32[44]};
    Full_Adder FA_1988(s1988, c1988, in1988_1, in1988_2, pp30[46]);
    wire[0:0] s1989, in1989_1, in1989_2;
    wire c1989;
    assign in1989_1 = {pp34[42]};
    assign in1989_2 = {pp35[41]};
    Full_Adder FA_1989(s1989, c1989, in1989_1, in1989_2, pp33[43]);
    wire[0:0] s1990, in1990_1, in1990_2;
    wire c1990;
    assign in1990_1 = {pp37[39]};
    assign in1990_2 = {pp38[38]};
    Full_Adder FA_1990(s1990, c1990, in1990_1, in1990_2, pp36[40]);
    wire[0:0] s1991, in1991_1, in1991_2;
    wire c1991;
    assign in1991_1 = {pp40[36]};
    assign in1991_2 = {pp41[35]};
    Full_Adder FA_1991(s1991, c1991, in1991_1, in1991_2, pp39[37]);
    wire[0:0] s1992, in1992_1, in1992_2;
    wire c1992;
    assign in1992_1 = {pp43[33]};
    assign in1992_2 = {pp44[32]};
    Full_Adder FA_1992(s1992, c1992, in1992_1, in1992_2, pp42[34]);
    wire[0:0] s1993, in1993_1, in1993_2;
    wire c1993;
    assign in1993_1 = {pp46[30]};
    assign in1993_2 = {pp47[29]};
    Full_Adder FA_1993(s1993, c1993, in1993_1, in1993_2, pp45[31]);
    wire[0:0] s1994, in1994_1, in1994_2;
    wire c1994;
    assign in1994_1 = {pp49[27]};
    assign in1994_2 = {pp50[26]};
    Full_Adder FA_1994(s1994, c1994, in1994_1, in1994_2, pp48[28]);
    wire[0:0] s1995, in1995_1, in1995_2;
    wire c1995;
    assign in1995_1 = {pp52[24]};
    assign in1995_2 = {pp53[23]};
    Full_Adder FA_1995(s1995, c1995, in1995_1, in1995_2, pp51[25]);
    wire[0:0] s1996, in1996_1, in1996_2;
    wire c1996;
    assign in1996_1 = {pp54[22]};
    assign in1996_2 = {pp55[21]};
    Half_Adder HA_1996(s1996, c1996, in1996_1, in1996_2);
    wire[0:0] s1997, in1997_1, in1997_2;
    wire c1997;
    assign in1997_1 = {pp1[76]};
    assign in1997_2 = {pp2[75]};
    Full_Adder FA_1997(s1997, c1997, in1997_1, in1997_2, pp0[77]);
    wire[0:0] s1998, in1998_1, in1998_2;
    wire c1998;
    assign in1998_1 = {pp4[73]};
    assign in1998_2 = {pp5[72]};
    Full_Adder FA_1998(s1998, c1998, in1998_1, in1998_2, pp3[74]);
    wire[0:0] s1999, in1999_1, in1999_2;
    wire c1999;
    assign in1999_1 = {pp7[70]};
    assign in1999_2 = {pp8[69]};
    Full_Adder FA_1999(s1999, c1999, in1999_1, in1999_2, pp6[71]);
    wire[0:0] s2000, in2000_1, in2000_2;
    wire c2000;
    assign in2000_1 = {pp10[67]};
    assign in2000_2 = {pp11[66]};
    Full_Adder FA_2000(s2000, c2000, in2000_1, in2000_2, pp9[68]);
    wire[0:0] s2001, in2001_1, in2001_2;
    wire c2001;
    assign in2001_1 = {pp13[64]};
    assign in2001_2 = {pp14[63]};
    Full_Adder FA_2001(s2001, c2001, in2001_1, in2001_2, pp12[65]);
    wire[0:0] s2002, in2002_1, in2002_2;
    wire c2002;
    assign in2002_1 = {pp16[61]};
    assign in2002_2 = {pp17[60]};
    Full_Adder FA_2002(s2002, c2002, in2002_1, in2002_2, pp15[62]);
    wire[0:0] s2003, in2003_1, in2003_2;
    wire c2003;
    assign in2003_1 = {pp19[58]};
    assign in2003_2 = {pp20[57]};
    Full_Adder FA_2003(s2003, c2003, in2003_1, in2003_2, pp18[59]);
    wire[0:0] s2004, in2004_1, in2004_2;
    wire c2004;
    assign in2004_1 = {pp22[55]};
    assign in2004_2 = {pp23[54]};
    Full_Adder FA_2004(s2004, c2004, in2004_1, in2004_2, pp21[56]);
    wire[0:0] s2005, in2005_1, in2005_2;
    wire c2005;
    assign in2005_1 = {pp25[52]};
    assign in2005_2 = {pp26[51]};
    Full_Adder FA_2005(s2005, c2005, in2005_1, in2005_2, pp24[53]);
    wire[0:0] s2006, in2006_1, in2006_2;
    wire c2006;
    assign in2006_1 = {pp28[49]};
    assign in2006_2 = {pp29[48]};
    Full_Adder FA_2006(s2006, c2006, in2006_1, in2006_2, pp27[50]);
    wire[0:0] s2007, in2007_1, in2007_2;
    wire c2007;
    assign in2007_1 = {pp31[46]};
    assign in2007_2 = {pp32[45]};
    Full_Adder FA_2007(s2007, c2007, in2007_1, in2007_2, pp30[47]);
    wire[0:0] s2008, in2008_1, in2008_2;
    wire c2008;
    assign in2008_1 = {pp34[43]};
    assign in2008_2 = {pp35[42]};
    Full_Adder FA_2008(s2008, c2008, in2008_1, in2008_2, pp33[44]);
    wire[0:0] s2009, in2009_1, in2009_2;
    wire c2009;
    assign in2009_1 = {pp37[40]};
    assign in2009_2 = {pp38[39]};
    Full_Adder FA_2009(s2009, c2009, in2009_1, in2009_2, pp36[41]);
    wire[0:0] s2010, in2010_1, in2010_2;
    wire c2010;
    assign in2010_1 = {pp40[37]};
    assign in2010_2 = {pp41[36]};
    Full_Adder FA_2010(s2010, c2010, in2010_1, in2010_2, pp39[38]);
    wire[0:0] s2011, in2011_1, in2011_2;
    wire c2011;
    assign in2011_1 = {pp43[34]};
    assign in2011_2 = {pp44[33]};
    Full_Adder FA_2011(s2011, c2011, in2011_1, in2011_2, pp42[35]);
    wire[0:0] s2012, in2012_1, in2012_2;
    wire c2012;
    assign in2012_1 = {pp46[31]};
    assign in2012_2 = {pp47[30]};
    Full_Adder FA_2012(s2012, c2012, in2012_1, in2012_2, pp45[32]);
    wire[0:0] s2013, in2013_1, in2013_2;
    wire c2013;
    assign in2013_1 = {pp49[28]};
    assign in2013_2 = {pp50[27]};
    Full_Adder FA_2013(s2013, c2013, in2013_1, in2013_2, pp48[29]);
    wire[0:0] s2014, in2014_1, in2014_2;
    wire c2014;
    assign in2014_1 = {pp52[25]};
    assign in2014_2 = {pp53[24]};
    Full_Adder FA_2014(s2014, c2014, in2014_1, in2014_2, pp51[26]);
    wire[0:0] s2015, in2015_1, in2015_2;
    wire c2015;
    assign in2015_1 = {pp55[22]};
    assign in2015_2 = {pp56[21]};
    Full_Adder FA_2015(s2015, c2015, in2015_1, in2015_2, pp54[23]);
    wire[0:0] s2016, in2016_1, in2016_2;
    wire c2016;
    assign in2016_1 = {pp57[20]};
    assign in2016_2 = {pp58[19]};
    Half_Adder HA_2016(s2016, c2016, in2016_1, in2016_2);
    wire[0:0] s2017, in2017_1, in2017_2;
    wire c2017;
    assign in2017_1 = {pp1[77]};
    assign in2017_2 = {pp2[76]};
    Full_Adder FA_2017(s2017, c2017, in2017_1, in2017_2, pp0[78]);
    wire[0:0] s2018, in2018_1, in2018_2;
    wire c2018;
    assign in2018_1 = {pp4[74]};
    assign in2018_2 = {pp5[73]};
    Full_Adder FA_2018(s2018, c2018, in2018_1, in2018_2, pp3[75]);
    wire[0:0] s2019, in2019_1, in2019_2;
    wire c2019;
    assign in2019_1 = {pp7[71]};
    assign in2019_2 = {pp8[70]};
    Full_Adder FA_2019(s2019, c2019, in2019_1, in2019_2, pp6[72]);
    wire[0:0] s2020, in2020_1, in2020_2;
    wire c2020;
    assign in2020_1 = {pp10[68]};
    assign in2020_2 = {pp11[67]};
    Full_Adder FA_2020(s2020, c2020, in2020_1, in2020_2, pp9[69]);
    wire[0:0] s2021, in2021_1, in2021_2;
    wire c2021;
    assign in2021_1 = {pp13[65]};
    assign in2021_2 = {pp14[64]};
    Full_Adder FA_2021(s2021, c2021, in2021_1, in2021_2, pp12[66]);
    wire[0:0] s2022, in2022_1, in2022_2;
    wire c2022;
    assign in2022_1 = {pp16[62]};
    assign in2022_2 = {pp17[61]};
    Full_Adder FA_2022(s2022, c2022, in2022_1, in2022_2, pp15[63]);
    wire[0:0] s2023, in2023_1, in2023_2;
    wire c2023;
    assign in2023_1 = {pp19[59]};
    assign in2023_2 = {pp20[58]};
    Full_Adder FA_2023(s2023, c2023, in2023_1, in2023_2, pp18[60]);
    wire[0:0] s2024, in2024_1, in2024_2;
    wire c2024;
    assign in2024_1 = {pp22[56]};
    assign in2024_2 = {pp23[55]};
    Full_Adder FA_2024(s2024, c2024, in2024_1, in2024_2, pp21[57]);
    wire[0:0] s2025, in2025_1, in2025_2;
    wire c2025;
    assign in2025_1 = {pp25[53]};
    assign in2025_2 = {pp26[52]};
    Full_Adder FA_2025(s2025, c2025, in2025_1, in2025_2, pp24[54]);
    wire[0:0] s2026, in2026_1, in2026_2;
    wire c2026;
    assign in2026_1 = {pp28[50]};
    assign in2026_2 = {pp29[49]};
    Full_Adder FA_2026(s2026, c2026, in2026_1, in2026_2, pp27[51]);
    wire[0:0] s2027, in2027_1, in2027_2;
    wire c2027;
    assign in2027_1 = {pp31[47]};
    assign in2027_2 = {pp32[46]};
    Full_Adder FA_2027(s2027, c2027, in2027_1, in2027_2, pp30[48]);
    wire[0:0] s2028, in2028_1, in2028_2;
    wire c2028;
    assign in2028_1 = {pp34[44]};
    assign in2028_2 = {pp35[43]};
    Full_Adder FA_2028(s2028, c2028, in2028_1, in2028_2, pp33[45]);
    wire[0:0] s2029, in2029_1, in2029_2;
    wire c2029;
    assign in2029_1 = {pp37[41]};
    assign in2029_2 = {pp38[40]};
    Full_Adder FA_2029(s2029, c2029, in2029_1, in2029_2, pp36[42]);
    wire[0:0] s2030, in2030_1, in2030_2;
    wire c2030;
    assign in2030_1 = {pp40[38]};
    assign in2030_2 = {pp41[37]};
    Full_Adder FA_2030(s2030, c2030, in2030_1, in2030_2, pp39[39]);
    wire[0:0] s2031, in2031_1, in2031_2;
    wire c2031;
    assign in2031_1 = {pp43[35]};
    assign in2031_2 = {pp44[34]};
    Full_Adder FA_2031(s2031, c2031, in2031_1, in2031_2, pp42[36]);
    wire[0:0] s2032, in2032_1, in2032_2;
    wire c2032;
    assign in2032_1 = {pp46[32]};
    assign in2032_2 = {pp47[31]};
    Full_Adder FA_2032(s2032, c2032, in2032_1, in2032_2, pp45[33]);
    wire[0:0] s2033, in2033_1, in2033_2;
    wire c2033;
    assign in2033_1 = {pp49[29]};
    assign in2033_2 = {pp50[28]};
    Full_Adder FA_2033(s2033, c2033, in2033_1, in2033_2, pp48[30]);
    wire[0:0] s2034, in2034_1, in2034_2;
    wire c2034;
    assign in2034_1 = {pp52[26]};
    assign in2034_2 = {pp53[25]};
    Full_Adder FA_2034(s2034, c2034, in2034_1, in2034_2, pp51[27]);
    wire[0:0] s2035, in2035_1, in2035_2;
    wire c2035;
    assign in2035_1 = {pp55[23]};
    assign in2035_2 = {pp56[22]};
    Full_Adder FA_2035(s2035, c2035, in2035_1, in2035_2, pp54[24]);
    wire[0:0] s2036, in2036_1, in2036_2;
    wire c2036;
    assign in2036_1 = {pp58[20]};
    assign in2036_2 = {pp59[19]};
    Full_Adder FA_2036(s2036, c2036, in2036_1, in2036_2, pp57[21]);
    wire[0:0] s2037, in2037_1, in2037_2;
    wire c2037;
    assign in2037_1 = {pp60[18]};
    assign in2037_2 = {pp61[17]};
    Half_Adder HA_2037(s2037, c2037, in2037_1, in2037_2);
    wire[0:0] s2038, in2038_1, in2038_2;
    wire c2038;
    assign in2038_1 = {pp1[78]};
    assign in2038_2 = {pp2[77]};
    Full_Adder FA_2038(s2038, c2038, in2038_1, in2038_2, pp0[79]);
    wire[0:0] s2039, in2039_1, in2039_2;
    wire c2039;
    assign in2039_1 = {pp4[75]};
    assign in2039_2 = {pp5[74]};
    Full_Adder FA_2039(s2039, c2039, in2039_1, in2039_2, pp3[76]);
    wire[0:0] s2040, in2040_1, in2040_2;
    wire c2040;
    assign in2040_1 = {pp7[72]};
    assign in2040_2 = {pp8[71]};
    Full_Adder FA_2040(s2040, c2040, in2040_1, in2040_2, pp6[73]);
    wire[0:0] s2041, in2041_1, in2041_2;
    wire c2041;
    assign in2041_1 = {pp10[69]};
    assign in2041_2 = {pp11[68]};
    Full_Adder FA_2041(s2041, c2041, in2041_1, in2041_2, pp9[70]);
    wire[0:0] s2042, in2042_1, in2042_2;
    wire c2042;
    assign in2042_1 = {pp13[66]};
    assign in2042_2 = {pp14[65]};
    Full_Adder FA_2042(s2042, c2042, in2042_1, in2042_2, pp12[67]);
    wire[0:0] s2043, in2043_1, in2043_2;
    wire c2043;
    assign in2043_1 = {pp16[63]};
    assign in2043_2 = {pp17[62]};
    Full_Adder FA_2043(s2043, c2043, in2043_1, in2043_2, pp15[64]);
    wire[0:0] s2044, in2044_1, in2044_2;
    wire c2044;
    assign in2044_1 = {pp19[60]};
    assign in2044_2 = {pp20[59]};
    Full_Adder FA_2044(s2044, c2044, in2044_1, in2044_2, pp18[61]);
    wire[0:0] s2045, in2045_1, in2045_2;
    wire c2045;
    assign in2045_1 = {pp22[57]};
    assign in2045_2 = {pp23[56]};
    Full_Adder FA_2045(s2045, c2045, in2045_1, in2045_2, pp21[58]);
    wire[0:0] s2046, in2046_1, in2046_2;
    wire c2046;
    assign in2046_1 = {pp25[54]};
    assign in2046_2 = {pp26[53]};
    Full_Adder FA_2046(s2046, c2046, in2046_1, in2046_2, pp24[55]);
    wire[0:0] s2047, in2047_1, in2047_2;
    wire c2047;
    assign in2047_1 = {pp28[51]};
    assign in2047_2 = {pp29[50]};
    Full_Adder FA_2047(s2047, c2047, in2047_1, in2047_2, pp27[52]);
    wire[0:0] s2048, in2048_1, in2048_2;
    wire c2048;
    assign in2048_1 = {pp31[48]};
    assign in2048_2 = {pp32[47]};
    Full_Adder FA_2048(s2048, c2048, in2048_1, in2048_2, pp30[49]);
    wire[0:0] s2049, in2049_1, in2049_2;
    wire c2049;
    assign in2049_1 = {pp34[45]};
    assign in2049_2 = {pp35[44]};
    Full_Adder FA_2049(s2049, c2049, in2049_1, in2049_2, pp33[46]);
    wire[0:0] s2050, in2050_1, in2050_2;
    wire c2050;
    assign in2050_1 = {pp37[42]};
    assign in2050_2 = {pp38[41]};
    Full_Adder FA_2050(s2050, c2050, in2050_1, in2050_2, pp36[43]);
    wire[0:0] s2051, in2051_1, in2051_2;
    wire c2051;
    assign in2051_1 = {pp40[39]};
    assign in2051_2 = {pp41[38]};
    Full_Adder FA_2051(s2051, c2051, in2051_1, in2051_2, pp39[40]);
    wire[0:0] s2052, in2052_1, in2052_2;
    wire c2052;
    assign in2052_1 = {pp43[36]};
    assign in2052_2 = {pp44[35]};
    Full_Adder FA_2052(s2052, c2052, in2052_1, in2052_2, pp42[37]);
    wire[0:0] s2053, in2053_1, in2053_2;
    wire c2053;
    assign in2053_1 = {pp46[33]};
    assign in2053_2 = {pp47[32]};
    Full_Adder FA_2053(s2053, c2053, in2053_1, in2053_2, pp45[34]);
    wire[0:0] s2054, in2054_1, in2054_2;
    wire c2054;
    assign in2054_1 = {pp49[30]};
    assign in2054_2 = {pp50[29]};
    Full_Adder FA_2054(s2054, c2054, in2054_1, in2054_2, pp48[31]);
    wire[0:0] s2055, in2055_1, in2055_2;
    wire c2055;
    assign in2055_1 = {pp52[27]};
    assign in2055_2 = {pp53[26]};
    Full_Adder FA_2055(s2055, c2055, in2055_1, in2055_2, pp51[28]);
    wire[0:0] s2056, in2056_1, in2056_2;
    wire c2056;
    assign in2056_1 = {pp55[24]};
    assign in2056_2 = {pp56[23]};
    Full_Adder FA_2056(s2056, c2056, in2056_1, in2056_2, pp54[25]);
    wire[0:0] s2057, in2057_1, in2057_2;
    wire c2057;
    assign in2057_1 = {pp58[21]};
    assign in2057_2 = {pp59[20]};
    Full_Adder FA_2057(s2057, c2057, in2057_1, in2057_2, pp57[22]);
    wire[0:0] s2058, in2058_1, in2058_2;
    wire c2058;
    assign in2058_1 = {pp61[18]};
    assign in2058_2 = {pp62[17]};
    Full_Adder FA_2058(s2058, c2058, in2058_1, in2058_2, pp60[19]);
    wire[0:0] s2059, in2059_1, in2059_2;
    wire c2059;
    assign in2059_1 = {pp63[16]};
    assign in2059_2 = {pp64[15]};
    Half_Adder HA_2059(s2059, c2059, in2059_1, in2059_2);
    wire[0:0] s2060, in2060_1, in2060_2;
    wire c2060;
    assign in2060_1 = {pp1[79]};
    assign in2060_2 = {pp2[78]};
    Full_Adder FA_2060(s2060, c2060, in2060_1, in2060_2, pp0[80]);
    wire[0:0] s2061, in2061_1, in2061_2;
    wire c2061;
    assign in2061_1 = {pp4[76]};
    assign in2061_2 = {pp5[75]};
    Full_Adder FA_2061(s2061, c2061, in2061_1, in2061_2, pp3[77]);
    wire[0:0] s2062, in2062_1, in2062_2;
    wire c2062;
    assign in2062_1 = {pp7[73]};
    assign in2062_2 = {pp8[72]};
    Full_Adder FA_2062(s2062, c2062, in2062_1, in2062_2, pp6[74]);
    wire[0:0] s2063, in2063_1, in2063_2;
    wire c2063;
    assign in2063_1 = {pp10[70]};
    assign in2063_2 = {pp11[69]};
    Full_Adder FA_2063(s2063, c2063, in2063_1, in2063_2, pp9[71]);
    wire[0:0] s2064, in2064_1, in2064_2;
    wire c2064;
    assign in2064_1 = {pp13[67]};
    assign in2064_2 = {pp14[66]};
    Full_Adder FA_2064(s2064, c2064, in2064_1, in2064_2, pp12[68]);
    wire[0:0] s2065, in2065_1, in2065_2;
    wire c2065;
    assign in2065_1 = {pp16[64]};
    assign in2065_2 = {pp17[63]};
    Full_Adder FA_2065(s2065, c2065, in2065_1, in2065_2, pp15[65]);
    wire[0:0] s2066, in2066_1, in2066_2;
    wire c2066;
    assign in2066_1 = {pp19[61]};
    assign in2066_2 = {pp20[60]};
    Full_Adder FA_2066(s2066, c2066, in2066_1, in2066_2, pp18[62]);
    wire[0:0] s2067, in2067_1, in2067_2;
    wire c2067;
    assign in2067_1 = {pp22[58]};
    assign in2067_2 = {pp23[57]};
    Full_Adder FA_2067(s2067, c2067, in2067_1, in2067_2, pp21[59]);
    wire[0:0] s2068, in2068_1, in2068_2;
    wire c2068;
    assign in2068_1 = {pp25[55]};
    assign in2068_2 = {pp26[54]};
    Full_Adder FA_2068(s2068, c2068, in2068_1, in2068_2, pp24[56]);
    wire[0:0] s2069, in2069_1, in2069_2;
    wire c2069;
    assign in2069_1 = {pp28[52]};
    assign in2069_2 = {pp29[51]};
    Full_Adder FA_2069(s2069, c2069, in2069_1, in2069_2, pp27[53]);
    wire[0:0] s2070, in2070_1, in2070_2;
    wire c2070;
    assign in2070_1 = {pp31[49]};
    assign in2070_2 = {pp32[48]};
    Full_Adder FA_2070(s2070, c2070, in2070_1, in2070_2, pp30[50]);
    wire[0:0] s2071, in2071_1, in2071_2;
    wire c2071;
    assign in2071_1 = {pp34[46]};
    assign in2071_2 = {pp35[45]};
    Full_Adder FA_2071(s2071, c2071, in2071_1, in2071_2, pp33[47]);
    wire[0:0] s2072, in2072_1, in2072_2;
    wire c2072;
    assign in2072_1 = {pp37[43]};
    assign in2072_2 = {pp38[42]};
    Full_Adder FA_2072(s2072, c2072, in2072_1, in2072_2, pp36[44]);
    wire[0:0] s2073, in2073_1, in2073_2;
    wire c2073;
    assign in2073_1 = {pp40[40]};
    assign in2073_2 = {pp41[39]};
    Full_Adder FA_2073(s2073, c2073, in2073_1, in2073_2, pp39[41]);
    wire[0:0] s2074, in2074_1, in2074_2;
    wire c2074;
    assign in2074_1 = {pp43[37]};
    assign in2074_2 = {pp44[36]};
    Full_Adder FA_2074(s2074, c2074, in2074_1, in2074_2, pp42[38]);
    wire[0:0] s2075, in2075_1, in2075_2;
    wire c2075;
    assign in2075_1 = {pp46[34]};
    assign in2075_2 = {pp47[33]};
    Full_Adder FA_2075(s2075, c2075, in2075_1, in2075_2, pp45[35]);
    wire[0:0] s2076, in2076_1, in2076_2;
    wire c2076;
    assign in2076_1 = {pp49[31]};
    assign in2076_2 = {pp50[30]};
    Full_Adder FA_2076(s2076, c2076, in2076_1, in2076_2, pp48[32]);
    wire[0:0] s2077, in2077_1, in2077_2;
    wire c2077;
    assign in2077_1 = {pp52[28]};
    assign in2077_2 = {pp53[27]};
    Full_Adder FA_2077(s2077, c2077, in2077_1, in2077_2, pp51[29]);
    wire[0:0] s2078, in2078_1, in2078_2;
    wire c2078;
    assign in2078_1 = {pp55[25]};
    assign in2078_2 = {pp56[24]};
    Full_Adder FA_2078(s2078, c2078, in2078_1, in2078_2, pp54[26]);
    wire[0:0] s2079, in2079_1, in2079_2;
    wire c2079;
    assign in2079_1 = {pp58[22]};
    assign in2079_2 = {pp59[21]};
    Full_Adder FA_2079(s2079, c2079, in2079_1, in2079_2, pp57[23]);
    wire[0:0] s2080, in2080_1, in2080_2;
    wire c2080;
    assign in2080_1 = {pp61[19]};
    assign in2080_2 = {pp62[18]};
    Full_Adder FA_2080(s2080, c2080, in2080_1, in2080_2, pp60[20]);
    wire[0:0] s2081, in2081_1, in2081_2;
    wire c2081;
    assign in2081_1 = {pp64[16]};
    assign in2081_2 = {pp65[15]};
    Full_Adder FA_2081(s2081, c2081, in2081_1, in2081_2, pp63[17]);
    wire[0:0] s2082, in2082_1, in2082_2;
    wire c2082;
    assign in2082_1 = {pp66[14]};
    assign in2082_2 = {pp67[13]};
    Half_Adder HA_2082(s2082, c2082, in2082_1, in2082_2);
    wire[0:0] s2083, in2083_1, in2083_2;
    wire c2083;
    assign in2083_1 = {pp1[80]};
    assign in2083_2 = {pp2[79]};
    Full_Adder FA_2083(s2083, c2083, in2083_1, in2083_2, pp0[81]);
    wire[0:0] s2084, in2084_1, in2084_2;
    wire c2084;
    assign in2084_1 = {pp4[77]};
    assign in2084_2 = {pp5[76]};
    Full_Adder FA_2084(s2084, c2084, in2084_1, in2084_2, pp3[78]);
    wire[0:0] s2085, in2085_1, in2085_2;
    wire c2085;
    assign in2085_1 = {pp7[74]};
    assign in2085_2 = {pp8[73]};
    Full_Adder FA_2085(s2085, c2085, in2085_1, in2085_2, pp6[75]);
    wire[0:0] s2086, in2086_1, in2086_2;
    wire c2086;
    assign in2086_1 = {pp10[71]};
    assign in2086_2 = {pp11[70]};
    Full_Adder FA_2086(s2086, c2086, in2086_1, in2086_2, pp9[72]);
    wire[0:0] s2087, in2087_1, in2087_2;
    wire c2087;
    assign in2087_1 = {pp13[68]};
    assign in2087_2 = {pp14[67]};
    Full_Adder FA_2087(s2087, c2087, in2087_1, in2087_2, pp12[69]);
    wire[0:0] s2088, in2088_1, in2088_2;
    wire c2088;
    assign in2088_1 = {pp16[65]};
    assign in2088_2 = {pp17[64]};
    Full_Adder FA_2088(s2088, c2088, in2088_1, in2088_2, pp15[66]);
    wire[0:0] s2089, in2089_1, in2089_2;
    wire c2089;
    assign in2089_1 = {pp19[62]};
    assign in2089_2 = {pp20[61]};
    Full_Adder FA_2089(s2089, c2089, in2089_1, in2089_2, pp18[63]);
    wire[0:0] s2090, in2090_1, in2090_2;
    wire c2090;
    assign in2090_1 = {pp22[59]};
    assign in2090_2 = {pp23[58]};
    Full_Adder FA_2090(s2090, c2090, in2090_1, in2090_2, pp21[60]);
    wire[0:0] s2091, in2091_1, in2091_2;
    wire c2091;
    assign in2091_1 = {pp25[56]};
    assign in2091_2 = {pp26[55]};
    Full_Adder FA_2091(s2091, c2091, in2091_1, in2091_2, pp24[57]);
    wire[0:0] s2092, in2092_1, in2092_2;
    wire c2092;
    assign in2092_1 = {pp28[53]};
    assign in2092_2 = {pp29[52]};
    Full_Adder FA_2092(s2092, c2092, in2092_1, in2092_2, pp27[54]);
    wire[0:0] s2093, in2093_1, in2093_2;
    wire c2093;
    assign in2093_1 = {pp31[50]};
    assign in2093_2 = {pp32[49]};
    Full_Adder FA_2093(s2093, c2093, in2093_1, in2093_2, pp30[51]);
    wire[0:0] s2094, in2094_1, in2094_2;
    wire c2094;
    assign in2094_1 = {pp34[47]};
    assign in2094_2 = {pp35[46]};
    Full_Adder FA_2094(s2094, c2094, in2094_1, in2094_2, pp33[48]);
    wire[0:0] s2095, in2095_1, in2095_2;
    wire c2095;
    assign in2095_1 = {pp37[44]};
    assign in2095_2 = {pp38[43]};
    Full_Adder FA_2095(s2095, c2095, in2095_1, in2095_2, pp36[45]);
    wire[0:0] s2096, in2096_1, in2096_2;
    wire c2096;
    assign in2096_1 = {pp40[41]};
    assign in2096_2 = {pp41[40]};
    Full_Adder FA_2096(s2096, c2096, in2096_1, in2096_2, pp39[42]);
    wire[0:0] s2097, in2097_1, in2097_2;
    wire c2097;
    assign in2097_1 = {pp43[38]};
    assign in2097_2 = {pp44[37]};
    Full_Adder FA_2097(s2097, c2097, in2097_1, in2097_2, pp42[39]);
    wire[0:0] s2098, in2098_1, in2098_2;
    wire c2098;
    assign in2098_1 = {pp46[35]};
    assign in2098_2 = {pp47[34]};
    Full_Adder FA_2098(s2098, c2098, in2098_1, in2098_2, pp45[36]);
    wire[0:0] s2099, in2099_1, in2099_2;
    wire c2099;
    assign in2099_1 = {pp49[32]};
    assign in2099_2 = {pp50[31]};
    Full_Adder FA_2099(s2099, c2099, in2099_1, in2099_2, pp48[33]);
    wire[0:0] s2100, in2100_1, in2100_2;
    wire c2100;
    assign in2100_1 = {pp52[29]};
    assign in2100_2 = {pp53[28]};
    Full_Adder FA_2100(s2100, c2100, in2100_1, in2100_2, pp51[30]);
    wire[0:0] s2101, in2101_1, in2101_2;
    wire c2101;
    assign in2101_1 = {pp55[26]};
    assign in2101_2 = {pp56[25]};
    Full_Adder FA_2101(s2101, c2101, in2101_1, in2101_2, pp54[27]);
    wire[0:0] s2102, in2102_1, in2102_2;
    wire c2102;
    assign in2102_1 = {pp58[23]};
    assign in2102_2 = {pp59[22]};
    Full_Adder FA_2102(s2102, c2102, in2102_1, in2102_2, pp57[24]);
    wire[0:0] s2103, in2103_1, in2103_2;
    wire c2103;
    assign in2103_1 = {pp61[20]};
    assign in2103_2 = {pp62[19]};
    Full_Adder FA_2103(s2103, c2103, in2103_1, in2103_2, pp60[21]);
    wire[0:0] s2104, in2104_1, in2104_2;
    wire c2104;
    assign in2104_1 = {pp64[17]};
    assign in2104_2 = {pp65[16]};
    Full_Adder FA_2104(s2104, c2104, in2104_1, in2104_2, pp63[18]);
    wire[0:0] s2105, in2105_1, in2105_2;
    wire c2105;
    assign in2105_1 = {pp67[14]};
    assign in2105_2 = {pp68[13]};
    Full_Adder FA_2105(s2105, c2105, in2105_1, in2105_2, pp66[15]);
    wire[0:0] s2106, in2106_1, in2106_2;
    wire c2106;
    assign in2106_1 = {pp69[12]};
    assign in2106_2 = {pp70[11]};
    Half_Adder HA_2106(s2106, c2106, in2106_1, in2106_2);
    wire[0:0] s2107, in2107_1, in2107_2;
    wire c2107;
    assign in2107_1 = {pp1[81]};
    assign in2107_2 = {pp2[80]};
    Full_Adder FA_2107(s2107, c2107, in2107_1, in2107_2, pp0[82]);
    wire[0:0] s2108, in2108_1, in2108_2;
    wire c2108;
    assign in2108_1 = {pp4[78]};
    assign in2108_2 = {pp5[77]};
    Full_Adder FA_2108(s2108, c2108, in2108_1, in2108_2, pp3[79]);
    wire[0:0] s2109, in2109_1, in2109_2;
    wire c2109;
    assign in2109_1 = {pp7[75]};
    assign in2109_2 = {pp8[74]};
    Full_Adder FA_2109(s2109, c2109, in2109_1, in2109_2, pp6[76]);
    wire[0:0] s2110, in2110_1, in2110_2;
    wire c2110;
    assign in2110_1 = {pp10[72]};
    assign in2110_2 = {pp11[71]};
    Full_Adder FA_2110(s2110, c2110, in2110_1, in2110_2, pp9[73]);
    wire[0:0] s2111, in2111_1, in2111_2;
    wire c2111;
    assign in2111_1 = {pp13[69]};
    assign in2111_2 = {pp14[68]};
    Full_Adder FA_2111(s2111, c2111, in2111_1, in2111_2, pp12[70]);
    wire[0:0] s2112, in2112_1, in2112_2;
    wire c2112;
    assign in2112_1 = {pp16[66]};
    assign in2112_2 = {pp17[65]};
    Full_Adder FA_2112(s2112, c2112, in2112_1, in2112_2, pp15[67]);
    wire[0:0] s2113, in2113_1, in2113_2;
    wire c2113;
    assign in2113_1 = {pp19[63]};
    assign in2113_2 = {pp20[62]};
    Full_Adder FA_2113(s2113, c2113, in2113_1, in2113_2, pp18[64]);
    wire[0:0] s2114, in2114_1, in2114_2;
    wire c2114;
    assign in2114_1 = {pp22[60]};
    assign in2114_2 = {pp23[59]};
    Full_Adder FA_2114(s2114, c2114, in2114_1, in2114_2, pp21[61]);
    wire[0:0] s2115, in2115_1, in2115_2;
    wire c2115;
    assign in2115_1 = {pp25[57]};
    assign in2115_2 = {pp26[56]};
    Full_Adder FA_2115(s2115, c2115, in2115_1, in2115_2, pp24[58]);
    wire[0:0] s2116, in2116_1, in2116_2;
    wire c2116;
    assign in2116_1 = {pp28[54]};
    assign in2116_2 = {pp29[53]};
    Full_Adder FA_2116(s2116, c2116, in2116_1, in2116_2, pp27[55]);
    wire[0:0] s2117, in2117_1, in2117_2;
    wire c2117;
    assign in2117_1 = {pp31[51]};
    assign in2117_2 = {pp32[50]};
    Full_Adder FA_2117(s2117, c2117, in2117_1, in2117_2, pp30[52]);
    wire[0:0] s2118, in2118_1, in2118_2;
    wire c2118;
    assign in2118_1 = {pp34[48]};
    assign in2118_2 = {pp35[47]};
    Full_Adder FA_2118(s2118, c2118, in2118_1, in2118_2, pp33[49]);
    wire[0:0] s2119, in2119_1, in2119_2;
    wire c2119;
    assign in2119_1 = {pp37[45]};
    assign in2119_2 = {pp38[44]};
    Full_Adder FA_2119(s2119, c2119, in2119_1, in2119_2, pp36[46]);
    wire[0:0] s2120, in2120_1, in2120_2;
    wire c2120;
    assign in2120_1 = {pp40[42]};
    assign in2120_2 = {pp41[41]};
    Full_Adder FA_2120(s2120, c2120, in2120_1, in2120_2, pp39[43]);
    wire[0:0] s2121, in2121_1, in2121_2;
    wire c2121;
    assign in2121_1 = {pp43[39]};
    assign in2121_2 = {pp44[38]};
    Full_Adder FA_2121(s2121, c2121, in2121_1, in2121_2, pp42[40]);
    wire[0:0] s2122, in2122_1, in2122_2;
    wire c2122;
    assign in2122_1 = {pp46[36]};
    assign in2122_2 = {pp47[35]};
    Full_Adder FA_2122(s2122, c2122, in2122_1, in2122_2, pp45[37]);
    wire[0:0] s2123, in2123_1, in2123_2;
    wire c2123;
    assign in2123_1 = {pp49[33]};
    assign in2123_2 = {pp50[32]};
    Full_Adder FA_2123(s2123, c2123, in2123_1, in2123_2, pp48[34]);
    wire[0:0] s2124, in2124_1, in2124_2;
    wire c2124;
    assign in2124_1 = {pp52[30]};
    assign in2124_2 = {pp53[29]};
    Full_Adder FA_2124(s2124, c2124, in2124_1, in2124_2, pp51[31]);
    wire[0:0] s2125, in2125_1, in2125_2;
    wire c2125;
    assign in2125_1 = {pp55[27]};
    assign in2125_2 = {pp56[26]};
    Full_Adder FA_2125(s2125, c2125, in2125_1, in2125_2, pp54[28]);
    wire[0:0] s2126, in2126_1, in2126_2;
    wire c2126;
    assign in2126_1 = {pp58[24]};
    assign in2126_2 = {pp59[23]};
    Full_Adder FA_2126(s2126, c2126, in2126_1, in2126_2, pp57[25]);
    wire[0:0] s2127, in2127_1, in2127_2;
    wire c2127;
    assign in2127_1 = {pp61[21]};
    assign in2127_2 = {pp62[20]};
    Full_Adder FA_2127(s2127, c2127, in2127_1, in2127_2, pp60[22]);
    wire[0:0] s2128, in2128_1, in2128_2;
    wire c2128;
    assign in2128_1 = {pp64[18]};
    assign in2128_2 = {pp65[17]};
    Full_Adder FA_2128(s2128, c2128, in2128_1, in2128_2, pp63[19]);
    wire[0:0] s2129, in2129_1, in2129_2;
    wire c2129;
    assign in2129_1 = {pp67[15]};
    assign in2129_2 = {pp68[14]};
    Full_Adder FA_2129(s2129, c2129, in2129_1, in2129_2, pp66[16]);
    wire[0:0] s2130, in2130_1, in2130_2;
    wire c2130;
    assign in2130_1 = {pp70[12]};
    assign in2130_2 = {pp71[11]};
    Full_Adder FA_2130(s2130, c2130, in2130_1, in2130_2, pp69[13]);
    wire[0:0] s2131, in2131_1, in2131_2;
    wire c2131;
    assign in2131_1 = {pp72[10]};
    assign in2131_2 = {pp73[9]};
    Half_Adder HA_2131(s2131, c2131, in2131_1, in2131_2);
    wire[0:0] s2132, in2132_1, in2132_2;
    wire c2132;
    assign in2132_1 = {pp1[82]};
    assign in2132_2 = {pp2[81]};
    Full_Adder FA_2132(s2132, c2132, in2132_1, in2132_2, pp0[83]);
    wire[0:0] s2133, in2133_1, in2133_2;
    wire c2133;
    assign in2133_1 = {pp4[79]};
    assign in2133_2 = {pp5[78]};
    Full_Adder FA_2133(s2133, c2133, in2133_1, in2133_2, pp3[80]);
    wire[0:0] s2134, in2134_1, in2134_2;
    wire c2134;
    assign in2134_1 = {pp7[76]};
    assign in2134_2 = {pp8[75]};
    Full_Adder FA_2134(s2134, c2134, in2134_1, in2134_2, pp6[77]);
    wire[0:0] s2135, in2135_1, in2135_2;
    wire c2135;
    assign in2135_1 = {pp10[73]};
    assign in2135_2 = {pp11[72]};
    Full_Adder FA_2135(s2135, c2135, in2135_1, in2135_2, pp9[74]);
    wire[0:0] s2136, in2136_1, in2136_2;
    wire c2136;
    assign in2136_1 = {pp13[70]};
    assign in2136_2 = {pp14[69]};
    Full_Adder FA_2136(s2136, c2136, in2136_1, in2136_2, pp12[71]);
    wire[0:0] s2137, in2137_1, in2137_2;
    wire c2137;
    assign in2137_1 = {pp16[67]};
    assign in2137_2 = {pp17[66]};
    Full_Adder FA_2137(s2137, c2137, in2137_1, in2137_2, pp15[68]);
    wire[0:0] s2138, in2138_1, in2138_2;
    wire c2138;
    assign in2138_1 = {pp19[64]};
    assign in2138_2 = {pp20[63]};
    Full_Adder FA_2138(s2138, c2138, in2138_1, in2138_2, pp18[65]);
    wire[0:0] s2139, in2139_1, in2139_2;
    wire c2139;
    assign in2139_1 = {pp22[61]};
    assign in2139_2 = {pp23[60]};
    Full_Adder FA_2139(s2139, c2139, in2139_1, in2139_2, pp21[62]);
    wire[0:0] s2140, in2140_1, in2140_2;
    wire c2140;
    assign in2140_1 = {pp25[58]};
    assign in2140_2 = {pp26[57]};
    Full_Adder FA_2140(s2140, c2140, in2140_1, in2140_2, pp24[59]);
    wire[0:0] s2141, in2141_1, in2141_2;
    wire c2141;
    assign in2141_1 = {pp28[55]};
    assign in2141_2 = {pp29[54]};
    Full_Adder FA_2141(s2141, c2141, in2141_1, in2141_2, pp27[56]);
    wire[0:0] s2142, in2142_1, in2142_2;
    wire c2142;
    assign in2142_1 = {pp31[52]};
    assign in2142_2 = {pp32[51]};
    Full_Adder FA_2142(s2142, c2142, in2142_1, in2142_2, pp30[53]);
    wire[0:0] s2143, in2143_1, in2143_2;
    wire c2143;
    assign in2143_1 = {pp34[49]};
    assign in2143_2 = {pp35[48]};
    Full_Adder FA_2143(s2143, c2143, in2143_1, in2143_2, pp33[50]);
    wire[0:0] s2144, in2144_1, in2144_2;
    wire c2144;
    assign in2144_1 = {pp37[46]};
    assign in2144_2 = {pp38[45]};
    Full_Adder FA_2144(s2144, c2144, in2144_1, in2144_2, pp36[47]);
    wire[0:0] s2145, in2145_1, in2145_2;
    wire c2145;
    assign in2145_1 = {pp40[43]};
    assign in2145_2 = {pp41[42]};
    Full_Adder FA_2145(s2145, c2145, in2145_1, in2145_2, pp39[44]);
    wire[0:0] s2146, in2146_1, in2146_2;
    wire c2146;
    assign in2146_1 = {pp43[40]};
    assign in2146_2 = {pp44[39]};
    Full_Adder FA_2146(s2146, c2146, in2146_1, in2146_2, pp42[41]);
    wire[0:0] s2147, in2147_1, in2147_2;
    wire c2147;
    assign in2147_1 = {pp46[37]};
    assign in2147_2 = {pp47[36]};
    Full_Adder FA_2147(s2147, c2147, in2147_1, in2147_2, pp45[38]);
    wire[0:0] s2148, in2148_1, in2148_2;
    wire c2148;
    assign in2148_1 = {pp49[34]};
    assign in2148_2 = {pp50[33]};
    Full_Adder FA_2148(s2148, c2148, in2148_1, in2148_2, pp48[35]);
    wire[0:0] s2149, in2149_1, in2149_2;
    wire c2149;
    assign in2149_1 = {pp52[31]};
    assign in2149_2 = {pp53[30]};
    Full_Adder FA_2149(s2149, c2149, in2149_1, in2149_2, pp51[32]);
    wire[0:0] s2150, in2150_1, in2150_2;
    wire c2150;
    assign in2150_1 = {pp55[28]};
    assign in2150_2 = {pp56[27]};
    Full_Adder FA_2150(s2150, c2150, in2150_1, in2150_2, pp54[29]);
    wire[0:0] s2151, in2151_1, in2151_2;
    wire c2151;
    assign in2151_1 = {pp58[25]};
    assign in2151_2 = {pp59[24]};
    Full_Adder FA_2151(s2151, c2151, in2151_1, in2151_2, pp57[26]);
    wire[0:0] s2152, in2152_1, in2152_2;
    wire c2152;
    assign in2152_1 = {pp61[22]};
    assign in2152_2 = {pp62[21]};
    Full_Adder FA_2152(s2152, c2152, in2152_1, in2152_2, pp60[23]);
    wire[0:0] s2153, in2153_1, in2153_2;
    wire c2153;
    assign in2153_1 = {pp64[19]};
    assign in2153_2 = {pp65[18]};
    Full_Adder FA_2153(s2153, c2153, in2153_1, in2153_2, pp63[20]);
    wire[0:0] s2154, in2154_1, in2154_2;
    wire c2154;
    assign in2154_1 = {pp67[16]};
    assign in2154_2 = {pp68[15]};
    Full_Adder FA_2154(s2154, c2154, in2154_1, in2154_2, pp66[17]);
    wire[0:0] s2155, in2155_1, in2155_2;
    wire c2155;
    assign in2155_1 = {pp70[13]};
    assign in2155_2 = {pp71[12]};
    Full_Adder FA_2155(s2155, c2155, in2155_1, in2155_2, pp69[14]);
    wire[0:0] s2156, in2156_1, in2156_2;
    wire c2156;
    assign in2156_1 = {pp73[10]};
    assign in2156_2 = {pp74[9]};
    Full_Adder FA_2156(s2156, c2156, in2156_1, in2156_2, pp72[11]);
    wire[0:0] s2157, in2157_1, in2157_2;
    wire c2157;
    assign in2157_1 = {pp75[8]};
    assign in2157_2 = {pp76[7]};
    Half_Adder HA_2157(s2157, c2157, in2157_1, in2157_2);
    wire[0:0] s2158, in2158_1, in2158_2;
    wire c2158;
    assign in2158_1 = {pp1[83]};
    assign in2158_2 = {pp2[82]};
    Full_Adder FA_2158(s2158, c2158, in2158_1, in2158_2, pp0[84]);
    wire[0:0] s2159, in2159_1, in2159_2;
    wire c2159;
    assign in2159_1 = {pp4[80]};
    assign in2159_2 = {pp5[79]};
    Full_Adder FA_2159(s2159, c2159, in2159_1, in2159_2, pp3[81]);
    wire[0:0] s2160, in2160_1, in2160_2;
    wire c2160;
    assign in2160_1 = {pp7[77]};
    assign in2160_2 = {pp8[76]};
    Full_Adder FA_2160(s2160, c2160, in2160_1, in2160_2, pp6[78]);
    wire[0:0] s2161, in2161_1, in2161_2;
    wire c2161;
    assign in2161_1 = {pp10[74]};
    assign in2161_2 = {pp11[73]};
    Full_Adder FA_2161(s2161, c2161, in2161_1, in2161_2, pp9[75]);
    wire[0:0] s2162, in2162_1, in2162_2;
    wire c2162;
    assign in2162_1 = {pp13[71]};
    assign in2162_2 = {pp14[70]};
    Full_Adder FA_2162(s2162, c2162, in2162_1, in2162_2, pp12[72]);
    wire[0:0] s2163, in2163_1, in2163_2;
    wire c2163;
    assign in2163_1 = {pp16[68]};
    assign in2163_2 = {pp17[67]};
    Full_Adder FA_2163(s2163, c2163, in2163_1, in2163_2, pp15[69]);
    wire[0:0] s2164, in2164_1, in2164_2;
    wire c2164;
    assign in2164_1 = {pp19[65]};
    assign in2164_2 = {pp20[64]};
    Full_Adder FA_2164(s2164, c2164, in2164_1, in2164_2, pp18[66]);
    wire[0:0] s2165, in2165_1, in2165_2;
    wire c2165;
    assign in2165_1 = {pp22[62]};
    assign in2165_2 = {pp23[61]};
    Full_Adder FA_2165(s2165, c2165, in2165_1, in2165_2, pp21[63]);
    wire[0:0] s2166, in2166_1, in2166_2;
    wire c2166;
    assign in2166_1 = {pp25[59]};
    assign in2166_2 = {pp26[58]};
    Full_Adder FA_2166(s2166, c2166, in2166_1, in2166_2, pp24[60]);
    wire[0:0] s2167, in2167_1, in2167_2;
    wire c2167;
    assign in2167_1 = {pp28[56]};
    assign in2167_2 = {pp29[55]};
    Full_Adder FA_2167(s2167, c2167, in2167_1, in2167_2, pp27[57]);
    wire[0:0] s2168, in2168_1, in2168_2;
    wire c2168;
    assign in2168_1 = {pp31[53]};
    assign in2168_2 = {pp32[52]};
    Full_Adder FA_2168(s2168, c2168, in2168_1, in2168_2, pp30[54]);
    wire[0:0] s2169, in2169_1, in2169_2;
    wire c2169;
    assign in2169_1 = {pp34[50]};
    assign in2169_2 = {pp35[49]};
    Full_Adder FA_2169(s2169, c2169, in2169_1, in2169_2, pp33[51]);
    wire[0:0] s2170, in2170_1, in2170_2;
    wire c2170;
    assign in2170_1 = {pp37[47]};
    assign in2170_2 = {pp38[46]};
    Full_Adder FA_2170(s2170, c2170, in2170_1, in2170_2, pp36[48]);
    wire[0:0] s2171, in2171_1, in2171_2;
    wire c2171;
    assign in2171_1 = {pp40[44]};
    assign in2171_2 = {pp41[43]};
    Full_Adder FA_2171(s2171, c2171, in2171_1, in2171_2, pp39[45]);
    wire[0:0] s2172, in2172_1, in2172_2;
    wire c2172;
    assign in2172_1 = {pp43[41]};
    assign in2172_2 = {pp44[40]};
    Full_Adder FA_2172(s2172, c2172, in2172_1, in2172_2, pp42[42]);
    wire[0:0] s2173, in2173_1, in2173_2;
    wire c2173;
    assign in2173_1 = {pp46[38]};
    assign in2173_2 = {pp47[37]};
    Full_Adder FA_2173(s2173, c2173, in2173_1, in2173_2, pp45[39]);
    wire[0:0] s2174, in2174_1, in2174_2;
    wire c2174;
    assign in2174_1 = {pp49[35]};
    assign in2174_2 = {pp50[34]};
    Full_Adder FA_2174(s2174, c2174, in2174_1, in2174_2, pp48[36]);
    wire[0:0] s2175, in2175_1, in2175_2;
    wire c2175;
    assign in2175_1 = {pp52[32]};
    assign in2175_2 = {pp53[31]};
    Full_Adder FA_2175(s2175, c2175, in2175_1, in2175_2, pp51[33]);
    wire[0:0] s2176, in2176_1, in2176_2;
    wire c2176;
    assign in2176_1 = {pp55[29]};
    assign in2176_2 = {pp56[28]};
    Full_Adder FA_2176(s2176, c2176, in2176_1, in2176_2, pp54[30]);
    wire[0:0] s2177, in2177_1, in2177_2;
    wire c2177;
    assign in2177_1 = {pp58[26]};
    assign in2177_2 = {pp59[25]};
    Full_Adder FA_2177(s2177, c2177, in2177_1, in2177_2, pp57[27]);
    wire[0:0] s2178, in2178_1, in2178_2;
    wire c2178;
    assign in2178_1 = {pp61[23]};
    assign in2178_2 = {pp62[22]};
    Full_Adder FA_2178(s2178, c2178, in2178_1, in2178_2, pp60[24]);
    wire[0:0] s2179, in2179_1, in2179_2;
    wire c2179;
    assign in2179_1 = {pp64[20]};
    assign in2179_2 = {pp65[19]};
    Full_Adder FA_2179(s2179, c2179, in2179_1, in2179_2, pp63[21]);
    wire[0:0] s2180, in2180_1, in2180_2;
    wire c2180;
    assign in2180_1 = {pp67[17]};
    assign in2180_2 = {pp68[16]};
    Full_Adder FA_2180(s2180, c2180, in2180_1, in2180_2, pp66[18]);
    wire[0:0] s2181, in2181_1, in2181_2;
    wire c2181;
    assign in2181_1 = {pp70[14]};
    assign in2181_2 = {pp71[13]};
    Full_Adder FA_2181(s2181, c2181, in2181_1, in2181_2, pp69[15]);
    wire[0:0] s2182, in2182_1, in2182_2;
    wire c2182;
    assign in2182_1 = {pp73[11]};
    assign in2182_2 = {pp74[10]};
    Full_Adder FA_2182(s2182, c2182, in2182_1, in2182_2, pp72[12]);
    wire[0:0] s2183, in2183_1, in2183_2;
    wire c2183;
    assign in2183_1 = {pp76[8]};
    assign in2183_2 = {pp77[7]};
    Full_Adder FA_2183(s2183, c2183, in2183_1, in2183_2, pp75[9]);
    wire[0:0] s2184, in2184_1, in2184_2;
    wire c2184;
    assign in2184_1 = {pp78[6]};
    assign in2184_2 = {pp79[5]};
    Half_Adder HA_2184(s2184, c2184, in2184_1, in2184_2);
    wire[0:0] s2185, in2185_1, in2185_2;
    wire c2185;
    assign in2185_1 = {pp1[84]};
    assign in2185_2 = {pp2[83]};
    Full_Adder FA_2185(s2185, c2185, in2185_1, in2185_2, pp0[85]);
    wire[0:0] s2186, in2186_1, in2186_2;
    wire c2186;
    assign in2186_1 = {pp4[81]};
    assign in2186_2 = {pp5[80]};
    Full_Adder FA_2186(s2186, c2186, in2186_1, in2186_2, pp3[82]);
    wire[0:0] s2187, in2187_1, in2187_2;
    wire c2187;
    assign in2187_1 = {pp7[78]};
    assign in2187_2 = {pp8[77]};
    Full_Adder FA_2187(s2187, c2187, in2187_1, in2187_2, pp6[79]);
    wire[0:0] s2188, in2188_1, in2188_2;
    wire c2188;
    assign in2188_1 = {pp10[75]};
    assign in2188_2 = {pp11[74]};
    Full_Adder FA_2188(s2188, c2188, in2188_1, in2188_2, pp9[76]);
    wire[0:0] s2189, in2189_1, in2189_2;
    wire c2189;
    assign in2189_1 = {pp13[72]};
    assign in2189_2 = {pp14[71]};
    Full_Adder FA_2189(s2189, c2189, in2189_1, in2189_2, pp12[73]);
    wire[0:0] s2190, in2190_1, in2190_2;
    wire c2190;
    assign in2190_1 = {pp16[69]};
    assign in2190_2 = {pp17[68]};
    Full_Adder FA_2190(s2190, c2190, in2190_1, in2190_2, pp15[70]);
    wire[0:0] s2191, in2191_1, in2191_2;
    wire c2191;
    assign in2191_1 = {pp19[66]};
    assign in2191_2 = {pp20[65]};
    Full_Adder FA_2191(s2191, c2191, in2191_1, in2191_2, pp18[67]);
    wire[0:0] s2192, in2192_1, in2192_2;
    wire c2192;
    assign in2192_1 = {pp22[63]};
    assign in2192_2 = {pp23[62]};
    Full_Adder FA_2192(s2192, c2192, in2192_1, in2192_2, pp21[64]);
    wire[0:0] s2193, in2193_1, in2193_2;
    wire c2193;
    assign in2193_1 = {pp25[60]};
    assign in2193_2 = {pp26[59]};
    Full_Adder FA_2193(s2193, c2193, in2193_1, in2193_2, pp24[61]);
    wire[0:0] s2194, in2194_1, in2194_2;
    wire c2194;
    assign in2194_1 = {pp28[57]};
    assign in2194_2 = {pp29[56]};
    Full_Adder FA_2194(s2194, c2194, in2194_1, in2194_2, pp27[58]);
    wire[0:0] s2195, in2195_1, in2195_2;
    wire c2195;
    assign in2195_1 = {pp31[54]};
    assign in2195_2 = {pp32[53]};
    Full_Adder FA_2195(s2195, c2195, in2195_1, in2195_2, pp30[55]);
    wire[0:0] s2196, in2196_1, in2196_2;
    wire c2196;
    assign in2196_1 = {pp34[51]};
    assign in2196_2 = {pp35[50]};
    Full_Adder FA_2196(s2196, c2196, in2196_1, in2196_2, pp33[52]);
    wire[0:0] s2197, in2197_1, in2197_2;
    wire c2197;
    assign in2197_1 = {pp37[48]};
    assign in2197_2 = {pp38[47]};
    Full_Adder FA_2197(s2197, c2197, in2197_1, in2197_2, pp36[49]);
    wire[0:0] s2198, in2198_1, in2198_2;
    wire c2198;
    assign in2198_1 = {pp40[45]};
    assign in2198_2 = {pp41[44]};
    Full_Adder FA_2198(s2198, c2198, in2198_1, in2198_2, pp39[46]);
    wire[0:0] s2199, in2199_1, in2199_2;
    wire c2199;
    assign in2199_1 = {pp43[42]};
    assign in2199_2 = {pp44[41]};
    Full_Adder FA_2199(s2199, c2199, in2199_1, in2199_2, pp42[43]);
    wire[0:0] s2200, in2200_1, in2200_2;
    wire c2200;
    assign in2200_1 = {pp46[39]};
    assign in2200_2 = {pp47[38]};
    Full_Adder FA_2200(s2200, c2200, in2200_1, in2200_2, pp45[40]);
    wire[0:0] s2201, in2201_1, in2201_2;
    wire c2201;
    assign in2201_1 = {pp49[36]};
    assign in2201_2 = {pp50[35]};
    Full_Adder FA_2201(s2201, c2201, in2201_1, in2201_2, pp48[37]);
    wire[0:0] s2202, in2202_1, in2202_2;
    wire c2202;
    assign in2202_1 = {pp52[33]};
    assign in2202_2 = {pp53[32]};
    Full_Adder FA_2202(s2202, c2202, in2202_1, in2202_2, pp51[34]);
    wire[0:0] s2203, in2203_1, in2203_2;
    wire c2203;
    assign in2203_1 = {pp55[30]};
    assign in2203_2 = {pp56[29]};
    Full_Adder FA_2203(s2203, c2203, in2203_1, in2203_2, pp54[31]);
    wire[0:0] s2204, in2204_1, in2204_2;
    wire c2204;
    assign in2204_1 = {pp58[27]};
    assign in2204_2 = {pp59[26]};
    Full_Adder FA_2204(s2204, c2204, in2204_1, in2204_2, pp57[28]);
    wire[0:0] s2205, in2205_1, in2205_2;
    wire c2205;
    assign in2205_1 = {pp61[24]};
    assign in2205_2 = {pp62[23]};
    Full_Adder FA_2205(s2205, c2205, in2205_1, in2205_2, pp60[25]);
    wire[0:0] s2206, in2206_1, in2206_2;
    wire c2206;
    assign in2206_1 = {pp64[21]};
    assign in2206_2 = {pp65[20]};
    Full_Adder FA_2206(s2206, c2206, in2206_1, in2206_2, pp63[22]);
    wire[0:0] s2207, in2207_1, in2207_2;
    wire c2207;
    assign in2207_1 = {pp67[18]};
    assign in2207_2 = {pp68[17]};
    Full_Adder FA_2207(s2207, c2207, in2207_1, in2207_2, pp66[19]);
    wire[0:0] s2208, in2208_1, in2208_2;
    wire c2208;
    assign in2208_1 = {pp70[15]};
    assign in2208_2 = {pp71[14]};
    Full_Adder FA_2208(s2208, c2208, in2208_1, in2208_2, pp69[16]);
    wire[0:0] s2209, in2209_1, in2209_2;
    wire c2209;
    assign in2209_1 = {pp73[12]};
    assign in2209_2 = {pp74[11]};
    Full_Adder FA_2209(s2209, c2209, in2209_1, in2209_2, pp72[13]);
    wire[0:0] s2210, in2210_1, in2210_2;
    wire c2210;
    assign in2210_1 = {pp76[9]};
    assign in2210_2 = {pp77[8]};
    Full_Adder FA_2210(s2210, c2210, in2210_1, in2210_2, pp75[10]);
    wire[0:0] s2211, in2211_1, in2211_2;
    wire c2211;
    assign in2211_1 = {pp79[6]};
    assign in2211_2 = {pp80[5]};
    Full_Adder FA_2211(s2211, c2211, in2211_1, in2211_2, pp78[7]);
    wire[0:0] s2212, in2212_1, in2212_2;
    wire c2212;
    assign in2212_1 = {pp81[4]};
    assign in2212_2 = {pp82[3]};
    Half_Adder HA_2212(s2212, c2212, in2212_1, in2212_2);
    wire[0:0] s2213, in2213_1, in2213_2;
    wire c2213;
    assign in2213_1 = {pp3[83]};
    assign in2213_2 = {pp4[82]};
    Full_Adder FA_2213(s2213, c2213, in2213_1, in2213_2, pp2[84]);
    wire[0:0] s2214, in2214_1, in2214_2;
    wire c2214;
    assign in2214_1 = {pp6[80]};
    assign in2214_2 = {pp7[79]};
    Full_Adder FA_2214(s2214, c2214, in2214_1, in2214_2, pp5[81]);
    wire[0:0] s2215, in2215_1, in2215_2;
    wire c2215;
    assign in2215_1 = {pp9[77]};
    assign in2215_2 = {pp10[76]};
    Full_Adder FA_2215(s2215, c2215, in2215_1, in2215_2, pp8[78]);
    wire[0:0] s2216, in2216_1, in2216_2;
    wire c2216;
    assign in2216_1 = {pp12[74]};
    assign in2216_2 = {pp13[73]};
    Full_Adder FA_2216(s2216, c2216, in2216_1, in2216_2, pp11[75]);
    wire[0:0] s2217, in2217_1, in2217_2;
    wire c2217;
    assign in2217_1 = {pp15[71]};
    assign in2217_2 = {pp16[70]};
    Full_Adder FA_2217(s2217, c2217, in2217_1, in2217_2, pp14[72]);
    wire[0:0] s2218, in2218_1, in2218_2;
    wire c2218;
    assign in2218_1 = {pp18[68]};
    assign in2218_2 = {pp19[67]};
    Full_Adder FA_2218(s2218, c2218, in2218_1, in2218_2, pp17[69]);
    wire[0:0] s2219, in2219_1, in2219_2;
    wire c2219;
    assign in2219_1 = {pp21[65]};
    assign in2219_2 = {pp22[64]};
    Full_Adder FA_2219(s2219, c2219, in2219_1, in2219_2, pp20[66]);
    wire[0:0] s2220, in2220_1, in2220_2;
    wire c2220;
    assign in2220_1 = {pp24[62]};
    assign in2220_2 = {pp25[61]};
    Full_Adder FA_2220(s2220, c2220, in2220_1, in2220_2, pp23[63]);
    wire[0:0] s2221, in2221_1, in2221_2;
    wire c2221;
    assign in2221_1 = {pp27[59]};
    assign in2221_2 = {pp28[58]};
    Full_Adder FA_2221(s2221, c2221, in2221_1, in2221_2, pp26[60]);
    wire[0:0] s2222, in2222_1, in2222_2;
    wire c2222;
    assign in2222_1 = {pp30[56]};
    assign in2222_2 = {pp31[55]};
    Full_Adder FA_2222(s2222, c2222, in2222_1, in2222_2, pp29[57]);
    wire[0:0] s2223, in2223_1, in2223_2;
    wire c2223;
    assign in2223_1 = {pp33[53]};
    assign in2223_2 = {pp34[52]};
    Full_Adder FA_2223(s2223, c2223, in2223_1, in2223_2, pp32[54]);
    wire[0:0] s2224, in2224_1, in2224_2;
    wire c2224;
    assign in2224_1 = {pp36[50]};
    assign in2224_2 = {pp37[49]};
    Full_Adder FA_2224(s2224, c2224, in2224_1, in2224_2, pp35[51]);
    wire[0:0] s2225, in2225_1, in2225_2;
    wire c2225;
    assign in2225_1 = {pp39[47]};
    assign in2225_2 = {pp40[46]};
    Full_Adder FA_2225(s2225, c2225, in2225_1, in2225_2, pp38[48]);
    wire[0:0] s2226, in2226_1, in2226_2;
    wire c2226;
    assign in2226_1 = {pp42[44]};
    assign in2226_2 = {pp43[43]};
    Full_Adder FA_2226(s2226, c2226, in2226_1, in2226_2, pp41[45]);
    wire[0:0] s2227, in2227_1, in2227_2;
    wire c2227;
    assign in2227_1 = {pp45[41]};
    assign in2227_2 = {pp46[40]};
    Full_Adder FA_2227(s2227, c2227, in2227_1, in2227_2, pp44[42]);
    wire[0:0] s2228, in2228_1, in2228_2;
    wire c2228;
    assign in2228_1 = {pp48[38]};
    assign in2228_2 = {pp49[37]};
    Full_Adder FA_2228(s2228, c2228, in2228_1, in2228_2, pp47[39]);
    wire[0:0] s2229, in2229_1, in2229_2;
    wire c2229;
    assign in2229_1 = {pp51[35]};
    assign in2229_2 = {pp52[34]};
    Full_Adder FA_2229(s2229, c2229, in2229_1, in2229_2, pp50[36]);
    wire[0:0] s2230, in2230_1, in2230_2;
    wire c2230;
    assign in2230_1 = {pp54[32]};
    assign in2230_2 = {pp55[31]};
    Full_Adder FA_2230(s2230, c2230, in2230_1, in2230_2, pp53[33]);
    wire[0:0] s2231, in2231_1, in2231_2;
    wire c2231;
    assign in2231_1 = {pp57[29]};
    assign in2231_2 = {pp58[28]};
    Full_Adder FA_2231(s2231, c2231, in2231_1, in2231_2, pp56[30]);
    wire[0:0] s2232, in2232_1, in2232_2;
    wire c2232;
    assign in2232_1 = {pp60[26]};
    assign in2232_2 = {pp61[25]};
    Full_Adder FA_2232(s2232, c2232, in2232_1, in2232_2, pp59[27]);
    wire[0:0] s2233, in2233_1, in2233_2;
    wire c2233;
    assign in2233_1 = {pp63[23]};
    assign in2233_2 = {pp64[22]};
    Full_Adder FA_2233(s2233, c2233, in2233_1, in2233_2, pp62[24]);
    wire[0:0] s2234, in2234_1, in2234_2;
    wire c2234;
    assign in2234_1 = {pp66[20]};
    assign in2234_2 = {pp67[19]};
    Full_Adder FA_2234(s2234, c2234, in2234_1, in2234_2, pp65[21]);
    wire[0:0] s2235, in2235_1, in2235_2;
    wire c2235;
    assign in2235_1 = {pp69[17]};
    assign in2235_2 = {pp70[16]};
    Full_Adder FA_2235(s2235, c2235, in2235_1, in2235_2, pp68[18]);
    wire[0:0] s2236, in2236_1, in2236_2;
    wire c2236;
    assign in2236_1 = {pp72[14]};
    assign in2236_2 = {pp73[13]};
    Full_Adder FA_2236(s2236, c2236, in2236_1, in2236_2, pp71[15]);
    wire[0:0] s2237, in2237_1, in2237_2;
    wire c2237;
    assign in2237_1 = {pp75[11]};
    assign in2237_2 = {pp76[10]};
    Full_Adder FA_2237(s2237, c2237, in2237_1, in2237_2, pp74[12]);
    wire[0:0] s2238, in2238_1, in2238_2;
    wire c2238;
    assign in2238_1 = {pp78[8]};
    assign in2238_2 = {pp79[7]};
    Full_Adder FA_2238(s2238, c2238, in2238_1, in2238_2, pp77[9]);
    wire[0:0] s2239, in2239_1, in2239_2;
    wire c2239;
    assign in2239_1 = {pp81[5]};
    assign in2239_2 = {pp82[4]};
    Full_Adder FA_2239(s2239, c2239, in2239_1, in2239_2, pp80[6]);
    wire[0:0] s2240, in2240_1, in2240_2;
    wire c2240;
    assign in2240_1 = {pp84[2]};
    assign in2240_2 = {pp85[1]};
    Full_Adder FA_2240(s2240, c2240, in2240_1, in2240_2, pp83[3]);
    wire[0:0] s2241, in2241_1, in2241_2;
    wire c2241;
    assign in2241_1 = {pp6[81]};
    assign in2241_2 = {pp7[80]};
    Full_Adder FA_2241(s2241, c2241, in2241_1, in2241_2, pp5[82]);
    wire[0:0] s2242, in2242_1, in2242_2;
    wire c2242;
    assign in2242_1 = {pp9[78]};
    assign in2242_2 = {pp10[77]};
    Full_Adder FA_2242(s2242, c2242, in2242_1, in2242_2, pp8[79]);
    wire[0:0] s2243, in2243_1, in2243_2;
    wire c2243;
    assign in2243_1 = {pp12[75]};
    assign in2243_2 = {pp13[74]};
    Full_Adder FA_2243(s2243, c2243, in2243_1, in2243_2, pp11[76]);
    wire[0:0] s2244, in2244_1, in2244_2;
    wire c2244;
    assign in2244_1 = {pp15[72]};
    assign in2244_2 = {pp16[71]};
    Full_Adder FA_2244(s2244, c2244, in2244_1, in2244_2, pp14[73]);
    wire[0:0] s2245, in2245_1, in2245_2;
    wire c2245;
    assign in2245_1 = {pp18[69]};
    assign in2245_2 = {pp19[68]};
    Full_Adder FA_2245(s2245, c2245, in2245_1, in2245_2, pp17[70]);
    wire[0:0] s2246, in2246_1, in2246_2;
    wire c2246;
    assign in2246_1 = {pp21[66]};
    assign in2246_2 = {pp22[65]};
    Full_Adder FA_2246(s2246, c2246, in2246_1, in2246_2, pp20[67]);
    wire[0:0] s2247, in2247_1, in2247_2;
    wire c2247;
    assign in2247_1 = {pp24[63]};
    assign in2247_2 = {pp25[62]};
    Full_Adder FA_2247(s2247, c2247, in2247_1, in2247_2, pp23[64]);
    wire[0:0] s2248, in2248_1, in2248_2;
    wire c2248;
    assign in2248_1 = {pp27[60]};
    assign in2248_2 = {pp28[59]};
    Full_Adder FA_2248(s2248, c2248, in2248_1, in2248_2, pp26[61]);
    wire[0:0] s2249, in2249_1, in2249_2;
    wire c2249;
    assign in2249_1 = {pp30[57]};
    assign in2249_2 = {pp31[56]};
    Full_Adder FA_2249(s2249, c2249, in2249_1, in2249_2, pp29[58]);
    wire[0:0] s2250, in2250_1, in2250_2;
    wire c2250;
    assign in2250_1 = {pp33[54]};
    assign in2250_2 = {pp34[53]};
    Full_Adder FA_2250(s2250, c2250, in2250_1, in2250_2, pp32[55]);
    wire[0:0] s2251, in2251_1, in2251_2;
    wire c2251;
    assign in2251_1 = {pp36[51]};
    assign in2251_2 = {pp37[50]};
    Full_Adder FA_2251(s2251, c2251, in2251_1, in2251_2, pp35[52]);
    wire[0:0] s2252, in2252_1, in2252_2;
    wire c2252;
    assign in2252_1 = {pp39[48]};
    assign in2252_2 = {pp40[47]};
    Full_Adder FA_2252(s2252, c2252, in2252_1, in2252_2, pp38[49]);
    wire[0:0] s2253, in2253_1, in2253_2;
    wire c2253;
    assign in2253_1 = {pp42[45]};
    assign in2253_2 = {pp43[44]};
    Full_Adder FA_2253(s2253, c2253, in2253_1, in2253_2, pp41[46]);
    wire[0:0] s2254, in2254_1, in2254_2;
    wire c2254;
    assign in2254_1 = {pp45[42]};
    assign in2254_2 = {pp46[41]};
    Full_Adder FA_2254(s2254, c2254, in2254_1, in2254_2, pp44[43]);
    wire[0:0] s2255, in2255_1, in2255_2;
    wire c2255;
    assign in2255_1 = {pp48[39]};
    assign in2255_2 = {pp49[38]};
    Full_Adder FA_2255(s2255, c2255, in2255_1, in2255_2, pp47[40]);
    wire[0:0] s2256, in2256_1, in2256_2;
    wire c2256;
    assign in2256_1 = {pp51[36]};
    assign in2256_2 = {pp52[35]};
    Full_Adder FA_2256(s2256, c2256, in2256_1, in2256_2, pp50[37]);
    wire[0:0] s2257, in2257_1, in2257_2;
    wire c2257;
    assign in2257_1 = {pp54[33]};
    assign in2257_2 = {pp55[32]};
    Full_Adder FA_2257(s2257, c2257, in2257_1, in2257_2, pp53[34]);
    wire[0:0] s2258, in2258_1, in2258_2;
    wire c2258;
    assign in2258_1 = {pp57[30]};
    assign in2258_2 = {pp58[29]};
    Full_Adder FA_2258(s2258, c2258, in2258_1, in2258_2, pp56[31]);
    wire[0:0] s2259, in2259_1, in2259_2;
    wire c2259;
    assign in2259_1 = {pp60[27]};
    assign in2259_2 = {pp61[26]};
    Full_Adder FA_2259(s2259, c2259, in2259_1, in2259_2, pp59[28]);
    wire[0:0] s2260, in2260_1, in2260_2;
    wire c2260;
    assign in2260_1 = {pp63[24]};
    assign in2260_2 = {pp64[23]};
    Full_Adder FA_2260(s2260, c2260, in2260_1, in2260_2, pp62[25]);
    wire[0:0] s2261, in2261_1, in2261_2;
    wire c2261;
    assign in2261_1 = {pp66[21]};
    assign in2261_2 = {pp67[20]};
    Full_Adder FA_2261(s2261, c2261, in2261_1, in2261_2, pp65[22]);
    wire[0:0] s2262, in2262_1, in2262_2;
    wire c2262;
    assign in2262_1 = {pp69[18]};
    assign in2262_2 = {pp70[17]};
    Full_Adder FA_2262(s2262, c2262, in2262_1, in2262_2, pp68[19]);
    wire[0:0] s2263, in2263_1, in2263_2;
    wire c2263;
    assign in2263_1 = {pp72[15]};
    assign in2263_2 = {pp73[14]};
    Full_Adder FA_2263(s2263, c2263, in2263_1, in2263_2, pp71[16]);
    wire[0:0] s2264, in2264_1, in2264_2;
    wire c2264;
    assign in2264_1 = {pp75[12]};
    assign in2264_2 = {pp76[11]};
    Full_Adder FA_2264(s2264, c2264, in2264_1, in2264_2, pp74[13]);
    wire[0:0] s2265, in2265_1, in2265_2;
    wire c2265;
    assign in2265_1 = {pp78[9]};
    assign in2265_2 = {pp79[8]};
    Full_Adder FA_2265(s2265, c2265, in2265_1, in2265_2, pp77[10]);
    wire[0:0] s2266, in2266_1, in2266_2;
    wire c2266;
    assign in2266_1 = {pp81[6]};
    assign in2266_2 = {pp82[5]};
    Full_Adder FA_2266(s2266, c2266, in2266_1, in2266_2, pp80[7]);
    wire[0:0] s2267, in2267_1, in2267_2;
    wire c2267;
    assign in2267_1 = {pp84[3]};
    assign in2267_2 = {pp85[2]};
    Full_Adder FA_2267(s2267, c2267, in2267_1, in2267_2, pp83[4]);
    wire[0:0] s2268, in2268_1, in2268_2;
    wire c2268;
    assign in2268_1 = {pp87[0]};
    assign in2268_2 = {c1};
    Full_Adder FA_2268(s2268, c2268, in2268_1, in2268_2, pp86[1]);
    wire[0:0] s2269, in2269_1, in2269_2;
    wire c2269;
    assign in2269_1 = {pp9[79]};
    assign in2269_2 = {pp10[78]};
    Full_Adder FA_2269(s2269, c2269, in2269_1, in2269_2, pp8[80]);
    wire[0:0] s2270, in2270_1, in2270_2;
    wire c2270;
    assign in2270_1 = {pp12[76]};
    assign in2270_2 = {pp13[75]};
    Full_Adder FA_2270(s2270, c2270, in2270_1, in2270_2, pp11[77]);
    wire[0:0] s2271, in2271_1, in2271_2;
    wire c2271;
    assign in2271_1 = {pp15[73]};
    assign in2271_2 = {pp16[72]};
    Full_Adder FA_2271(s2271, c2271, in2271_1, in2271_2, pp14[74]);
    wire[0:0] s2272, in2272_1, in2272_2;
    wire c2272;
    assign in2272_1 = {pp18[70]};
    assign in2272_2 = {pp19[69]};
    Full_Adder FA_2272(s2272, c2272, in2272_1, in2272_2, pp17[71]);
    wire[0:0] s2273, in2273_1, in2273_2;
    wire c2273;
    assign in2273_1 = {pp21[67]};
    assign in2273_2 = {pp22[66]};
    Full_Adder FA_2273(s2273, c2273, in2273_1, in2273_2, pp20[68]);
    wire[0:0] s2274, in2274_1, in2274_2;
    wire c2274;
    assign in2274_1 = {pp24[64]};
    assign in2274_2 = {pp25[63]};
    Full_Adder FA_2274(s2274, c2274, in2274_1, in2274_2, pp23[65]);
    wire[0:0] s2275, in2275_1, in2275_2;
    wire c2275;
    assign in2275_1 = {pp27[61]};
    assign in2275_2 = {pp28[60]};
    Full_Adder FA_2275(s2275, c2275, in2275_1, in2275_2, pp26[62]);
    wire[0:0] s2276, in2276_1, in2276_2;
    wire c2276;
    assign in2276_1 = {pp30[58]};
    assign in2276_2 = {pp31[57]};
    Full_Adder FA_2276(s2276, c2276, in2276_1, in2276_2, pp29[59]);
    wire[0:0] s2277, in2277_1, in2277_2;
    wire c2277;
    assign in2277_1 = {pp33[55]};
    assign in2277_2 = {pp34[54]};
    Full_Adder FA_2277(s2277, c2277, in2277_1, in2277_2, pp32[56]);
    wire[0:0] s2278, in2278_1, in2278_2;
    wire c2278;
    assign in2278_1 = {pp36[52]};
    assign in2278_2 = {pp37[51]};
    Full_Adder FA_2278(s2278, c2278, in2278_1, in2278_2, pp35[53]);
    wire[0:0] s2279, in2279_1, in2279_2;
    wire c2279;
    assign in2279_1 = {pp39[49]};
    assign in2279_2 = {pp40[48]};
    Full_Adder FA_2279(s2279, c2279, in2279_1, in2279_2, pp38[50]);
    wire[0:0] s2280, in2280_1, in2280_2;
    wire c2280;
    assign in2280_1 = {pp42[46]};
    assign in2280_2 = {pp43[45]};
    Full_Adder FA_2280(s2280, c2280, in2280_1, in2280_2, pp41[47]);
    wire[0:0] s2281, in2281_1, in2281_2;
    wire c2281;
    assign in2281_1 = {pp45[43]};
    assign in2281_2 = {pp46[42]};
    Full_Adder FA_2281(s2281, c2281, in2281_1, in2281_2, pp44[44]);
    wire[0:0] s2282, in2282_1, in2282_2;
    wire c2282;
    assign in2282_1 = {pp48[40]};
    assign in2282_2 = {pp49[39]};
    Full_Adder FA_2282(s2282, c2282, in2282_1, in2282_2, pp47[41]);
    wire[0:0] s2283, in2283_1, in2283_2;
    wire c2283;
    assign in2283_1 = {pp51[37]};
    assign in2283_2 = {pp52[36]};
    Full_Adder FA_2283(s2283, c2283, in2283_1, in2283_2, pp50[38]);
    wire[0:0] s2284, in2284_1, in2284_2;
    wire c2284;
    assign in2284_1 = {pp54[34]};
    assign in2284_2 = {pp55[33]};
    Full_Adder FA_2284(s2284, c2284, in2284_1, in2284_2, pp53[35]);
    wire[0:0] s2285, in2285_1, in2285_2;
    wire c2285;
    assign in2285_1 = {pp57[31]};
    assign in2285_2 = {pp58[30]};
    Full_Adder FA_2285(s2285, c2285, in2285_1, in2285_2, pp56[32]);
    wire[0:0] s2286, in2286_1, in2286_2;
    wire c2286;
    assign in2286_1 = {pp60[28]};
    assign in2286_2 = {pp61[27]};
    Full_Adder FA_2286(s2286, c2286, in2286_1, in2286_2, pp59[29]);
    wire[0:0] s2287, in2287_1, in2287_2;
    wire c2287;
    assign in2287_1 = {pp63[25]};
    assign in2287_2 = {pp64[24]};
    Full_Adder FA_2287(s2287, c2287, in2287_1, in2287_2, pp62[26]);
    wire[0:0] s2288, in2288_1, in2288_2;
    wire c2288;
    assign in2288_1 = {pp66[22]};
    assign in2288_2 = {pp67[21]};
    Full_Adder FA_2288(s2288, c2288, in2288_1, in2288_2, pp65[23]);
    wire[0:0] s2289, in2289_1, in2289_2;
    wire c2289;
    assign in2289_1 = {pp69[19]};
    assign in2289_2 = {pp70[18]};
    Full_Adder FA_2289(s2289, c2289, in2289_1, in2289_2, pp68[20]);
    wire[0:0] s2290, in2290_1, in2290_2;
    wire c2290;
    assign in2290_1 = {pp72[16]};
    assign in2290_2 = {pp73[15]};
    Full_Adder FA_2290(s2290, c2290, in2290_1, in2290_2, pp71[17]);
    wire[0:0] s2291, in2291_1, in2291_2;
    wire c2291;
    assign in2291_1 = {pp75[13]};
    assign in2291_2 = {pp76[12]};
    Full_Adder FA_2291(s2291, c2291, in2291_1, in2291_2, pp74[14]);
    wire[0:0] s2292, in2292_1, in2292_2;
    wire c2292;
    assign in2292_1 = {pp78[10]};
    assign in2292_2 = {pp79[9]};
    Full_Adder FA_2292(s2292, c2292, in2292_1, in2292_2, pp77[11]);
    wire[0:0] s2293, in2293_1, in2293_2;
    wire c2293;
    assign in2293_1 = {pp81[7]};
    assign in2293_2 = {pp82[6]};
    Full_Adder FA_2293(s2293, c2293, in2293_1, in2293_2, pp80[8]);
    wire[0:0] s2294, in2294_1, in2294_2;
    wire c2294;
    assign in2294_1 = {pp84[4]};
    assign in2294_2 = {pp85[3]};
    Full_Adder FA_2294(s2294, c2294, in2294_1, in2294_2, pp83[5]);
    wire[0:0] s2295, in2295_1, in2295_2;
    wire c2295;
    assign in2295_1 = {pp87[1]};
    assign in2295_2 = {pp88[0]};
    Full_Adder FA_2295(s2295, c2295, in2295_1, in2295_2, pp86[2]);
    wire[0:0] s2296, in2296_1, in2296_2;
    wire c2296;
    assign in2296_1 = {c3};
    assign in2296_2 = {s4[0]};
    Full_Adder FA_2296(s2296, c2296, in2296_1, in2296_2, c2);
    wire[0:0] s2297, in2297_1, in2297_2;
    wire c2297;
    assign in2297_1 = {pp12[77]};
    assign in2297_2 = {pp13[76]};
    Full_Adder FA_2297(s2297, c2297, in2297_1, in2297_2, pp11[78]);
    wire[0:0] s2298, in2298_1, in2298_2;
    wire c2298;
    assign in2298_1 = {pp15[74]};
    assign in2298_2 = {pp16[73]};
    Full_Adder FA_2298(s2298, c2298, in2298_1, in2298_2, pp14[75]);
    wire[0:0] s2299, in2299_1, in2299_2;
    wire c2299;
    assign in2299_1 = {pp18[71]};
    assign in2299_2 = {pp19[70]};
    Full_Adder FA_2299(s2299, c2299, in2299_1, in2299_2, pp17[72]);
    wire[0:0] s2300, in2300_1, in2300_2;
    wire c2300;
    assign in2300_1 = {pp21[68]};
    assign in2300_2 = {pp22[67]};
    Full_Adder FA_2300(s2300, c2300, in2300_1, in2300_2, pp20[69]);
    wire[0:0] s2301, in2301_1, in2301_2;
    wire c2301;
    assign in2301_1 = {pp24[65]};
    assign in2301_2 = {pp25[64]};
    Full_Adder FA_2301(s2301, c2301, in2301_1, in2301_2, pp23[66]);
    wire[0:0] s2302, in2302_1, in2302_2;
    wire c2302;
    assign in2302_1 = {pp27[62]};
    assign in2302_2 = {pp28[61]};
    Full_Adder FA_2302(s2302, c2302, in2302_1, in2302_2, pp26[63]);
    wire[0:0] s2303, in2303_1, in2303_2;
    wire c2303;
    assign in2303_1 = {pp30[59]};
    assign in2303_2 = {pp31[58]};
    Full_Adder FA_2303(s2303, c2303, in2303_1, in2303_2, pp29[60]);
    wire[0:0] s2304, in2304_1, in2304_2;
    wire c2304;
    assign in2304_1 = {pp33[56]};
    assign in2304_2 = {pp34[55]};
    Full_Adder FA_2304(s2304, c2304, in2304_1, in2304_2, pp32[57]);
    wire[0:0] s2305, in2305_1, in2305_2;
    wire c2305;
    assign in2305_1 = {pp36[53]};
    assign in2305_2 = {pp37[52]};
    Full_Adder FA_2305(s2305, c2305, in2305_1, in2305_2, pp35[54]);
    wire[0:0] s2306, in2306_1, in2306_2;
    wire c2306;
    assign in2306_1 = {pp39[50]};
    assign in2306_2 = {pp40[49]};
    Full_Adder FA_2306(s2306, c2306, in2306_1, in2306_2, pp38[51]);
    wire[0:0] s2307, in2307_1, in2307_2;
    wire c2307;
    assign in2307_1 = {pp42[47]};
    assign in2307_2 = {pp43[46]};
    Full_Adder FA_2307(s2307, c2307, in2307_1, in2307_2, pp41[48]);
    wire[0:0] s2308, in2308_1, in2308_2;
    wire c2308;
    assign in2308_1 = {pp45[44]};
    assign in2308_2 = {pp46[43]};
    Full_Adder FA_2308(s2308, c2308, in2308_1, in2308_2, pp44[45]);
    wire[0:0] s2309, in2309_1, in2309_2;
    wire c2309;
    assign in2309_1 = {pp48[41]};
    assign in2309_2 = {pp49[40]};
    Full_Adder FA_2309(s2309, c2309, in2309_1, in2309_2, pp47[42]);
    wire[0:0] s2310, in2310_1, in2310_2;
    wire c2310;
    assign in2310_1 = {pp51[38]};
    assign in2310_2 = {pp52[37]};
    Full_Adder FA_2310(s2310, c2310, in2310_1, in2310_2, pp50[39]);
    wire[0:0] s2311, in2311_1, in2311_2;
    wire c2311;
    assign in2311_1 = {pp54[35]};
    assign in2311_2 = {pp55[34]};
    Full_Adder FA_2311(s2311, c2311, in2311_1, in2311_2, pp53[36]);
    wire[0:0] s2312, in2312_1, in2312_2;
    wire c2312;
    assign in2312_1 = {pp57[32]};
    assign in2312_2 = {pp58[31]};
    Full_Adder FA_2312(s2312, c2312, in2312_1, in2312_2, pp56[33]);
    wire[0:0] s2313, in2313_1, in2313_2;
    wire c2313;
    assign in2313_1 = {pp60[29]};
    assign in2313_2 = {pp61[28]};
    Full_Adder FA_2313(s2313, c2313, in2313_1, in2313_2, pp59[30]);
    wire[0:0] s2314, in2314_1, in2314_2;
    wire c2314;
    assign in2314_1 = {pp63[26]};
    assign in2314_2 = {pp64[25]};
    Full_Adder FA_2314(s2314, c2314, in2314_1, in2314_2, pp62[27]);
    wire[0:0] s2315, in2315_1, in2315_2;
    wire c2315;
    assign in2315_1 = {pp66[23]};
    assign in2315_2 = {pp67[22]};
    Full_Adder FA_2315(s2315, c2315, in2315_1, in2315_2, pp65[24]);
    wire[0:0] s2316, in2316_1, in2316_2;
    wire c2316;
    assign in2316_1 = {pp69[20]};
    assign in2316_2 = {pp70[19]};
    Full_Adder FA_2316(s2316, c2316, in2316_1, in2316_2, pp68[21]);
    wire[0:0] s2317, in2317_1, in2317_2;
    wire c2317;
    assign in2317_1 = {pp72[17]};
    assign in2317_2 = {pp73[16]};
    Full_Adder FA_2317(s2317, c2317, in2317_1, in2317_2, pp71[18]);
    wire[0:0] s2318, in2318_1, in2318_2;
    wire c2318;
    assign in2318_1 = {pp75[14]};
    assign in2318_2 = {pp76[13]};
    Full_Adder FA_2318(s2318, c2318, in2318_1, in2318_2, pp74[15]);
    wire[0:0] s2319, in2319_1, in2319_2;
    wire c2319;
    assign in2319_1 = {pp78[11]};
    assign in2319_2 = {pp79[10]};
    Full_Adder FA_2319(s2319, c2319, in2319_1, in2319_2, pp77[12]);
    wire[0:0] s2320, in2320_1, in2320_2;
    wire c2320;
    assign in2320_1 = {pp81[8]};
    assign in2320_2 = {pp82[7]};
    Full_Adder FA_2320(s2320, c2320, in2320_1, in2320_2, pp80[9]);
    wire[0:0] s2321, in2321_1, in2321_2;
    wire c2321;
    assign in2321_1 = {pp84[5]};
    assign in2321_2 = {pp85[4]};
    Full_Adder FA_2321(s2321, c2321, in2321_1, in2321_2, pp83[6]);
    wire[0:0] s2322, in2322_1, in2322_2;
    wire c2322;
    assign in2322_1 = {pp87[2]};
    assign in2322_2 = {pp88[1]};
    Full_Adder FA_2322(s2322, c2322, in2322_1, in2322_2, pp86[3]);
    wire[0:0] s2323, in2323_1, in2323_2;
    wire c2323;
    assign in2323_1 = {c4};
    assign in2323_2 = {c5};
    Full_Adder FA_2323(s2323, c2323, in2323_1, in2323_2, pp89[0]);
    wire[0:0] s2324, in2324_1, in2324_2;
    wire c2324;
    assign in2324_1 = {s7[0]};
    assign in2324_2 = {s8[0]};
    Full_Adder FA_2324(s2324, c2324, in2324_1, in2324_2, c6);
    wire[0:0] s2325, in2325_1, in2325_2;
    wire c2325;
    assign in2325_1 = {pp15[75]};
    assign in2325_2 = {pp16[74]};
    Full_Adder FA_2325(s2325, c2325, in2325_1, in2325_2, pp14[76]);
    wire[0:0] s2326, in2326_1, in2326_2;
    wire c2326;
    assign in2326_1 = {pp18[72]};
    assign in2326_2 = {pp19[71]};
    Full_Adder FA_2326(s2326, c2326, in2326_1, in2326_2, pp17[73]);
    wire[0:0] s2327, in2327_1, in2327_2;
    wire c2327;
    assign in2327_1 = {pp21[69]};
    assign in2327_2 = {pp22[68]};
    Full_Adder FA_2327(s2327, c2327, in2327_1, in2327_2, pp20[70]);
    wire[0:0] s2328, in2328_1, in2328_2;
    wire c2328;
    assign in2328_1 = {pp24[66]};
    assign in2328_2 = {pp25[65]};
    Full_Adder FA_2328(s2328, c2328, in2328_1, in2328_2, pp23[67]);
    wire[0:0] s2329, in2329_1, in2329_2;
    wire c2329;
    assign in2329_1 = {pp27[63]};
    assign in2329_2 = {pp28[62]};
    Full_Adder FA_2329(s2329, c2329, in2329_1, in2329_2, pp26[64]);
    wire[0:0] s2330, in2330_1, in2330_2;
    wire c2330;
    assign in2330_1 = {pp30[60]};
    assign in2330_2 = {pp31[59]};
    Full_Adder FA_2330(s2330, c2330, in2330_1, in2330_2, pp29[61]);
    wire[0:0] s2331, in2331_1, in2331_2;
    wire c2331;
    assign in2331_1 = {pp33[57]};
    assign in2331_2 = {pp34[56]};
    Full_Adder FA_2331(s2331, c2331, in2331_1, in2331_2, pp32[58]);
    wire[0:0] s2332, in2332_1, in2332_2;
    wire c2332;
    assign in2332_1 = {pp36[54]};
    assign in2332_2 = {pp37[53]};
    Full_Adder FA_2332(s2332, c2332, in2332_1, in2332_2, pp35[55]);
    wire[0:0] s2333, in2333_1, in2333_2;
    wire c2333;
    assign in2333_1 = {pp39[51]};
    assign in2333_2 = {pp40[50]};
    Full_Adder FA_2333(s2333, c2333, in2333_1, in2333_2, pp38[52]);
    wire[0:0] s2334, in2334_1, in2334_2;
    wire c2334;
    assign in2334_1 = {pp42[48]};
    assign in2334_2 = {pp43[47]};
    Full_Adder FA_2334(s2334, c2334, in2334_1, in2334_2, pp41[49]);
    wire[0:0] s2335, in2335_1, in2335_2;
    wire c2335;
    assign in2335_1 = {pp45[45]};
    assign in2335_2 = {pp46[44]};
    Full_Adder FA_2335(s2335, c2335, in2335_1, in2335_2, pp44[46]);
    wire[0:0] s2336, in2336_1, in2336_2;
    wire c2336;
    assign in2336_1 = {pp48[42]};
    assign in2336_2 = {pp49[41]};
    Full_Adder FA_2336(s2336, c2336, in2336_1, in2336_2, pp47[43]);
    wire[0:0] s2337, in2337_1, in2337_2;
    wire c2337;
    assign in2337_1 = {pp51[39]};
    assign in2337_2 = {pp52[38]};
    Full_Adder FA_2337(s2337, c2337, in2337_1, in2337_2, pp50[40]);
    wire[0:0] s2338, in2338_1, in2338_2;
    wire c2338;
    assign in2338_1 = {pp54[36]};
    assign in2338_2 = {pp55[35]};
    Full_Adder FA_2338(s2338, c2338, in2338_1, in2338_2, pp53[37]);
    wire[0:0] s2339, in2339_1, in2339_2;
    wire c2339;
    assign in2339_1 = {pp57[33]};
    assign in2339_2 = {pp58[32]};
    Full_Adder FA_2339(s2339, c2339, in2339_1, in2339_2, pp56[34]);
    wire[0:0] s2340, in2340_1, in2340_2;
    wire c2340;
    assign in2340_1 = {pp60[30]};
    assign in2340_2 = {pp61[29]};
    Full_Adder FA_2340(s2340, c2340, in2340_1, in2340_2, pp59[31]);
    wire[0:0] s2341, in2341_1, in2341_2;
    wire c2341;
    assign in2341_1 = {pp63[27]};
    assign in2341_2 = {pp64[26]};
    Full_Adder FA_2341(s2341, c2341, in2341_1, in2341_2, pp62[28]);
    wire[0:0] s2342, in2342_1, in2342_2;
    wire c2342;
    assign in2342_1 = {pp66[24]};
    assign in2342_2 = {pp67[23]};
    Full_Adder FA_2342(s2342, c2342, in2342_1, in2342_2, pp65[25]);
    wire[0:0] s2343, in2343_1, in2343_2;
    wire c2343;
    assign in2343_1 = {pp69[21]};
    assign in2343_2 = {pp70[20]};
    Full_Adder FA_2343(s2343, c2343, in2343_1, in2343_2, pp68[22]);
    wire[0:0] s2344, in2344_1, in2344_2;
    wire c2344;
    assign in2344_1 = {pp72[18]};
    assign in2344_2 = {pp73[17]};
    Full_Adder FA_2344(s2344, c2344, in2344_1, in2344_2, pp71[19]);
    wire[0:0] s2345, in2345_1, in2345_2;
    wire c2345;
    assign in2345_1 = {pp75[15]};
    assign in2345_2 = {pp76[14]};
    Full_Adder FA_2345(s2345, c2345, in2345_1, in2345_2, pp74[16]);
    wire[0:0] s2346, in2346_1, in2346_2;
    wire c2346;
    assign in2346_1 = {pp78[12]};
    assign in2346_2 = {pp79[11]};
    Full_Adder FA_2346(s2346, c2346, in2346_1, in2346_2, pp77[13]);
    wire[0:0] s2347, in2347_1, in2347_2;
    wire c2347;
    assign in2347_1 = {pp81[9]};
    assign in2347_2 = {pp82[8]};
    Full_Adder FA_2347(s2347, c2347, in2347_1, in2347_2, pp80[10]);
    wire[0:0] s2348, in2348_1, in2348_2;
    wire c2348;
    assign in2348_1 = {pp84[6]};
    assign in2348_2 = {pp85[5]};
    Full_Adder FA_2348(s2348, c2348, in2348_1, in2348_2, pp83[7]);
    wire[0:0] s2349, in2349_1, in2349_2;
    wire c2349;
    assign in2349_1 = {pp87[3]};
    assign in2349_2 = {pp88[2]};
    Full_Adder FA_2349(s2349, c2349, in2349_1, in2349_2, pp86[4]);
    wire[0:0] s2350, in2350_1, in2350_2;
    wire c2350;
    assign in2350_1 = {pp90[0]};
    assign in2350_2 = {c7};
    Full_Adder FA_2350(s2350, c2350, in2350_1, in2350_2, pp89[1]);
    wire[0:0] s2351, in2351_1, in2351_2;
    wire c2351;
    assign in2351_1 = {c9};
    assign in2351_2 = {c10};
    Full_Adder FA_2351(s2351, c2351, in2351_1, in2351_2, c8);
    wire[0:0] s2352, in2352_1, in2352_2;
    wire c2352;
    assign in2352_1 = {s12[0]};
    assign in2352_2 = {s13[0]};
    Full_Adder FA_2352(s2352, c2352, in2352_1, in2352_2, s11[0]);
    wire[0:0] s2353, in2353_1, in2353_2;
    wire c2353;
    assign in2353_1 = {pp18[73]};
    assign in2353_2 = {pp19[72]};
    Full_Adder FA_2353(s2353, c2353, in2353_1, in2353_2, pp17[74]);
    wire[0:0] s2354, in2354_1, in2354_2;
    wire c2354;
    assign in2354_1 = {pp21[70]};
    assign in2354_2 = {pp22[69]};
    Full_Adder FA_2354(s2354, c2354, in2354_1, in2354_2, pp20[71]);
    wire[0:0] s2355, in2355_1, in2355_2;
    wire c2355;
    assign in2355_1 = {pp24[67]};
    assign in2355_2 = {pp25[66]};
    Full_Adder FA_2355(s2355, c2355, in2355_1, in2355_2, pp23[68]);
    wire[0:0] s2356, in2356_1, in2356_2;
    wire c2356;
    assign in2356_1 = {pp27[64]};
    assign in2356_2 = {pp28[63]};
    Full_Adder FA_2356(s2356, c2356, in2356_1, in2356_2, pp26[65]);
    wire[0:0] s2357, in2357_1, in2357_2;
    wire c2357;
    assign in2357_1 = {pp30[61]};
    assign in2357_2 = {pp31[60]};
    Full_Adder FA_2357(s2357, c2357, in2357_1, in2357_2, pp29[62]);
    wire[0:0] s2358, in2358_1, in2358_2;
    wire c2358;
    assign in2358_1 = {pp33[58]};
    assign in2358_2 = {pp34[57]};
    Full_Adder FA_2358(s2358, c2358, in2358_1, in2358_2, pp32[59]);
    wire[0:0] s2359, in2359_1, in2359_2;
    wire c2359;
    assign in2359_1 = {pp36[55]};
    assign in2359_2 = {pp37[54]};
    Full_Adder FA_2359(s2359, c2359, in2359_1, in2359_2, pp35[56]);
    wire[0:0] s2360, in2360_1, in2360_2;
    wire c2360;
    assign in2360_1 = {pp39[52]};
    assign in2360_2 = {pp40[51]};
    Full_Adder FA_2360(s2360, c2360, in2360_1, in2360_2, pp38[53]);
    wire[0:0] s2361, in2361_1, in2361_2;
    wire c2361;
    assign in2361_1 = {pp42[49]};
    assign in2361_2 = {pp43[48]};
    Full_Adder FA_2361(s2361, c2361, in2361_1, in2361_2, pp41[50]);
    wire[0:0] s2362, in2362_1, in2362_2;
    wire c2362;
    assign in2362_1 = {pp45[46]};
    assign in2362_2 = {pp46[45]};
    Full_Adder FA_2362(s2362, c2362, in2362_1, in2362_2, pp44[47]);
    wire[0:0] s2363, in2363_1, in2363_2;
    wire c2363;
    assign in2363_1 = {pp48[43]};
    assign in2363_2 = {pp49[42]};
    Full_Adder FA_2363(s2363, c2363, in2363_1, in2363_2, pp47[44]);
    wire[0:0] s2364, in2364_1, in2364_2;
    wire c2364;
    assign in2364_1 = {pp51[40]};
    assign in2364_2 = {pp52[39]};
    Full_Adder FA_2364(s2364, c2364, in2364_1, in2364_2, pp50[41]);
    wire[0:0] s2365, in2365_1, in2365_2;
    wire c2365;
    assign in2365_1 = {pp54[37]};
    assign in2365_2 = {pp55[36]};
    Full_Adder FA_2365(s2365, c2365, in2365_1, in2365_2, pp53[38]);
    wire[0:0] s2366, in2366_1, in2366_2;
    wire c2366;
    assign in2366_1 = {pp57[34]};
    assign in2366_2 = {pp58[33]};
    Full_Adder FA_2366(s2366, c2366, in2366_1, in2366_2, pp56[35]);
    wire[0:0] s2367, in2367_1, in2367_2;
    wire c2367;
    assign in2367_1 = {pp60[31]};
    assign in2367_2 = {pp61[30]};
    Full_Adder FA_2367(s2367, c2367, in2367_1, in2367_2, pp59[32]);
    wire[0:0] s2368, in2368_1, in2368_2;
    wire c2368;
    assign in2368_1 = {pp63[28]};
    assign in2368_2 = {pp64[27]};
    Full_Adder FA_2368(s2368, c2368, in2368_1, in2368_2, pp62[29]);
    wire[0:0] s2369, in2369_1, in2369_2;
    wire c2369;
    assign in2369_1 = {pp66[25]};
    assign in2369_2 = {pp67[24]};
    Full_Adder FA_2369(s2369, c2369, in2369_1, in2369_2, pp65[26]);
    wire[0:0] s2370, in2370_1, in2370_2;
    wire c2370;
    assign in2370_1 = {pp69[22]};
    assign in2370_2 = {pp70[21]};
    Full_Adder FA_2370(s2370, c2370, in2370_1, in2370_2, pp68[23]);
    wire[0:0] s2371, in2371_1, in2371_2;
    wire c2371;
    assign in2371_1 = {pp72[19]};
    assign in2371_2 = {pp73[18]};
    Full_Adder FA_2371(s2371, c2371, in2371_1, in2371_2, pp71[20]);
    wire[0:0] s2372, in2372_1, in2372_2;
    wire c2372;
    assign in2372_1 = {pp75[16]};
    assign in2372_2 = {pp76[15]};
    Full_Adder FA_2372(s2372, c2372, in2372_1, in2372_2, pp74[17]);
    wire[0:0] s2373, in2373_1, in2373_2;
    wire c2373;
    assign in2373_1 = {pp78[13]};
    assign in2373_2 = {pp79[12]};
    Full_Adder FA_2373(s2373, c2373, in2373_1, in2373_2, pp77[14]);
    wire[0:0] s2374, in2374_1, in2374_2;
    wire c2374;
    assign in2374_1 = {pp81[10]};
    assign in2374_2 = {pp82[9]};
    Full_Adder FA_2374(s2374, c2374, in2374_1, in2374_2, pp80[11]);
    wire[0:0] s2375, in2375_1, in2375_2;
    wire c2375;
    assign in2375_1 = {pp84[7]};
    assign in2375_2 = {pp85[6]};
    Full_Adder FA_2375(s2375, c2375, in2375_1, in2375_2, pp83[8]);
    wire[0:0] s2376, in2376_1, in2376_2;
    wire c2376;
    assign in2376_1 = {pp87[4]};
    assign in2376_2 = {pp88[3]};
    Full_Adder FA_2376(s2376, c2376, in2376_1, in2376_2, pp86[5]);
    wire[0:0] s2377, in2377_1, in2377_2;
    wire c2377;
    assign in2377_1 = {pp90[1]};
    assign in2377_2 = {pp91[0]};
    Full_Adder FA_2377(s2377, c2377, in2377_1, in2377_2, pp89[2]);
    wire[0:0] s2378, in2378_1, in2378_2;
    wire c2378;
    assign in2378_1 = {c12};
    assign in2378_2 = {c13};
    Full_Adder FA_2378(s2378, c2378, in2378_1, in2378_2, c11);
    wire[0:0] s2379, in2379_1, in2379_2;
    wire c2379;
    assign in2379_1 = {c15};
    assign in2379_2 = {s16[0]};
    Full_Adder FA_2379(s2379, c2379, in2379_1, in2379_2, c14);
    wire[0:0] s2380, in2380_1, in2380_2;
    wire c2380;
    assign in2380_1 = {s18[0]};
    assign in2380_2 = {s19[0]};
    Full_Adder FA_2380(s2380, c2380, in2380_1, in2380_2, s17[0]);
    wire[0:0] s2381, in2381_1, in2381_2;
    wire c2381;
    assign in2381_1 = {pp21[71]};
    assign in2381_2 = {pp22[70]};
    Full_Adder FA_2381(s2381, c2381, in2381_1, in2381_2, pp20[72]);
    wire[0:0] s2382, in2382_1, in2382_2;
    wire c2382;
    assign in2382_1 = {pp24[68]};
    assign in2382_2 = {pp25[67]};
    Full_Adder FA_2382(s2382, c2382, in2382_1, in2382_2, pp23[69]);
    wire[0:0] s2383, in2383_1, in2383_2;
    wire c2383;
    assign in2383_1 = {pp27[65]};
    assign in2383_2 = {pp28[64]};
    Full_Adder FA_2383(s2383, c2383, in2383_1, in2383_2, pp26[66]);
    wire[0:0] s2384, in2384_1, in2384_2;
    wire c2384;
    assign in2384_1 = {pp30[62]};
    assign in2384_2 = {pp31[61]};
    Full_Adder FA_2384(s2384, c2384, in2384_1, in2384_2, pp29[63]);
    wire[0:0] s2385, in2385_1, in2385_2;
    wire c2385;
    assign in2385_1 = {pp33[59]};
    assign in2385_2 = {pp34[58]};
    Full_Adder FA_2385(s2385, c2385, in2385_1, in2385_2, pp32[60]);
    wire[0:0] s2386, in2386_1, in2386_2;
    wire c2386;
    assign in2386_1 = {pp36[56]};
    assign in2386_2 = {pp37[55]};
    Full_Adder FA_2386(s2386, c2386, in2386_1, in2386_2, pp35[57]);
    wire[0:0] s2387, in2387_1, in2387_2;
    wire c2387;
    assign in2387_1 = {pp39[53]};
    assign in2387_2 = {pp40[52]};
    Full_Adder FA_2387(s2387, c2387, in2387_1, in2387_2, pp38[54]);
    wire[0:0] s2388, in2388_1, in2388_2;
    wire c2388;
    assign in2388_1 = {pp42[50]};
    assign in2388_2 = {pp43[49]};
    Full_Adder FA_2388(s2388, c2388, in2388_1, in2388_2, pp41[51]);
    wire[0:0] s2389, in2389_1, in2389_2;
    wire c2389;
    assign in2389_1 = {pp45[47]};
    assign in2389_2 = {pp46[46]};
    Full_Adder FA_2389(s2389, c2389, in2389_1, in2389_2, pp44[48]);
    wire[0:0] s2390, in2390_1, in2390_2;
    wire c2390;
    assign in2390_1 = {pp48[44]};
    assign in2390_2 = {pp49[43]};
    Full_Adder FA_2390(s2390, c2390, in2390_1, in2390_2, pp47[45]);
    wire[0:0] s2391, in2391_1, in2391_2;
    wire c2391;
    assign in2391_1 = {pp51[41]};
    assign in2391_2 = {pp52[40]};
    Full_Adder FA_2391(s2391, c2391, in2391_1, in2391_2, pp50[42]);
    wire[0:0] s2392, in2392_1, in2392_2;
    wire c2392;
    assign in2392_1 = {pp54[38]};
    assign in2392_2 = {pp55[37]};
    Full_Adder FA_2392(s2392, c2392, in2392_1, in2392_2, pp53[39]);
    wire[0:0] s2393, in2393_1, in2393_2;
    wire c2393;
    assign in2393_1 = {pp57[35]};
    assign in2393_2 = {pp58[34]};
    Full_Adder FA_2393(s2393, c2393, in2393_1, in2393_2, pp56[36]);
    wire[0:0] s2394, in2394_1, in2394_2;
    wire c2394;
    assign in2394_1 = {pp60[32]};
    assign in2394_2 = {pp61[31]};
    Full_Adder FA_2394(s2394, c2394, in2394_1, in2394_2, pp59[33]);
    wire[0:0] s2395, in2395_1, in2395_2;
    wire c2395;
    assign in2395_1 = {pp63[29]};
    assign in2395_2 = {pp64[28]};
    Full_Adder FA_2395(s2395, c2395, in2395_1, in2395_2, pp62[30]);
    wire[0:0] s2396, in2396_1, in2396_2;
    wire c2396;
    assign in2396_1 = {pp66[26]};
    assign in2396_2 = {pp67[25]};
    Full_Adder FA_2396(s2396, c2396, in2396_1, in2396_2, pp65[27]);
    wire[0:0] s2397, in2397_1, in2397_2;
    wire c2397;
    assign in2397_1 = {pp69[23]};
    assign in2397_2 = {pp70[22]};
    Full_Adder FA_2397(s2397, c2397, in2397_1, in2397_2, pp68[24]);
    wire[0:0] s2398, in2398_1, in2398_2;
    wire c2398;
    assign in2398_1 = {pp72[20]};
    assign in2398_2 = {pp73[19]};
    Full_Adder FA_2398(s2398, c2398, in2398_1, in2398_2, pp71[21]);
    wire[0:0] s2399, in2399_1, in2399_2;
    wire c2399;
    assign in2399_1 = {pp75[17]};
    assign in2399_2 = {pp76[16]};
    Full_Adder FA_2399(s2399, c2399, in2399_1, in2399_2, pp74[18]);
    wire[0:0] s2400, in2400_1, in2400_2;
    wire c2400;
    assign in2400_1 = {pp78[14]};
    assign in2400_2 = {pp79[13]};
    Full_Adder FA_2400(s2400, c2400, in2400_1, in2400_2, pp77[15]);
    wire[0:0] s2401, in2401_1, in2401_2;
    wire c2401;
    assign in2401_1 = {pp81[11]};
    assign in2401_2 = {pp82[10]};
    Full_Adder FA_2401(s2401, c2401, in2401_1, in2401_2, pp80[12]);
    wire[0:0] s2402, in2402_1, in2402_2;
    wire c2402;
    assign in2402_1 = {pp84[8]};
    assign in2402_2 = {pp85[7]};
    Full_Adder FA_2402(s2402, c2402, in2402_1, in2402_2, pp83[9]);
    wire[0:0] s2403, in2403_1, in2403_2;
    wire c2403;
    assign in2403_1 = {pp87[5]};
    assign in2403_2 = {pp88[4]};
    Full_Adder FA_2403(s2403, c2403, in2403_1, in2403_2, pp86[6]);
    wire[0:0] s2404, in2404_1, in2404_2;
    wire c2404;
    assign in2404_1 = {pp90[2]};
    assign in2404_2 = {pp91[1]};
    Full_Adder FA_2404(s2404, c2404, in2404_1, in2404_2, pp89[3]);
    wire[0:0] s2405, in2405_1, in2405_2;
    wire c2405;
    assign in2405_1 = {c16};
    assign in2405_2 = {c17};
    Full_Adder FA_2405(s2405, c2405, in2405_1, in2405_2, pp92[0]);
    wire[0:0] s2406, in2406_1, in2406_2;
    wire c2406;
    assign in2406_1 = {c19};
    assign in2406_2 = {c20};
    Full_Adder FA_2406(s2406, c2406, in2406_1, in2406_2, c18);
    wire[0:0] s2407, in2407_1, in2407_2;
    wire c2407;
    assign in2407_1 = {s22[0]};
    assign in2407_2 = {s23[0]};
    Full_Adder FA_2407(s2407, c2407, in2407_1, in2407_2, c21);
    wire[0:0] s2408, in2408_1, in2408_2;
    wire c2408;
    assign in2408_1 = {s25[0]};
    assign in2408_2 = {s26[0]};
    Full_Adder FA_2408(s2408, c2408, in2408_1, in2408_2, s24[0]);
    wire[0:0] s2409, in2409_1, in2409_2;
    wire c2409;
    assign in2409_1 = {pp24[69]};
    assign in2409_2 = {pp25[68]};
    Full_Adder FA_2409(s2409, c2409, in2409_1, in2409_2, pp23[70]);
    wire[0:0] s2410, in2410_1, in2410_2;
    wire c2410;
    assign in2410_1 = {pp27[66]};
    assign in2410_2 = {pp28[65]};
    Full_Adder FA_2410(s2410, c2410, in2410_1, in2410_2, pp26[67]);
    wire[0:0] s2411, in2411_1, in2411_2;
    wire c2411;
    assign in2411_1 = {pp30[63]};
    assign in2411_2 = {pp31[62]};
    Full_Adder FA_2411(s2411, c2411, in2411_1, in2411_2, pp29[64]);
    wire[0:0] s2412, in2412_1, in2412_2;
    wire c2412;
    assign in2412_1 = {pp33[60]};
    assign in2412_2 = {pp34[59]};
    Full_Adder FA_2412(s2412, c2412, in2412_1, in2412_2, pp32[61]);
    wire[0:0] s2413, in2413_1, in2413_2;
    wire c2413;
    assign in2413_1 = {pp36[57]};
    assign in2413_2 = {pp37[56]};
    Full_Adder FA_2413(s2413, c2413, in2413_1, in2413_2, pp35[58]);
    wire[0:0] s2414, in2414_1, in2414_2;
    wire c2414;
    assign in2414_1 = {pp39[54]};
    assign in2414_2 = {pp40[53]};
    Full_Adder FA_2414(s2414, c2414, in2414_1, in2414_2, pp38[55]);
    wire[0:0] s2415, in2415_1, in2415_2;
    wire c2415;
    assign in2415_1 = {pp42[51]};
    assign in2415_2 = {pp43[50]};
    Full_Adder FA_2415(s2415, c2415, in2415_1, in2415_2, pp41[52]);
    wire[0:0] s2416, in2416_1, in2416_2;
    wire c2416;
    assign in2416_1 = {pp45[48]};
    assign in2416_2 = {pp46[47]};
    Full_Adder FA_2416(s2416, c2416, in2416_1, in2416_2, pp44[49]);
    wire[0:0] s2417, in2417_1, in2417_2;
    wire c2417;
    assign in2417_1 = {pp48[45]};
    assign in2417_2 = {pp49[44]};
    Full_Adder FA_2417(s2417, c2417, in2417_1, in2417_2, pp47[46]);
    wire[0:0] s2418, in2418_1, in2418_2;
    wire c2418;
    assign in2418_1 = {pp51[42]};
    assign in2418_2 = {pp52[41]};
    Full_Adder FA_2418(s2418, c2418, in2418_1, in2418_2, pp50[43]);
    wire[0:0] s2419, in2419_1, in2419_2;
    wire c2419;
    assign in2419_1 = {pp54[39]};
    assign in2419_2 = {pp55[38]};
    Full_Adder FA_2419(s2419, c2419, in2419_1, in2419_2, pp53[40]);
    wire[0:0] s2420, in2420_1, in2420_2;
    wire c2420;
    assign in2420_1 = {pp57[36]};
    assign in2420_2 = {pp58[35]};
    Full_Adder FA_2420(s2420, c2420, in2420_1, in2420_2, pp56[37]);
    wire[0:0] s2421, in2421_1, in2421_2;
    wire c2421;
    assign in2421_1 = {pp60[33]};
    assign in2421_2 = {pp61[32]};
    Full_Adder FA_2421(s2421, c2421, in2421_1, in2421_2, pp59[34]);
    wire[0:0] s2422, in2422_1, in2422_2;
    wire c2422;
    assign in2422_1 = {pp63[30]};
    assign in2422_2 = {pp64[29]};
    Full_Adder FA_2422(s2422, c2422, in2422_1, in2422_2, pp62[31]);
    wire[0:0] s2423, in2423_1, in2423_2;
    wire c2423;
    assign in2423_1 = {pp66[27]};
    assign in2423_2 = {pp67[26]};
    Full_Adder FA_2423(s2423, c2423, in2423_1, in2423_2, pp65[28]);
    wire[0:0] s2424, in2424_1, in2424_2;
    wire c2424;
    assign in2424_1 = {pp69[24]};
    assign in2424_2 = {pp70[23]};
    Full_Adder FA_2424(s2424, c2424, in2424_1, in2424_2, pp68[25]);
    wire[0:0] s2425, in2425_1, in2425_2;
    wire c2425;
    assign in2425_1 = {pp72[21]};
    assign in2425_2 = {pp73[20]};
    Full_Adder FA_2425(s2425, c2425, in2425_1, in2425_2, pp71[22]);
    wire[0:0] s2426, in2426_1, in2426_2;
    wire c2426;
    assign in2426_1 = {pp75[18]};
    assign in2426_2 = {pp76[17]};
    Full_Adder FA_2426(s2426, c2426, in2426_1, in2426_2, pp74[19]);
    wire[0:0] s2427, in2427_1, in2427_2;
    wire c2427;
    assign in2427_1 = {pp78[15]};
    assign in2427_2 = {pp79[14]};
    Full_Adder FA_2427(s2427, c2427, in2427_1, in2427_2, pp77[16]);
    wire[0:0] s2428, in2428_1, in2428_2;
    wire c2428;
    assign in2428_1 = {pp81[12]};
    assign in2428_2 = {pp82[11]};
    Full_Adder FA_2428(s2428, c2428, in2428_1, in2428_2, pp80[13]);
    wire[0:0] s2429, in2429_1, in2429_2;
    wire c2429;
    assign in2429_1 = {pp84[9]};
    assign in2429_2 = {pp85[8]};
    Full_Adder FA_2429(s2429, c2429, in2429_1, in2429_2, pp83[10]);
    wire[0:0] s2430, in2430_1, in2430_2;
    wire c2430;
    assign in2430_1 = {pp87[6]};
    assign in2430_2 = {pp88[5]};
    Full_Adder FA_2430(s2430, c2430, in2430_1, in2430_2, pp86[7]);
    wire[0:0] s2431, in2431_1, in2431_2;
    wire c2431;
    assign in2431_1 = {pp90[3]};
    assign in2431_2 = {pp91[2]};
    Full_Adder FA_2431(s2431, c2431, in2431_1, in2431_2, pp89[4]);
    wire[0:0] s2432, in2432_1, in2432_2;
    wire c2432;
    assign in2432_1 = {pp93[0]};
    assign in2432_2 = {c22};
    Full_Adder FA_2432(s2432, c2432, in2432_1, in2432_2, pp92[1]);
    wire[0:0] s2433, in2433_1, in2433_2;
    wire c2433;
    assign in2433_1 = {c24};
    assign in2433_2 = {c25};
    Full_Adder FA_2433(s2433, c2433, in2433_1, in2433_2, c23);
    wire[0:0] s2434, in2434_1, in2434_2;
    wire c2434;
    assign in2434_1 = {c27};
    assign in2434_2 = {c28};
    Full_Adder FA_2434(s2434, c2434, in2434_1, in2434_2, c26);
    wire[0:0] s2435, in2435_1, in2435_2;
    wire c2435;
    assign in2435_1 = {s30[0]};
    assign in2435_2 = {s31[0]};
    Full_Adder FA_2435(s2435, c2435, in2435_1, in2435_2, s29[0]);
    wire[0:0] s2436, in2436_1, in2436_2;
    wire c2436;
    assign in2436_1 = {s33[0]};
    assign in2436_2 = {s34[0]};
    Full_Adder FA_2436(s2436, c2436, in2436_1, in2436_2, s32[0]);
    wire[0:0] s2437, in2437_1, in2437_2;
    wire c2437;
    assign in2437_1 = {pp27[67]};
    assign in2437_2 = {pp28[66]};
    Full_Adder FA_2437(s2437, c2437, in2437_1, in2437_2, pp26[68]);
    wire[0:0] s2438, in2438_1, in2438_2;
    wire c2438;
    assign in2438_1 = {pp30[64]};
    assign in2438_2 = {pp31[63]};
    Full_Adder FA_2438(s2438, c2438, in2438_1, in2438_2, pp29[65]);
    wire[0:0] s2439, in2439_1, in2439_2;
    wire c2439;
    assign in2439_1 = {pp33[61]};
    assign in2439_2 = {pp34[60]};
    Full_Adder FA_2439(s2439, c2439, in2439_1, in2439_2, pp32[62]);
    wire[0:0] s2440, in2440_1, in2440_2;
    wire c2440;
    assign in2440_1 = {pp36[58]};
    assign in2440_2 = {pp37[57]};
    Full_Adder FA_2440(s2440, c2440, in2440_1, in2440_2, pp35[59]);
    wire[0:0] s2441, in2441_1, in2441_2;
    wire c2441;
    assign in2441_1 = {pp39[55]};
    assign in2441_2 = {pp40[54]};
    Full_Adder FA_2441(s2441, c2441, in2441_1, in2441_2, pp38[56]);
    wire[0:0] s2442, in2442_1, in2442_2;
    wire c2442;
    assign in2442_1 = {pp42[52]};
    assign in2442_2 = {pp43[51]};
    Full_Adder FA_2442(s2442, c2442, in2442_1, in2442_2, pp41[53]);
    wire[0:0] s2443, in2443_1, in2443_2;
    wire c2443;
    assign in2443_1 = {pp45[49]};
    assign in2443_2 = {pp46[48]};
    Full_Adder FA_2443(s2443, c2443, in2443_1, in2443_2, pp44[50]);
    wire[0:0] s2444, in2444_1, in2444_2;
    wire c2444;
    assign in2444_1 = {pp48[46]};
    assign in2444_2 = {pp49[45]};
    Full_Adder FA_2444(s2444, c2444, in2444_1, in2444_2, pp47[47]);
    wire[0:0] s2445, in2445_1, in2445_2;
    wire c2445;
    assign in2445_1 = {pp51[43]};
    assign in2445_2 = {pp52[42]};
    Full_Adder FA_2445(s2445, c2445, in2445_1, in2445_2, pp50[44]);
    wire[0:0] s2446, in2446_1, in2446_2;
    wire c2446;
    assign in2446_1 = {pp54[40]};
    assign in2446_2 = {pp55[39]};
    Full_Adder FA_2446(s2446, c2446, in2446_1, in2446_2, pp53[41]);
    wire[0:0] s2447, in2447_1, in2447_2;
    wire c2447;
    assign in2447_1 = {pp57[37]};
    assign in2447_2 = {pp58[36]};
    Full_Adder FA_2447(s2447, c2447, in2447_1, in2447_2, pp56[38]);
    wire[0:0] s2448, in2448_1, in2448_2;
    wire c2448;
    assign in2448_1 = {pp60[34]};
    assign in2448_2 = {pp61[33]};
    Full_Adder FA_2448(s2448, c2448, in2448_1, in2448_2, pp59[35]);
    wire[0:0] s2449, in2449_1, in2449_2;
    wire c2449;
    assign in2449_1 = {pp63[31]};
    assign in2449_2 = {pp64[30]};
    Full_Adder FA_2449(s2449, c2449, in2449_1, in2449_2, pp62[32]);
    wire[0:0] s2450, in2450_1, in2450_2;
    wire c2450;
    assign in2450_1 = {pp66[28]};
    assign in2450_2 = {pp67[27]};
    Full_Adder FA_2450(s2450, c2450, in2450_1, in2450_2, pp65[29]);
    wire[0:0] s2451, in2451_1, in2451_2;
    wire c2451;
    assign in2451_1 = {pp69[25]};
    assign in2451_2 = {pp70[24]};
    Full_Adder FA_2451(s2451, c2451, in2451_1, in2451_2, pp68[26]);
    wire[0:0] s2452, in2452_1, in2452_2;
    wire c2452;
    assign in2452_1 = {pp72[22]};
    assign in2452_2 = {pp73[21]};
    Full_Adder FA_2452(s2452, c2452, in2452_1, in2452_2, pp71[23]);
    wire[0:0] s2453, in2453_1, in2453_2;
    wire c2453;
    assign in2453_1 = {pp75[19]};
    assign in2453_2 = {pp76[18]};
    Full_Adder FA_2453(s2453, c2453, in2453_1, in2453_2, pp74[20]);
    wire[0:0] s2454, in2454_1, in2454_2;
    wire c2454;
    assign in2454_1 = {pp78[16]};
    assign in2454_2 = {pp79[15]};
    Full_Adder FA_2454(s2454, c2454, in2454_1, in2454_2, pp77[17]);
    wire[0:0] s2455, in2455_1, in2455_2;
    wire c2455;
    assign in2455_1 = {pp81[13]};
    assign in2455_2 = {pp82[12]};
    Full_Adder FA_2455(s2455, c2455, in2455_1, in2455_2, pp80[14]);
    wire[0:0] s2456, in2456_1, in2456_2;
    wire c2456;
    assign in2456_1 = {pp84[10]};
    assign in2456_2 = {pp85[9]};
    Full_Adder FA_2456(s2456, c2456, in2456_1, in2456_2, pp83[11]);
    wire[0:0] s2457, in2457_1, in2457_2;
    wire c2457;
    assign in2457_1 = {pp87[7]};
    assign in2457_2 = {pp88[6]};
    Full_Adder FA_2457(s2457, c2457, in2457_1, in2457_2, pp86[8]);
    wire[0:0] s2458, in2458_1, in2458_2;
    wire c2458;
    assign in2458_1 = {pp90[4]};
    assign in2458_2 = {pp91[3]};
    Full_Adder FA_2458(s2458, c2458, in2458_1, in2458_2, pp89[5]);
    wire[0:0] s2459, in2459_1, in2459_2;
    wire c2459;
    assign in2459_1 = {pp93[1]};
    assign in2459_2 = {pp94[0]};
    Full_Adder FA_2459(s2459, c2459, in2459_1, in2459_2, pp92[2]);
    wire[0:0] s2460, in2460_1, in2460_2;
    wire c2460;
    assign in2460_1 = {c30};
    assign in2460_2 = {c31};
    Full_Adder FA_2460(s2460, c2460, in2460_1, in2460_2, c29);
    wire[0:0] s2461, in2461_1, in2461_2;
    wire c2461;
    assign in2461_1 = {c33};
    assign in2461_2 = {c34};
    Full_Adder FA_2461(s2461, c2461, in2461_1, in2461_2, c32);
    wire[0:0] s2462, in2462_1, in2462_2;
    wire c2462;
    assign in2462_1 = {c36};
    assign in2462_2 = {s37[0]};
    Full_Adder FA_2462(s2462, c2462, in2462_1, in2462_2, c35);
    wire[0:0] s2463, in2463_1, in2463_2;
    wire c2463;
    assign in2463_1 = {s39[0]};
    assign in2463_2 = {s40[0]};
    Full_Adder FA_2463(s2463, c2463, in2463_1, in2463_2, s38[0]);
    wire[0:0] s2464, in2464_1, in2464_2;
    wire c2464;
    assign in2464_1 = {s42[0]};
    assign in2464_2 = {s43[0]};
    Full_Adder FA_2464(s2464, c2464, in2464_1, in2464_2, s41[0]);
    wire[0:0] s2465, in2465_1, in2465_2;
    wire c2465;
    assign in2465_1 = {pp30[65]};
    assign in2465_2 = {pp31[64]};
    Full_Adder FA_2465(s2465, c2465, in2465_1, in2465_2, pp29[66]);
    wire[0:0] s2466, in2466_1, in2466_2;
    wire c2466;
    assign in2466_1 = {pp33[62]};
    assign in2466_2 = {pp34[61]};
    Full_Adder FA_2466(s2466, c2466, in2466_1, in2466_2, pp32[63]);
    wire[0:0] s2467, in2467_1, in2467_2;
    wire c2467;
    assign in2467_1 = {pp36[59]};
    assign in2467_2 = {pp37[58]};
    Full_Adder FA_2467(s2467, c2467, in2467_1, in2467_2, pp35[60]);
    wire[0:0] s2468, in2468_1, in2468_2;
    wire c2468;
    assign in2468_1 = {pp39[56]};
    assign in2468_2 = {pp40[55]};
    Full_Adder FA_2468(s2468, c2468, in2468_1, in2468_2, pp38[57]);
    wire[0:0] s2469, in2469_1, in2469_2;
    wire c2469;
    assign in2469_1 = {pp42[53]};
    assign in2469_2 = {pp43[52]};
    Full_Adder FA_2469(s2469, c2469, in2469_1, in2469_2, pp41[54]);
    wire[0:0] s2470, in2470_1, in2470_2;
    wire c2470;
    assign in2470_1 = {pp45[50]};
    assign in2470_2 = {pp46[49]};
    Full_Adder FA_2470(s2470, c2470, in2470_1, in2470_2, pp44[51]);
    wire[0:0] s2471, in2471_1, in2471_2;
    wire c2471;
    assign in2471_1 = {pp48[47]};
    assign in2471_2 = {pp49[46]};
    Full_Adder FA_2471(s2471, c2471, in2471_1, in2471_2, pp47[48]);
    wire[0:0] s2472, in2472_1, in2472_2;
    wire c2472;
    assign in2472_1 = {pp51[44]};
    assign in2472_2 = {pp52[43]};
    Full_Adder FA_2472(s2472, c2472, in2472_1, in2472_2, pp50[45]);
    wire[0:0] s2473, in2473_1, in2473_2;
    wire c2473;
    assign in2473_1 = {pp54[41]};
    assign in2473_2 = {pp55[40]};
    Full_Adder FA_2473(s2473, c2473, in2473_1, in2473_2, pp53[42]);
    wire[0:0] s2474, in2474_1, in2474_2;
    wire c2474;
    assign in2474_1 = {pp57[38]};
    assign in2474_2 = {pp58[37]};
    Full_Adder FA_2474(s2474, c2474, in2474_1, in2474_2, pp56[39]);
    wire[0:0] s2475, in2475_1, in2475_2;
    wire c2475;
    assign in2475_1 = {pp60[35]};
    assign in2475_2 = {pp61[34]};
    Full_Adder FA_2475(s2475, c2475, in2475_1, in2475_2, pp59[36]);
    wire[0:0] s2476, in2476_1, in2476_2;
    wire c2476;
    assign in2476_1 = {pp63[32]};
    assign in2476_2 = {pp64[31]};
    Full_Adder FA_2476(s2476, c2476, in2476_1, in2476_2, pp62[33]);
    wire[0:0] s2477, in2477_1, in2477_2;
    wire c2477;
    assign in2477_1 = {pp66[29]};
    assign in2477_2 = {pp67[28]};
    Full_Adder FA_2477(s2477, c2477, in2477_1, in2477_2, pp65[30]);
    wire[0:0] s2478, in2478_1, in2478_2;
    wire c2478;
    assign in2478_1 = {pp69[26]};
    assign in2478_2 = {pp70[25]};
    Full_Adder FA_2478(s2478, c2478, in2478_1, in2478_2, pp68[27]);
    wire[0:0] s2479, in2479_1, in2479_2;
    wire c2479;
    assign in2479_1 = {pp72[23]};
    assign in2479_2 = {pp73[22]};
    Full_Adder FA_2479(s2479, c2479, in2479_1, in2479_2, pp71[24]);
    wire[0:0] s2480, in2480_1, in2480_2;
    wire c2480;
    assign in2480_1 = {pp75[20]};
    assign in2480_2 = {pp76[19]};
    Full_Adder FA_2480(s2480, c2480, in2480_1, in2480_2, pp74[21]);
    wire[0:0] s2481, in2481_1, in2481_2;
    wire c2481;
    assign in2481_1 = {pp78[17]};
    assign in2481_2 = {pp79[16]};
    Full_Adder FA_2481(s2481, c2481, in2481_1, in2481_2, pp77[18]);
    wire[0:0] s2482, in2482_1, in2482_2;
    wire c2482;
    assign in2482_1 = {pp81[14]};
    assign in2482_2 = {pp82[13]};
    Full_Adder FA_2482(s2482, c2482, in2482_1, in2482_2, pp80[15]);
    wire[0:0] s2483, in2483_1, in2483_2;
    wire c2483;
    assign in2483_1 = {pp84[11]};
    assign in2483_2 = {pp85[10]};
    Full_Adder FA_2483(s2483, c2483, in2483_1, in2483_2, pp83[12]);
    wire[0:0] s2484, in2484_1, in2484_2;
    wire c2484;
    assign in2484_1 = {pp87[8]};
    assign in2484_2 = {pp88[7]};
    Full_Adder FA_2484(s2484, c2484, in2484_1, in2484_2, pp86[9]);
    wire[0:0] s2485, in2485_1, in2485_2;
    wire c2485;
    assign in2485_1 = {pp90[5]};
    assign in2485_2 = {pp91[4]};
    Full_Adder FA_2485(s2485, c2485, in2485_1, in2485_2, pp89[6]);
    wire[0:0] s2486, in2486_1, in2486_2;
    wire c2486;
    assign in2486_1 = {pp93[2]};
    assign in2486_2 = {pp94[1]};
    Full_Adder FA_2486(s2486, c2486, in2486_1, in2486_2, pp92[3]);
    wire[0:0] s2487, in2487_1, in2487_2;
    wire c2487;
    assign in2487_1 = {c37};
    assign in2487_2 = {c38};
    Full_Adder FA_2487(s2487, c2487, in2487_1, in2487_2, pp95[0]);
    wire[0:0] s2488, in2488_1, in2488_2;
    wire c2488;
    assign in2488_1 = {c40};
    assign in2488_2 = {c41};
    Full_Adder FA_2488(s2488, c2488, in2488_1, in2488_2, c39);
    wire[0:0] s2489, in2489_1, in2489_2;
    wire c2489;
    assign in2489_1 = {c43};
    assign in2489_2 = {c44};
    Full_Adder FA_2489(s2489, c2489, in2489_1, in2489_2, c42);
    wire[0:0] s2490, in2490_1, in2490_2;
    wire c2490;
    assign in2490_1 = {s46[0]};
    assign in2490_2 = {s47[0]};
    Full_Adder FA_2490(s2490, c2490, in2490_1, in2490_2, c45);
    wire[0:0] s2491, in2491_1, in2491_2;
    wire c2491;
    assign in2491_1 = {s49[0]};
    assign in2491_2 = {s50[0]};
    Full_Adder FA_2491(s2491, c2491, in2491_1, in2491_2, s48[0]);
    wire[0:0] s2492, in2492_1, in2492_2;
    wire c2492;
    assign in2492_1 = {s52[0]};
    assign in2492_2 = {s53[0]};
    Full_Adder FA_2492(s2492, c2492, in2492_1, in2492_2, s51[0]);
    wire[0:0] s2493, in2493_1, in2493_2;
    wire c2493;
    assign in2493_1 = {pp33[63]};
    assign in2493_2 = {pp34[62]};
    Full_Adder FA_2493(s2493, c2493, in2493_1, in2493_2, pp32[64]);
    wire[0:0] s2494, in2494_1, in2494_2;
    wire c2494;
    assign in2494_1 = {pp36[60]};
    assign in2494_2 = {pp37[59]};
    Full_Adder FA_2494(s2494, c2494, in2494_1, in2494_2, pp35[61]);
    wire[0:0] s2495, in2495_1, in2495_2;
    wire c2495;
    assign in2495_1 = {pp39[57]};
    assign in2495_2 = {pp40[56]};
    Full_Adder FA_2495(s2495, c2495, in2495_1, in2495_2, pp38[58]);
    wire[0:0] s2496, in2496_1, in2496_2;
    wire c2496;
    assign in2496_1 = {pp42[54]};
    assign in2496_2 = {pp43[53]};
    Full_Adder FA_2496(s2496, c2496, in2496_1, in2496_2, pp41[55]);
    wire[0:0] s2497, in2497_1, in2497_2;
    wire c2497;
    assign in2497_1 = {pp45[51]};
    assign in2497_2 = {pp46[50]};
    Full_Adder FA_2497(s2497, c2497, in2497_1, in2497_2, pp44[52]);
    wire[0:0] s2498, in2498_1, in2498_2;
    wire c2498;
    assign in2498_1 = {pp48[48]};
    assign in2498_2 = {pp49[47]};
    Full_Adder FA_2498(s2498, c2498, in2498_1, in2498_2, pp47[49]);
    wire[0:0] s2499, in2499_1, in2499_2;
    wire c2499;
    assign in2499_1 = {pp51[45]};
    assign in2499_2 = {pp52[44]};
    Full_Adder FA_2499(s2499, c2499, in2499_1, in2499_2, pp50[46]);
    wire[0:0] s2500, in2500_1, in2500_2;
    wire c2500;
    assign in2500_1 = {pp54[42]};
    assign in2500_2 = {pp55[41]};
    Full_Adder FA_2500(s2500, c2500, in2500_1, in2500_2, pp53[43]);
    wire[0:0] s2501, in2501_1, in2501_2;
    wire c2501;
    assign in2501_1 = {pp57[39]};
    assign in2501_2 = {pp58[38]};
    Full_Adder FA_2501(s2501, c2501, in2501_1, in2501_2, pp56[40]);
    wire[0:0] s2502, in2502_1, in2502_2;
    wire c2502;
    assign in2502_1 = {pp60[36]};
    assign in2502_2 = {pp61[35]};
    Full_Adder FA_2502(s2502, c2502, in2502_1, in2502_2, pp59[37]);
    wire[0:0] s2503, in2503_1, in2503_2;
    wire c2503;
    assign in2503_1 = {pp63[33]};
    assign in2503_2 = {pp64[32]};
    Full_Adder FA_2503(s2503, c2503, in2503_1, in2503_2, pp62[34]);
    wire[0:0] s2504, in2504_1, in2504_2;
    wire c2504;
    assign in2504_1 = {pp66[30]};
    assign in2504_2 = {pp67[29]};
    Full_Adder FA_2504(s2504, c2504, in2504_1, in2504_2, pp65[31]);
    wire[0:0] s2505, in2505_1, in2505_2;
    wire c2505;
    assign in2505_1 = {pp69[27]};
    assign in2505_2 = {pp70[26]};
    Full_Adder FA_2505(s2505, c2505, in2505_1, in2505_2, pp68[28]);
    wire[0:0] s2506, in2506_1, in2506_2;
    wire c2506;
    assign in2506_1 = {pp72[24]};
    assign in2506_2 = {pp73[23]};
    Full_Adder FA_2506(s2506, c2506, in2506_1, in2506_2, pp71[25]);
    wire[0:0] s2507, in2507_1, in2507_2;
    wire c2507;
    assign in2507_1 = {pp75[21]};
    assign in2507_2 = {pp76[20]};
    Full_Adder FA_2507(s2507, c2507, in2507_1, in2507_2, pp74[22]);
    wire[0:0] s2508, in2508_1, in2508_2;
    wire c2508;
    assign in2508_1 = {pp78[18]};
    assign in2508_2 = {pp79[17]};
    Full_Adder FA_2508(s2508, c2508, in2508_1, in2508_2, pp77[19]);
    wire[0:0] s2509, in2509_1, in2509_2;
    wire c2509;
    assign in2509_1 = {pp81[15]};
    assign in2509_2 = {pp82[14]};
    Full_Adder FA_2509(s2509, c2509, in2509_1, in2509_2, pp80[16]);
    wire[0:0] s2510, in2510_1, in2510_2;
    wire c2510;
    assign in2510_1 = {pp84[12]};
    assign in2510_2 = {pp85[11]};
    Full_Adder FA_2510(s2510, c2510, in2510_1, in2510_2, pp83[13]);
    wire[0:0] s2511, in2511_1, in2511_2;
    wire c2511;
    assign in2511_1 = {pp87[9]};
    assign in2511_2 = {pp88[8]};
    Full_Adder FA_2511(s2511, c2511, in2511_1, in2511_2, pp86[10]);
    wire[0:0] s2512, in2512_1, in2512_2;
    wire c2512;
    assign in2512_1 = {pp90[6]};
    assign in2512_2 = {pp91[5]};
    Full_Adder FA_2512(s2512, c2512, in2512_1, in2512_2, pp89[7]);
    wire[0:0] s2513, in2513_1, in2513_2;
    wire c2513;
    assign in2513_1 = {pp93[3]};
    assign in2513_2 = {pp94[2]};
    Full_Adder FA_2513(s2513, c2513, in2513_1, in2513_2, pp92[4]);
    wire[0:0] s2514, in2514_1, in2514_2;
    wire c2514;
    assign in2514_1 = {pp96[0]};
    assign in2514_2 = {c46};
    Full_Adder FA_2514(s2514, c2514, in2514_1, in2514_2, pp95[1]);
    wire[0:0] s2515, in2515_1, in2515_2;
    wire c2515;
    assign in2515_1 = {c48};
    assign in2515_2 = {c49};
    Full_Adder FA_2515(s2515, c2515, in2515_1, in2515_2, c47);
    wire[0:0] s2516, in2516_1, in2516_2;
    wire c2516;
    assign in2516_1 = {c51};
    assign in2516_2 = {c52};
    Full_Adder FA_2516(s2516, c2516, in2516_1, in2516_2, c50);
    wire[0:0] s2517, in2517_1, in2517_2;
    wire c2517;
    assign in2517_1 = {c54};
    assign in2517_2 = {c55};
    Full_Adder FA_2517(s2517, c2517, in2517_1, in2517_2, c53);
    wire[0:0] s2518, in2518_1, in2518_2;
    wire c2518;
    assign in2518_1 = {s57[0]};
    assign in2518_2 = {s58[0]};
    Full_Adder FA_2518(s2518, c2518, in2518_1, in2518_2, s56[0]);
    wire[0:0] s2519, in2519_1, in2519_2;
    wire c2519;
    assign in2519_1 = {s60[0]};
    assign in2519_2 = {s61[0]};
    Full_Adder FA_2519(s2519, c2519, in2519_1, in2519_2, s59[0]);
    wire[0:0] s2520, in2520_1, in2520_2;
    wire c2520;
    assign in2520_1 = {s63[0]};
    assign in2520_2 = {s64[0]};
    Full_Adder FA_2520(s2520, c2520, in2520_1, in2520_2, s62[0]);
    wire[0:0] s2521, in2521_1, in2521_2;
    wire c2521;
    assign in2521_1 = {pp36[61]};
    assign in2521_2 = {pp37[60]};
    Full_Adder FA_2521(s2521, c2521, in2521_1, in2521_2, pp35[62]);
    wire[0:0] s2522, in2522_1, in2522_2;
    wire c2522;
    assign in2522_1 = {pp39[58]};
    assign in2522_2 = {pp40[57]};
    Full_Adder FA_2522(s2522, c2522, in2522_1, in2522_2, pp38[59]);
    wire[0:0] s2523, in2523_1, in2523_2;
    wire c2523;
    assign in2523_1 = {pp42[55]};
    assign in2523_2 = {pp43[54]};
    Full_Adder FA_2523(s2523, c2523, in2523_1, in2523_2, pp41[56]);
    wire[0:0] s2524, in2524_1, in2524_2;
    wire c2524;
    assign in2524_1 = {pp45[52]};
    assign in2524_2 = {pp46[51]};
    Full_Adder FA_2524(s2524, c2524, in2524_1, in2524_2, pp44[53]);
    wire[0:0] s2525, in2525_1, in2525_2;
    wire c2525;
    assign in2525_1 = {pp48[49]};
    assign in2525_2 = {pp49[48]};
    Full_Adder FA_2525(s2525, c2525, in2525_1, in2525_2, pp47[50]);
    wire[0:0] s2526, in2526_1, in2526_2;
    wire c2526;
    assign in2526_1 = {pp51[46]};
    assign in2526_2 = {pp52[45]};
    Full_Adder FA_2526(s2526, c2526, in2526_1, in2526_2, pp50[47]);
    wire[0:0] s2527, in2527_1, in2527_2;
    wire c2527;
    assign in2527_1 = {pp54[43]};
    assign in2527_2 = {pp55[42]};
    Full_Adder FA_2527(s2527, c2527, in2527_1, in2527_2, pp53[44]);
    wire[0:0] s2528, in2528_1, in2528_2;
    wire c2528;
    assign in2528_1 = {pp57[40]};
    assign in2528_2 = {pp58[39]};
    Full_Adder FA_2528(s2528, c2528, in2528_1, in2528_2, pp56[41]);
    wire[0:0] s2529, in2529_1, in2529_2;
    wire c2529;
    assign in2529_1 = {pp60[37]};
    assign in2529_2 = {pp61[36]};
    Full_Adder FA_2529(s2529, c2529, in2529_1, in2529_2, pp59[38]);
    wire[0:0] s2530, in2530_1, in2530_2;
    wire c2530;
    assign in2530_1 = {pp63[34]};
    assign in2530_2 = {pp64[33]};
    Full_Adder FA_2530(s2530, c2530, in2530_1, in2530_2, pp62[35]);
    wire[0:0] s2531, in2531_1, in2531_2;
    wire c2531;
    assign in2531_1 = {pp66[31]};
    assign in2531_2 = {pp67[30]};
    Full_Adder FA_2531(s2531, c2531, in2531_1, in2531_2, pp65[32]);
    wire[0:0] s2532, in2532_1, in2532_2;
    wire c2532;
    assign in2532_1 = {pp69[28]};
    assign in2532_2 = {pp70[27]};
    Full_Adder FA_2532(s2532, c2532, in2532_1, in2532_2, pp68[29]);
    wire[0:0] s2533, in2533_1, in2533_2;
    wire c2533;
    assign in2533_1 = {pp72[25]};
    assign in2533_2 = {pp73[24]};
    Full_Adder FA_2533(s2533, c2533, in2533_1, in2533_2, pp71[26]);
    wire[0:0] s2534, in2534_1, in2534_2;
    wire c2534;
    assign in2534_1 = {pp75[22]};
    assign in2534_2 = {pp76[21]};
    Full_Adder FA_2534(s2534, c2534, in2534_1, in2534_2, pp74[23]);
    wire[0:0] s2535, in2535_1, in2535_2;
    wire c2535;
    assign in2535_1 = {pp78[19]};
    assign in2535_2 = {pp79[18]};
    Full_Adder FA_2535(s2535, c2535, in2535_1, in2535_2, pp77[20]);
    wire[0:0] s2536, in2536_1, in2536_2;
    wire c2536;
    assign in2536_1 = {pp81[16]};
    assign in2536_2 = {pp82[15]};
    Full_Adder FA_2536(s2536, c2536, in2536_1, in2536_2, pp80[17]);
    wire[0:0] s2537, in2537_1, in2537_2;
    wire c2537;
    assign in2537_1 = {pp84[13]};
    assign in2537_2 = {pp85[12]};
    Full_Adder FA_2537(s2537, c2537, in2537_1, in2537_2, pp83[14]);
    wire[0:0] s2538, in2538_1, in2538_2;
    wire c2538;
    assign in2538_1 = {pp87[10]};
    assign in2538_2 = {pp88[9]};
    Full_Adder FA_2538(s2538, c2538, in2538_1, in2538_2, pp86[11]);
    wire[0:0] s2539, in2539_1, in2539_2;
    wire c2539;
    assign in2539_1 = {pp90[7]};
    assign in2539_2 = {pp91[6]};
    Full_Adder FA_2539(s2539, c2539, in2539_1, in2539_2, pp89[8]);
    wire[0:0] s2540, in2540_1, in2540_2;
    wire c2540;
    assign in2540_1 = {pp93[4]};
    assign in2540_2 = {pp94[3]};
    Full_Adder FA_2540(s2540, c2540, in2540_1, in2540_2, pp92[5]);
    wire[0:0] s2541, in2541_1, in2541_2;
    wire c2541;
    assign in2541_1 = {pp96[1]};
    assign in2541_2 = {pp97[0]};
    Full_Adder FA_2541(s2541, c2541, in2541_1, in2541_2, pp95[2]);
    wire[0:0] s2542, in2542_1, in2542_2;
    wire c2542;
    assign in2542_1 = {c57};
    assign in2542_2 = {c58};
    Full_Adder FA_2542(s2542, c2542, in2542_1, in2542_2, c56);
    wire[0:0] s2543, in2543_1, in2543_2;
    wire c2543;
    assign in2543_1 = {c60};
    assign in2543_2 = {c61};
    Full_Adder FA_2543(s2543, c2543, in2543_1, in2543_2, c59);
    wire[0:0] s2544, in2544_1, in2544_2;
    wire c2544;
    assign in2544_1 = {c63};
    assign in2544_2 = {c64};
    Full_Adder FA_2544(s2544, c2544, in2544_1, in2544_2, c62);
    wire[0:0] s2545, in2545_1, in2545_2;
    wire c2545;
    assign in2545_1 = {c66};
    assign in2545_2 = {s67[0]};
    Full_Adder FA_2545(s2545, c2545, in2545_1, in2545_2, c65);
    wire[0:0] s2546, in2546_1, in2546_2;
    wire c2546;
    assign in2546_1 = {s69[0]};
    assign in2546_2 = {s70[0]};
    Full_Adder FA_2546(s2546, c2546, in2546_1, in2546_2, s68[0]);
    wire[0:0] s2547, in2547_1, in2547_2;
    wire c2547;
    assign in2547_1 = {s72[0]};
    assign in2547_2 = {s73[0]};
    Full_Adder FA_2547(s2547, c2547, in2547_1, in2547_2, s71[0]);
    wire[0:0] s2548, in2548_1, in2548_2;
    wire c2548;
    assign in2548_1 = {s75[0]};
    assign in2548_2 = {s76[0]};
    Full_Adder FA_2548(s2548, c2548, in2548_1, in2548_2, s74[0]);
    wire[0:0] s2549, in2549_1, in2549_2;
    wire c2549;
    assign in2549_1 = {pp39[59]};
    assign in2549_2 = {pp40[58]};
    Full_Adder FA_2549(s2549, c2549, in2549_1, in2549_2, pp38[60]);
    wire[0:0] s2550, in2550_1, in2550_2;
    wire c2550;
    assign in2550_1 = {pp42[56]};
    assign in2550_2 = {pp43[55]};
    Full_Adder FA_2550(s2550, c2550, in2550_1, in2550_2, pp41[57]);
    wire[0:0] s2551, in2551_1, in2551_2;
    wire c2551;
    assign in2551_1 = {pp45[53]};
    assign in2551_2 = {pp46[52]};
    Full_Adder FA_2551(s2551, c2551, in2551_1, in2551_2, pp44[54]);
    wire[0:0] s2552, in2552_1, in2552_2;
    wire c2552;
    assign in2552_1 = {pp48[50]};
    assign in2552_2 = {pp49[49]};
    Full_Adder FA_2552(s2552, c2552, in2552_1, in2552_2, pp47[51]);
    wire[0:0] s2553, in2553_1, in2553_2;
    wire c2553;
    assign in2553_1 = {pp51[47]};
    assign in2553_2 = {pp52[46]};
    Full_Adder FA_2553(s2553, c2553, in2553_1, in2553_2, pp50[48]);
    wire[0:0] s2554, in2554_1, in2554_2;
    wire c2554;
    assign in2554_1 = {pp54[44]};
    assign in2554_2 = {pp55[43]};
    Full_Adder FA_2554(s2554, c2554, in2554_1, in2554_2, pp53[45]);
    wire[0:0] s2555, in2555_1, in2555_2;
    wire c2555;
    assign in2555_1 = {pp57[41]};
    assign in2555_2 = {pp58[40]};
    Full_Adder FA_2555(s2555, c2555, in2555_1, in2555_2, pp56[42]);
    wire[0:0] s2556, in2556_1, in2556_2;
    wire c2556;
    assign in2556_1 = {pp60[38]};
    assign in2556_2 = {pp61[37]};
    Full_Adder FA_2556(s2556, c2556, in2556_1, in2556_2, pp59[39]);
    wire[0:0] s2557, in2557_1, in2557_2;
    wire c2557;
    assign in2557_1 = {pp63[35]};
    assign in2557_2 = {pp64[34]};
    Full_Adder FA_2557(s2557, c2557, in2557_1, in2557_2, pp62[36]);
    wire[0:0] s2558, in2558_1, in2558_2;
    wire c2558;
    assign in2558_1 = {pp66[32]};
    assign in2558_2 = {pp67[31]};
    Full_Adder FA_2558(s2558, c2558, in2558_1, in2558_2, pp65[33]);
    wire[0:0] s2559, in2559_1, in2559_2;
    wire c2559;
    assign in2559_1 = {pp69[29]};
    assign in2559_2 = {pp70[28]};
    Full_Adder FA_2559(s2559, c2559, in2559_1, in2559_2, pp68[30]);
    wire[0:0] s2560, in2560_1, in2560_2;
    wire c2560;
    assign in2560_1 = {pp72[26]};
    assign in2560_2 = {pp73[25]};
    Full_Adder FA_2560(s2560, c2560, in2560_1, in2560_2, pp71[27]);
    wire[0:0] s2561, in2561_1, in2561_2;
    wire c2561;
    assign in2561_1 = {pp75[23]};
    assign in2561_2 = {pp76[22]};
    Full_Adder FA_2561(s2561, c2561, in2561_1, in2561_2, pp74[24]);
    wire[0:0] s2562, in2562_1, in2562_2;
    wire c2562;
    assign in2562_1 = {pp78[20]};
    assign in2562_2 = {pp79[19]};
    Full_Adder FA_2562(s2562, c2562, in2562_1, in2562_2, pp77[21]);
    wire[0:0] s2563, in2563_1, in2563_2;
    wire c2563;
    assign in2563_1 = {pp81[17]};
    assign in2563_2 = {pp82[16]};
    Full_Adder FA_2563(s2563, c2563, in2563_1, in2563_2, pp80[18]);
    wire[0:0] s2564, in2564_1, in2564_2;
    wire c2564;
    assign in2564_1 = {pp84[14]};
    assign in2564_2 = {pp85[13]};
    Full_Adder FA_2564(s2564, c2564, in2564_1, in2564_2, pp83[15]);
    wire[0:0] s2565, in2565_1, in2565_2;
    wire c2565;
    assign in2565_1 = {pp87[11]};
    assign in2565_2 = {pp88[10]};
    Full_Adder FA_2565(s2565, c2565, in2565_1, in2565_2, pp86[12]);
    wire[0:0] s2566, in2566_1, in2566_2;
    wire c2566;
    assign in2566_1 = {pp90[8]};
    assign in2566_2 = {pp91[7]};
    Full_Adder FA_2566(s2566, c2566, in2566_1, in2566_2, pp89[9]);
    wire[0:0] s2567, in2567_1, in2567_2;
    wire c2567;
    assign in2567_1 = {pp93[5]};
    assign in2567_2 = {pp94[4]};
    Full_Adder FA_2567(s2567, c2567, in2567_1, in2567_2, pp92[6]);
    wire[0:0] s2568, in2568_1, in2568_2;
    wire c2568;
    assign in2568_1 = {pp96[2]};
    assign in2568_2 = {pp97[1]};
    Full_Adder FA_2568(s2568, c2568, in2568_1, in2568_2, pp95[3]);
    wire[0:0] s2569, in2569_1, in2569_2;
    wire c2569;
    assign in2569_1 = {c67};
    assign in2569_2 = {c68};
    Full_Adder FA_2569(s2569, c2569, in2569_1, in2569_2, pp98[0]);
    wire[0:0] s2570, in2570_1, in2570_2;
    wire c2570;
    assign in2570_1 = {c70};
    assign in2570_2 = {c71};
    Full_Adder FA_2570(s2570, c2570, in2570_1, in2570_2, c69);
    wire[0:0] s2571, in2571_1, in2571_2;
    wire c2571;
    assign in2571_1 = {c73};
    assign in2571_2 = {c74};
    Full_Adder FA_2571(s2571, c2571, in2571_1, in2571_2, c72);
    wire[0:0] s2572, in2572_1, in2572_2;
    wire c2572;
    assign in2572_1 = {c76};
    assign in2572_2 = {c77};
    Full_Adder FA_2572(s2572, c2572, in2572_1, in2572_2, c75);
    wire[0:0] s2573, in2573_1, in2573_2;
    wire c2573;
    assign in2573_1 = {s79[0]};
    assign in2573_2 = {s80[0]};
    Full_Adder FA_2573(s2573, c2573, in2573_1, in2573_2, c78);
    wire[0:0] s2574, in2574_1, in2574_2;
    wire c2574;
    assign in2574_1 = {s82[0]};
    assign in2574_2 = {s83[0]};
    Full_Adder FA_2574(s2574, c2574, in2574_1, in2574_2, s81[0]);
    wire[0:0] s2575, in2575_1, in2575_2;
    wire c2575;
    assign in2575_1 = {s85[0]};
    assign in2575_2 = {s86[0]};
    Full_Adder FA_2575(s2575, c2575, in2575_1, in2575_2, s84[0]);
    wire[0:0] s2576, in2576_1, in2576_2;
    wire c2576;
    assign in2576_1 = {s88[0]};
    assign in2576_2 = {s89[0]};
    Full_Adder FA_2576(s2576, c2576, in2576_1, in2576_2, s87[0]);
    wire[0:0] s2577, in2577_1, in2577_2;
    wire c2577;
    assign in2577_1 = {pp42[57]};
    assign in2577_2 = {pp43[56]};
    Full_Adder FA_2577(s2577, c2577, in2577_1, in2577_2, pp41[58]);
    wire[0:0] s2578, in2578_1, in2578_2;
    wire c2578;
    assign in2578_1 = {pp45[54]};
    assign in2578_2 = {pp46[53]};
    Full_Adder FA_2578(s2578, c2578, in2578_1, in2578_2, pp44[55]);
    wire[0:0] s2579, in2579_1, in2579_2;
    wire c2579;
    assign in2579_1 = {pp48[51]};
    assign in2579_2 = {pp49[50]};
    Full_Adder FA_2579(s2579, c2579, in2579_1, in2579_2, pp47[52]);
    wire[0:0] s2580, in2580_1, in2580_2;
    wire c2580;
    assign in2580_1 = {pp51[48]};
    assign in2580_2 = {pp52[47]};
    Full_Adder FA_2580(s2580, c2580, in2580_1, in2580_2, pp50[49]);
    wire[0:0] s2581, in2581_1, in2581_2;
    wire c2581;
    assign in2581_1 = {pp54[45]};
    assign in2581_2 = {pp55[44]};
    Full_Adder FA_2581(s2581, c2581, in2581_1, in2581_2, pp53[46]);
    wire[0:0] s2582, in2582_1, in2582_2;
    wire c2582;
    assign in2582_1 = {pp57[42]};
    assign in2582_2 = {pp58[41]};
    Full_Adder FA_2582(s2582, c2582, in2582_1, in2582_2, pp56[43]);
    wire[0:0] s2583, in2583_1, in2583_2;
    wire c2583;
    assign in2583_1 = {pp60[39]};
    assign in2583_2 = {pp61[38]};
    Full_Adder FA_2583(s2583, c2583, in2583_1, in2583_2, pp59[40]);
    wire[0:0] s2584, in2584_1, in2584_2;
    wire c2584;
    assign in2584_1 = {pp63[36]};
    assign in2584_2 = {pp64[35]};
    Full_Adder FA_2584(s2584, c2584, in2584_1, in2584_2, pp62[37]);
    wire[0:0] s2585, in2585_1, in2585_2;
    wire c2585;
    assign in2585_1 = {pp66[33]};
    assign in2585_2 = {pp67[32]};
    Full_Adder FA_2585(s2585, c2585, in2585_1, in2585_2, pp65[34]);
    wire[0:0] s2586, in2586_1, in2586_2;
    wire c2586;
    assign in2586_1 = {pp69[30]};
    assign in2586_2 = {pp70[29]};
    Full_Adder FA_2586(s2586, c2586, in2586_1, in2586_2, pp68[31]);
    wire[0:0] s2587, in2587_1, in2587_2;
    wire c2587;
    assign in2587_1 = {pp72[27]};
    assign in2587_2 = {pp73[26]};
    Full_Adder FA_2587(s2587, c2587, in2587_1, in2587_2, pp71[28]);
    wire[0:0] s2588, in2588_1, in2588_2;
    wire c2588;
    assign in2588_1 = {pp75[24]};
    assign in2588_2 = {pp76[23]};
    Full_Adder FA_2588(s2588, c2588, in2588_1, in2588_2, pp74[25]);
    wire[0:0] s2589, in2589_1, in2589_2;
    wire c2589;
    assign in2589_1 = {pp78[21]};
    assign in2589_2 = {pp79[20]};
    Full_Adder FA_2589(s2589, c2589, in2589_1, in2589_2, pp77[22]);
    wire[0:0] s2590, in2590_1, in2590_2;
    wire c2590;
    assign in2590_1 = {pp81[18]};
    assign in2590_2 = {pp82[17]};
    Full_Adder FA_2590(s2590, c2590, in2590_1, in2590_2, pp80[19]);
    wire[0:0] s2591, in2591_1, in2591_2;
    wire c2591;
    assign in2591_1 = {pp84[15]};
    assign in2591_2 = {pp85[14]};
    Full_Adder FA_2591(s2591, c2591, in2591_1, in2591_2, pp83[16]);
    wire[0:0] s2592, in2592_1, in2592_2;
    wire c2592;
    assign in2592_1 = {pp87[12]};
    assign in2592_2 = {pp88[11]};
    Full_Adder FA_2592(s2592, c2592, in2592_1, in2592_2, pp86[13]);
    wire[0:0] s2593, in2593_1, in2593_2;
    wire c2593;
    assign in2593_1 = {pp90[9]};
    assign in2593_2 = {pp91[8]};
    Full_Adder FA_2593(s2593, c2593, in2593_1, in2593_2, pp89[10]);
    wire[0:0] s2594, in2594_1, in2594_2;
    wire c2594;
    assign in2594_1 = {pp93[6]};
    assign in2594_2 = {pp94[5]};
    Full_Adder FA_2594(s2594, c2594, in2594_1, in2594_2, pp92[7]);
    wire[0:0] s2595, in2595_1, in2595_2;
    wire c2595;
    assign in2595_1 = {pp96[3]};
    assign in2595_2 = {pp97[2]};
    Full_Adder FA_2595(s2595, c2595, in2595_1, in2595_2, pp95[4]);
    wire[0:0] s2596, in2596_1, in2596_2;
    wire c2596;
    assign in2596_1 = {pp99[0]};
    assign in2596_2 = {c79};
    Full_Adder FA_2596(s2596, c2596, in2596_1, in2596_2, pp98[1]);
    wire[0:0] s2597, in2597_1, in2597_2;
    wire c2597;
    assign in2597_1 = {c81};
    assign in2597_2 = {c82};
    Full_Adder FA_2597(s2597, c2597, in2597_1, in2597_2, c80);
    wire[0:0] s2598, in2598_1, in2598_2;
    wire c2598;
    assign in2598_1 = {c84};
    assign in2598_2 = {c85};
    Full_Adder FA_2598(s2598, c2598, in2598_1, in2598_2, c83);
    wire[0:0] s2599, in2599_1, in2599_2;
    wire c2599;
    assign in2599_1 = {c87};
    assign in2599_2 = {c88};
    Full_Adder FA_2599(s2599, c2599, in2599_1, in2599_2, c86);
    wire[0:0] s2600, in2600_1, in2600_2;
    wire c2600;
    assign in2600_1 = {c90};
    assign in2600_2 = {c91};
    Full_Adder FA_2600(s2600, c2600, in2600_1, in2600_2, c89);
    wire[0:0] s2601, in2601_1, in2601_2;
    wire c2601;
    assign in2601_1 = {s93[0]};
    assign in2601_2 = {s94[0]};
    Full_Adder FA_2601(s2601, c2601, in2601_1, in2601_2, s92[0]);
    wire[0:0] s2602, in2602_1, in2602_2;
    wire c2602;
    assign in2602_1 = {s96[0]};
    assign in2602_2 = {s97[0]};
    Full_Adder FA_2602(s2602, c2602, in2602_1, in2602_2, s95[0]);
    wire[0:0] s2603, in2603_1, in2603_2;
    wire c2603;
    assign in2603_1 = {s99[0]};
    assign in2603_2 = {s100[0]};
    Full_Adder FA_2603(s2603, c2603, in2603_1, in2603_2, s98[0]);
    wire[0:0] s2604, in2604_1, in2604_2;
    wire c2604;
    assign in2604_1 = {s102[0]};
    assign in2604_2 = {s103[0]};
    Full_Adder FA_2604(s2604, c2604, in2604_1, in2604_2, s101[0]);
    wire[0:0] s2605, in2605_1, in2605_2;
    wire c2605;
    assign in2605_1 = {pp45[55]};
    assign in2605_2 = {pp46[54]};
    Full_Adder FA_2605(s2605, c2605, in2605_1, in2605_2, pp44[56]);
    wire[0:0] s2606, in2606_1, in2606_2;
    wire c2606;
    assign in2606_1 = {pp48[52]};
    assign in2606_2 = {pp49[51]};
    Full_Adder FA_2606(s2606, c2606, in2606_1, in2606_2, pp47[53]);
    wire[0:0] s2607, in2607_1, in2607_2;
    wire c2607;
    assign in2607_1 = {pp51[49]};
    assign in2607_2 = {pp52[48]};
    Full_Adder FA_2607(s2607, c2607, in2607_1, in2607_2, pp50[50]);
    wire[0:0] s2608, in2608_1, in2608_2;
    wire c2608;
    assign in2608_1 = {pp54[46]};
    assign in2608_2 = {pp55[45]};
    Full_Adder FA_2608(s2608, c2608, in2608_1, in2608_2, pp53[47]);
    wire[0:0] s2609, in2609_1, in2609_2;
    wire c2609;
    assign in2609_1 = {pp57[43]};
    assign in2609_2 = {pp58[42]};
    Full_Adder FA_2609(s2609, c2609, in2609_1, in2609_2, pp56[44]);
    wire[0:0] s2610, in2610_1, in2610_2;
    wire c2610;
    assign in2610_1 = {pp60[40]};
    assign in2610_2 = {pp61[39]};
    Full_Adder FA_2610(s2610, c2610, in2610_1, in2610_2, pp59[41]);
    wire[0:0] s2611, in2611_1, in2611_2;
    wire c2611;
    assign in2611_1 = {pp63[37]};
    assign in2611_2 = {pp64[36]};
    Full_Adder FA_2611(s2611, c2611, in2611_1, in2611_2, pp62[38]);
    wire[0:0] s2612, in2612_1, in2612_2;
    wire c2612;
    assign in2612_1 = {pp66[34]};
    assign in2612_2 = {pp67[33]};
    Full_Adder FA_2612(s2612, c2612, in2612_1, in2612_2, pp65[35]);
    wire[0:0] s2613, in2613_1, in2613_2;
    wire c2613;
    assign in2613_1 = {pp69[31]};
    assign in2613_2 = {pp70[30]};
    Full_Adder FA_2613(s2613, c2613, in2613_1, in2613_2, pp68[32]);
    wire[0:0] s2614, in2614_1, in2614_2;
    wire c2614;
    assign in2614_1 = {pp72[28]};
    assign in2614_2 = {pp73[27]};
    Full_Adder FA_2614(s2614, c2614, in2614_1, in2614_2, pp71[29]);
    wire[0:0] s2615, in2615_1, in2615_2;
    wire c2615;
    assign in2615_1 = {pp75[25]};
    assign in2615_2 = {pp76[24]};
    Full_Adder FA_2615(s2615, c2615, in2615_1, in2615_2, pp74[26]);
    wire[0:0] s2616, in2616_1, in2616_2;
    wire c2616;
    assign in2616_1 = {pp78[22]};
    assign in2616_2 = {pp79[21]};
    Full_Adder FA_2616(s2616, c2616, in2616_1, in2616_2, pp77[23]);
    wire[0:0] s2617, in2617_1, in2617_2;
    wire c2617;
    assign in2617_1 = {pp81[19]};
    assign in2617_2 = {pp82[18]};
    Full_Adder FA_2617(s2617, c2617, in2617_1, in2617_2, pp80[20]);
    wire[0:0] s2618, in2618_1, in2618_2;
    wire c2618;
    assign in2618_1 = {pp84[16]};
    assign in2618_2 = {pp85[15]};
    Full_Adder FA_2618(s2618, c2618, in2618_1, in2618_2, pp83[17]);
    wire[0:0] s2619, in2619_1, in2619_2;
    wire c2619;
    assign in2619_1 = {pp87[13]};
    assign in2619_2 = {pp88[12]};
    Full_Adder FA_2619(s2619, c2619, in2619_1, in2619_2, pp86[14]);
    wire[0:0] s2620, in2620_1, in2620_2;
    wire c2620;
    assign in2620_1 = {pp90[10]};
    assign in2620_2 = {pp91[9]};
    Full_Adder FA_2620(s2620, c2620, in2620_1, in2620_2, pp89[11]);
    wire[0:0] s2621, in2621_1, in2621_2;
    wire c2621;
    assign in2621_1 = {pp93[7]};
    assign in2621_2 = {pp94[6]};
    Full_Adder FA_2621(s2621, c2621, in2621_1, in2621_2, pp92[8]);
    wire[0:0] s2622, in2622_1, in2622_2;
    wire c2622;
    assign in2622_1 = {pp96[4]};
    assign in2622_2 = {pp97[3]};
    Full_Adder FA_2622(s2622, c2622, in2622_1, in2622_2, pp95[5]);
    wire[0:0] s2623, in2623_1, in2623_2;
    wire c2623;
    assign in2623_1 = {pp99[1]};
    assign in2623_2 = {pp100[0]};
    Full_Adder FA_2623(s2623, c2623, in2623_1, in2623_2, pp98[2]);
    wire[0:0] s2624, in2624_1, in2624_2;
    wire c2624;
    assign in2624_1 = {c93};
    assign in2624_2 = {c94};
    Full_Adder FA_2624(s2624, c2624, in2624_1, in2624_2, c92);
    wire[0:0] s2625, in2625_1, in2625_2;
    wire c2625;
    assign in2625_1 = {c96};
    assign in2625_2 = {c97};
    Full_Adder FA_2625(s2625, c2625, in2625_1, in2625_2, c95);
    wire[0:0] s2626, in2626_1, in2626_2;
    wire c2626;
    assign in2626_1 = {c99};
    assign in2626_2 = {c100};
    Full_Adder FA_2626(s2626, c2626, in2626_1, in2626_2, c98);
    wire[0:0] s2627, in2627_1, in2627_2;
    wire c2627;
    assign in2627_1 = {c102};
    assign in2627_2 = {c103};
    Full_Adder FA_2627(s2627, c2627, in2627_1, in2627_2, c101);
    wire[0:0] s2628, in2628_1, in2628_2;
    wire c2628;
    assign in2628_1 = {c105};
    assign in2628_2 = {s106[0]};
    Full_Adder FA_2628(s2628, c2628, in2628_1, in2628_2, c104);
    wire[0:0] s2629, in2629_1, in2629_2;
    wire c2629;
    assign in2629_1 = {s108[0]};
    assign in2629_2 = {s109[0]};
    Full_Adder FA_2629(s2629, c2629, in2629_1, in2629_2, s107[0]);
    wire[0:0] s2630, in2630_1, in2630_2;
    wire c2630;
    assign in2630_1 = {s111[0]};
    assign in2630_2 = {s112[0]};
    Full_Adder FA_2630(s2630, c2630, in2630_1, in2630_2, s110[0]);
    wire[0:0] s2631, in2631_1, in2631_2;
    wire c2631;
    assign in2631_1 = {s114[0]};
    assign in2631_2 = {s115[0]};
    Full_Adder FA_2631(s2631, c2631, in2631_1, in2631_2, s113[0]);
    wire[0:0] s2632, in2632_1, in2632_2;
    wire c2632;
    assign in2632_1 = {s117[0]};
    assign in2632_2 = {s118[0]};
    Full_Adder FA_2632(s2632, c2632, in2632_1, in2632_2, s116[0]);
    wire[0:0] s2633, in2633_1, in2633_2;
    wire c2633;
    assign in2633_1 = {pp48[53]};
    assign in2633_2 = {pp49[52]};
    Full_Adder FA_2633(s2633, c2633, in2633_1, in2633_2, pp47[54]);
    wire[0:0] s2634, in2634_1, in2634_2;
    wire c2634;
    assign in2634_1 = {pp51[50]};
    assign in2634_2 = {pp52[49]};
    Full_Adder FA_2634(s2634, c2634, in2634_1, in2634_2, pp50[51]);
    wire[0:0] s2635, in2635_1, in2635_2;
    wire c2635;
    assign in2635_1 = {pp54[47]};
    assign in2635_2 = {pp55[46]};
    Full_Adder FA_2635(s2635, c2635, in2635_1, in2635_2, pp53[48]);
    wire[0:0] s2636, in2636_1, in2636_2;
    wire c2636;
    assign in2636_1 = {pp57[44]};
    assign in2636_2 = {pp58[43]};
    Full_Adder FA_2636(s2636, c2636, in2636_1, in2636_2, pp56[45]);
    wire[0:0] s2637, in2637_1, in2637_2;
    wire c2637;
    assign in2637_1 = {pp60[41]};
    assign in2637_2 = {pp61[40]};
    Full_Adder FA_2637(s2637, c2637, in2637_1, in2637_2, pp59[42]);
    wire[0:0] s2638, in2638_1, in2638_2;
    wire c2638;
    assign in2638_1 = {pp63[38]};
    assign in2638_2 = {pp64[37]};
    Full_Adder FA_2638(s2638, c2638, in2638_1, in2638_2, pp62[39]);
    wire[0:0] s2639, in2639_1, in2639_2;
    wire c2639;
    assign in2639_1 = {pp66[35]};
    assign in2639_2 = {pp67[34]};
    Full_Adder FA_2639(s2639, c2639, in2639_1, in2639_2, pp65[36]);
    wire[0:0] s2640, in2640_1, in2640_2;
    wire c2640;
    assign in2640_1 = {pp69[32]};
    assign in2640_2 = {pp70[31]};
    Full_Adder FA_2640(s2640, c2640, in2640_1, in2640_2, pp68[33]);
    wire[0:0] s2641, in2641_1, in2641_2;
    wire c2641;
    assign in2641_1 = {pp72[29]};
    assign in2641_2 = {pp73[28]};
    Full_Adder FA_2641(s2641, c2641, in2641_1, in2641_2, pp71[30]);
    wire[0:0] s2642, in2642_1, in2642_2;
    wire c2642;
    assign in2642_1 = {pp75[26]};
    assign in2642_2 = {pp76[25]};
    Full_Adder FA_2642(s2642, c2642, in2642_1, in2642_2, pp74[27]);
    wire[0:0] s2643, in2643_1, in2643_2;
    wire c2643;
    assign in2643_1 = {pp78[23]};
    assign in2643_2 = {pp79[22]};
    Full_Adder FA_2643(s2643, c2643, in2643_1, in2643_2, pp77[24]);
    wire[0:0] s2644, in2644_1, in2644_2;
    wire c2644;
    assign in2644_1 = {pp81[20]};
    assign in2644_2 = {pp82[19]};
    Full_Adder FA_2644(s2644, c2644, in2644_1, in2644_2, pp80[21]);
    wire[0:0] s2645, in2645_1, in2645_2;
    wire c2645;
    assign in2645_1 = {pp84[17]};
    assign in2645_2 = {pp85[16]};
    Full_Adder FA_2645(s2645, c2645, in2645_1, in2645_2, pp83[18]);
    wire[0:0] s2646, in2646_1, in2646_2;
    wire c2646;
    assign in2646_1 = {pp87[14]};
    assign in2646_2 = {pp88[13]};
    Full_Adder FA_2646(s2646, c2646, in2646_1, in2646_2, pp86[15]);
    wire[0:0] s2647, in2647_1, in2647_2;
    wire c2647;
    assign in2647_1 = {pp90[11]};
    assign in2647_2 = {pp91[10]};
    Full_Adder FA_2647(s2647, c2647, in2647_1, in2647_2, pp89[12]);
    wire[0:0] s2648, in2648_1, in2648_2;
    wire c2648;
    assign in2648_1 = {pp93[8]};
    assign in2648_2 = {pp94[7]};
    Full_Adder FA_2648(s2648, c2648, in2648_1, in2648_2, pp92[9]);
    wire[0:0] s2649, in2649_1, in2649_2;
    wire c2649;
    assign in2649_1 = {pp96[5]};
    assign in2649_2 = {pp97[4]};
    Full_Adder FA_2649(s2649, c2649, in2649_1, in2649_2, pp95[6]);
    wire[0:0] s2650, in2650_1, in2650_2;
    wire c2650;
    assign in2650_1 = {pp99[2]};
    assign in2650_2 = {pp100[1]};
    Full_Adder FA_2650(s2650, c2650, in2650_1, in2650_2, pp98[3]);
    wire[0:0] s2651, in2651_1, in2651_2;
    wire c2651;
    assign in2651_1 = {c106};
    assign in2651_2 = {c107};
    Full_Adder FA_2651(s2651, c2651, in2651_1, in2651_2, pp101[0]);
    wire[0:0] s2652, in2652_1, in2652_2;
    wire c2652;
    assign in2652_1 = {c109};
    assign in2652_2 = {c110};
    Full_Adder FA_2652(s2652, c2652, in2652_1, in2652_2, c108);
    wire[0:0] s2653, in2653_1, in2653_2;
    wire c2653;
    assign in2653_1 = {c112};
    assign in2653_2 = {c113};
    Full_Adder FA_2653(s2653, c2653, in2653_1, in2653_2, c111);
    wire[0:0] s2654, in2654_1, in2654_2;
    wire c2654;
    assign in2654_1 = {c115};
    assign in2654_2 = {c116};
    Full_Adder FA_2654(s2654, c2654, in2654_1, in2654_2, c114);
    wire[0:0] s2655, in2655_1, in2655_2;
    wire c2655;
    assign in2655_1 = {c118};
    assign in2655_2 = {c119};
    Full_Adder FA_2655(s2655, c2655, in2655_1, in2655_2, c117);
    wire[0:0] s2656, in2656_1, in2656_2;
    wire c2656;
    assign in2656_1 = {s121[0]};
    assign in2656_2 = {s122[0]};
    Full_Adder FA_2656(s2656, c2656, in2656_1, in2656_2, c120);
    wire[0:0] s2657, in2657_1, in2657_2;
    wire c2657;
    assign in2657_1 = {s124[0]};
    assign in2657_2 = {s125[0]};
    Full_Adder FA_2657(s2657, c2657, in2657_1, in2657_2, s123[0]);
    wire[0:0] s2658, in2658_1, in2658_2;
    wire c2658;
    assign in2658_1 = {s127[0]};
    assign in2658_2 = {s128[0]};
    Full_Adder FA_2658(s2658, c2658, in2658_1, in2658_2, s126[0]);
    wire[0:0] s2659, in2659_1, in2659_2;
    wire c2659;
    assign in2659_1 = {s130[0]};
    assign in2659_2 = {s131[0]};
    Full_Adder FA_2659(s2659, c2659, in2659_1, in2659_2, s129[0]);
    wire[0:0] s2660, in2660_1, in2660_2;
    wire c2660;
    assign in2660_1 = {s133[0]};
    assign in2660_2 = {s134[0]};
    Full_Adder FA_2660(s2660, c2660, in2660_1, in2660_2, s132[0]);
    wire[0:0] s2661, in2661_1, in2661_2;
    wire c2661;
    assign in2661_1 = {pp51[51]};
    assign in2661_2 = {pp52[50]};
    Full_Adder FA_2661(s2661, c2661, in2661_1, in2661_2, pp50[52]);
    wire[0:0] s2662, in2662_1, in2662_2;
    wire c2662;
    assign in2662_1 = {pp54[48]};
    assign in2662_2 = {pp55[47]};
    Full_Adder FA_2662(s2662, c2662, in2662_1, in2662_2, pp53[49]);
    wire[0:0] s2663, in2663_1, in2663_2;
    wire c2663;
    assign in2663_1 = {pp57[45]};
    assign in2663_2 = {pp58[44]};
    Full_Adder FA_2663(s2663, c2663, in2663_1, in2663_2, pp56[46]);
    wire[0:0] s2664, in2664_1, in2664_2;
    wire c2664;
    assign in2664_1 = {pp60[42]};
    assign in2664_2 = {pp61[41]};
    Full_Adder FA_2664(s2664, c2664, in2664_1, in2664_2, pp59[43]);
    wire[0:0] s2665, in2665_1, in2665_2;
    wire c2665;
    assign in2665_1 = {pp63[39]};
    assign in2665_2 = {pp64[38]};
    Full_Adder FA_2665(s2665, c2665, in2665_1, in2665_2, pp62[40]);
    wire[0:0] s2666, in2666_1, in2666_2;
    wire c2666;
    assign in2666_1 = {pp66[36]};
    assign in2666_2 = {pp67[35]};
    Full_Adder FA_2666(s2666, c2666, in2666_1, in2666_2, pp65[37]);
    wire[0:0] s2667, in2667_1, in2667_2;
    wire c2667;
    assign in2667_1 = {pp69[33]};
    assign in2667_2 = {pp70[32]};
    Full_Adder FA_2667(s2667, c2667, in2667_1, in2667_2, pp68[34]);
    wire[0:0] s2668, in2668_1, in2668_2;
    wire c2668;
    assign in2668_1 = {pp72[30]};
    assign in2668_2 = {pp73[29]};
    Full_Adder FA_2668(s2668, c2668, in2668_1, in2668_2, pp71[31]);
    wire[0:0] s2669, in2669_1, in2669_2;
    wire c2669;
    assign in2669_1 = {pp75[27]};
    assign in2669_2 = {pp76[26]};
    Full_Adder FA_2669(s2669, c2669, in2669_1, in2669_2, pp74[28]);
    wire[0:0] s2670, in2670_1, in2670_2;
    wire c2670;
    assign in2670_1 = {pp78[24]};
    assign in2670_2 = {pp79[23]};
    Full_Adder FA_2670(s2670, c2670, in2670_1, in2670_2, pp77[25]);
    wire[0:0] s2671, in2671_1, in2671_2;
    wire c2671;
    assign in2671_1 = {pp81[21]};
    assign in2671_2 = {pp82[20]};
    Full_Adder FA_2671(s2671, c2671, in2671_1, in2671_2, pp80[22]);
    wire[0:0] s2672, in2672_1, in2672_2;
    wire c2672;
    assign in2672_1 = {pp84[18]};
    assign in2672_2 = {pp85[17]};
    Full_Adder FA_2672(s2672, c2672, in2672_1, in2672_2, pp83[19]);
    wire[0:0] s2673, in2673_1, in2673_2;
    wire c2673;
    assign in2673_1 = {pp87[15]};
    assign in2673_2 = {pp88[14]};
    Full_Adder FA_2673(s2673, c2673, in2673_1, in2673_2, pp86[16]);
    wire[0:0] s2674, in2674_1, in2674_2;
    wire c2674;
    assign in2674_1 = {pp90[12]};
    assign in2674_2 = {pp91[11]};
    Full_Adder FA_2674(s2674, c2674, in2674_1, in2674_2, pp89[13]);
    wire[0:0] s2675, in2675_1, in2675_2;
    wire c2675;
    assign in2675_1 = {pp93[9]};
    assign in2675_2 = {pp94[8]};
    Full_Adder FA_2675(s2675, c2675, in2675_1, in2675_2, pp92[10]);
    wire[0:0] s2676, in2676_1, in2676_2;
    wire c2676;
    assign in2676_1 = {pp96[6]};
    assign in2676_2 = {pp97[5]};
    Full_Adder FA_2676(s2676, c2676, in2676_1, in2676_2, pp95[7]);
    wire[0:0] s2677, in2677_1, in2677_2;
    wire c2677;
    assign in2677_1 = {pp99[3]};
    assign in2677_2 = {pp100[2]};
    Full_Adder FA_2677(s2677, c2677, in2677_1, in2677_2, pp98[4]);
    wire[0:0] s2678, in2678_1, in2678_2;
    wire c2678;
    assign in2678_1 = {pp102[0]};
    assign in2678_2 = {c121};
    Full_Adder FA_2678(s2678, c2678, in2678_1, in2678_2, pp101[1]);
    wire[0:0] s2679, in2679_1, in2679_2;
    wire c2679;
    assign in2679_1 = {c123};
    assign in2679_2 = {c124};
    Full_Adder FA_2679(s2679, c2679, in2679_1, in2679_2, c122);
    wire[0:0] s2680, in2680_1, in2680_2;
    wire c2680;
    assign in2680_1 = {c126};
    assign in2680_2 = {c127};
    Full_Adder FA_2680(s2680, c2680, in2680_1, in2680_2, c125);
    wire[0:0] s2681, in2681_1, in2681_2;
    wire c2681;
    assign in2681_1 = {c129};
    assign in2681_2 = {c130};
    Full_Adder FA_2681(s2681, c2681, in2681_1, in2681_2, c128);
    wire[0:0] s2682, in2682_1, in2682_2;
    wire c2682;
    assign in2682_1 = {c132};
    assign in2682_2 = {c133};
    Full_Adder FA_2682(s2682, c2682, in2682_1, in2682_2, c131);
    wire[0:0] s2683, in2683_1, in2683_2;
    wire c2683;
    assign in2683_1 = {c135};
    assign in2683_2 = {c136};
    Full_Adder FA_2683(s2683, c2683, in2683_1, in2683_2, c134);
    wire[0:0] s2684, in2684_1, in2684_2;
    wire c2684;
    assign in2684_1 = {s138[0]};
    assign in2684_2 = {s139[0]};
    Full_Adder FA_2684(s2684, c2684, in2684_1, in2684_2, s137[0]);
    wire[0:0] s2685, in2685_1, in2685_2;
    wire c2685;
    assign in2685_1 = {s141[0]};
    assign in2685_2 = {s142[0]};
    Full_Adder FA_2685(s2685, c2685, in2685_1, in2685_2, s140[0]);
    wire[0:0] s2686, in2686_1, in2686_2;
    wire c2686;
    assign in2686_1 = {s144[0]};
    assign in2686_2 = {s145[0]};
    Full_Adder FA_2686(s2686, c2686, in2686_1, in2686_2, s143[0]);
    wire[0:0] s2687, in2687_1, in2687_2;
    wire c2687;
    assign in2687_1 = {s147[0]};
    assign in2687_2 = {s148[0]};
    Full_Adder FA_2687(s2687, c2687, in2687_1, in2687_2, s146[0]);
    wire[0:0] s2688, in2688_1, in2688_2;
    wire c2688;
    assign in2688_1 = {s150[0]};
    assign in2688_2 = {s151[0]};
    Full_Adder FA_2688(s2688, c2688, in2688_1, in2688_2, s149[0]);
    wire[0:0] s2689, in2689_1, in2689_2;
    wire c2689;
    assign in2689_1 = {pp54[49]};
    assign in2689_2 = {pp55[48]};
    Full_Adder FA_2689(s2689, c2689, in2689_1, in2689_2, pp53[50]);
    wire[0:0] s2690, in2690_1, in2690_2;
    wire c2690;
    assign in2690_1 = {pp57[46]};
    assign in2690_2 = {pp58[45]};
    Full_Adder FA_2690(s2690, c2690, in2690_1, in2690_2, pp56[47]);
    wire[0:0] s2691, in2691_1, in2691_2;
    wire c2691;
    assign in2691_1 = {pp60[43]};
    assign in2691_2 = {pp61[42]};
    Full_Adder FA_2691(s2691, c2691, in2691_1, in2691_2, pp59[44]);
    wire[0:0] s2692, in2692_1, in2692_2;
    wire c2692;
    assign in2692_1 = {pp63[40]};
    assign in2692_2 = {pp64[39]};
    Full_Adder FA_2692(s2692, c2692, in2692_1, in2692_2, pp62[41]);
    wire[0:0] s2693, in2693_1, in2693_2;
    wire c2693;
    assign in2693_1 = {pp66[37]};
    assign in2693_2 = {pp67[36]};
    Full_Adder FA_2693(s2693, c2693, in2693_1, in2693_2, pp65[38]);
    wire[0:0] s2694, in2694_1, in2694_2;
    wire c2694;
    assign in2694_1 = {pp69[34]};
    assign in2694_2 = {pp70[33]};
    Full_Adder FA_2694(s2694, c2694, in2694_1, in2694_2, pp68[35]);
    wire[0:0] s2695, in2695_1, in2695_2;
    wire c2695;
    assign in2695_1 = {pp72[31]};
    assign in2695_2 = {pp73[30]};
    Full_Adder FA_2695(s2695, c2695, in2695_1, in2695_2, pp71[32]);
    wire[0:0] s2696, in2696_1, in2696_2;
    wire c2696;
    assign in2696_1 = {pp75[28]};
    assign in2696_2 = {pp76[27]};
    Full_Adder FA_2696(s2696, c2696, in2696_1, in2696_2, pp74[29]);
    wire[0:0] s2697, in2697_1, in2697_2;
    wire c2697;
    assign in2697_1 = {pp78[25]};
    assign in2697_2 = {pp79[24]};
    Full_Adder FA_2697(s2697, c2697, in2697_1, in2697_2, pp77[26]);
    wire[0:0] s2698, in2698_1, in2698_2;
    wire c2698;
    assign in2698_1 = {pp81[22]};
    assign in2698_2 = {pp82[21]};
    Full_Adder FA_2698(s2698, c2698, in2698_1, in2698_2, pp80[23]);
    wire[0:0] s2699, in2699_1, in2699_2;
    wire c2699;
    assign in2699_1 = {pp84[19]};
    assign in2699_2 = {pp85[18]};
    Full_Adder FA_2699(s2699, c2699, in2699_1, in2699_2, pp83[20]);
    wire[0:0] s2700, in2700_1, in2700_2;
    wire c2700;
    assign in2700_1 = {pp87[16]};
    assign in2700_2 = {pp88[15]};
    Full_Adder FA_2700(s2700, c2700, in2700_1, in2700_2, pp86[17]);
    wire[0:0] s2701, in2701_1, in2701_2;
    wire c2701;
    assign in2701_1 = {pp90[13]};
    assign in2701_2 = {pp91[12]};
    Full_Adder FA_2701(s2701, c2701, in2701_1, in2701_2, pp89[14]);
    wire[0:0] s2702, in2702_1, in2702_2;
    wire c2702;
    assign in2702_1 = {pp93[10]};
    assign in2702_2 = {pp94[9]};
    Full_Adder FA_2702(s2702, c2702, in2702_1, in2702_2, pp92[11]);
    wire[0:0] s2703, in2703_1, in2703_2;
    wire c2703;
    assign in2703_1 = {pp96[7]};
    assign in2703_2 = {pp97[6]};
    Full_Adder FA_2703(s2703, c2703, in2703_1, in2703_2, pp95[8]);
    wire[0:0] s2704, in2704_1, in2704_2;
    wire c2704;
    assign in2704_1 = {pp99[4]};
    assign in2704_2 = {pp100[3]};
    Full_Adder FA_2704(s2704, c2704, in2704_1, in2704_2, pp98[5]);
    wire[0:0] s2705, in2705_1, in2705_2;
    wire c2705;
    assign in2705_1 = {pp102[1]};
    assign in2705_2 = {pp103[0]};
    Full_Adder FA_2705(s2705, c2705, in2705_1, in2705_2, pp101[2]);
    wire[0:0] s2706, in2706_1, in2706_2;
    wire c2706;
    assign in2706_1 = {c138};
    assign in2706_2 = {c139};
    Full_Adder FA_2706(s2706, c2706, in2706_1, in2706_2, c137);
    wire[0:0] s2707, in2707_1, in2707_2;
    wire c2707;
    assign in2707_1 = {c141};
    assign in2707_2 = {c142};
    Full_Adder FA_2707(s2707, c2707, in2707_1, in2707_2, c140);
    wire[0:0] s2708, in2708_1, in2708_2;
    wire c2708;
    assign in2708_1 = {c144};
    assign in2708_2 = {c145};
    Full_Adder FA_2708(s2708, c2708, in2708_1, in2708_2, c143);
    wire[0:0] s2709, in2709_1, in2709_2;
    wire c2709;
    assign in2709_1 = {c147};
    assign in2709_2 = {c148};
    Full_Adder FA_2709(s2709, c2709, in2709_1, in2709_2, c146);
    wire[0:0] s2710, in2710_1, in2710_2;
    wire c2710;
    assign in2710_1 = {c150};
    assign in2710_2 = {c151};
    Full_Adder FA_2710(s2710, c2710, in2710_1, in2710_2, c149);
    wire[0:0] s2711, in2711_1, in2711_2;
    wire c2711;
    assign in2711_1 = {c153};
    assign in2711_2 = {s154[0]};
    Full_Adder FA_2711(s2711, c2711, in2711_1, in2711_2, c152);
    wire[0:0] s2712, in2712_1, in2712_2;
    wire c2712;
    assign in2712_1 = {s156[0]};
    assign in2712_2 = {s157[0]};
    Full_Adder FA_2712(s2712, c2712, in2712_1, in2712_2, s155[0]);
    wire[0:0] s2713, in2713_1, in2713_2;
    wire c2713;
    assign in2713_1 = {s159[0]};
    assign in2713_2 = {s160[0]};
    Full_Adder FA_2713(s2713, c2713, in2713_1, in2713_2, s158[0]);
    wire[0:0] s2714, in2714_1, in2714_2;
    wire c2714;
    assign in2714_1 = {s162[0]};
    assign in2714_2 = {s163[0]};
    Full_Adder FA_2714(s2714, c2714, in2714_1, in2714_2, s161[0]);
    wire[0:0] s2715, in2715_1, in2715_2;
    wire c2715;
    assign in2715_1 = {s165[0]};
    assign in2715_2 = {s166[0]};
    Full_Adder FA_2715(s2715, c2715, in2715_1, in2715_2, s164[0]);
    wire[0:0] s2716, in2716_1, in2716_2;
    wire c2716;
    assign in2716_1 = {s168[0]};
    assign in2716_2 = {s169[0]};
    Full_Adder FA_2716(s2716, c2716, in2716_1, in2716_2, s167[0]);
    wire[0:0] s2717, in2717_1, in2717_2;
    wire c2717;
    assign in2717_1 = {pp57[47]};
    assign in2717_2 = {pp58[46]};
    Full_Adder FA_2717(s2717, c2717, in2717_1, in2717_2, pp56[48]);
    wire[0:0] s2718, in2718_1, in2718_2;
    wire c2718;
    assign in2718_1 = {pp60[44]};
    assign in2718_2 = {pp61[43]};
    Full_Adder FA_2718(s2718, c2718, in2718_1, in2718_2, pp59[45]);
    wire[0:0] s2719, in2719_1, in2719_2;
    wire c2719;
    assign in2719_1 = {pp63[41]};
    assign in2719_2 = {pp64[40]};
    Full_Adder FA_2719(s2719, c2719, in2719_1, in2719_2, pp62[42]);
    wire[0:0] s2720, in2720_1, in2720_2;
    wire c2720;
    assign in2720_1 = {pp66[38]};
    assign in2720_2 = {pp67[37]};
    Full_Adder FA_2720(s2720, c2720, in2720_1, in2720_2, pp65[39]);
    wire[0:0] s2721, in2721_1, in2721_2;
    wire c2721;
    assign in2721_1 = {pp69[35]};
    assign in2721_2 = {pp70[34]};
    Full_Adder FA_2721(s2721, c2721, in2721_1, in2721_2, pp68[36]);
    wire[0:0] s2722, in2722_1, in2722_2;
    wire c2722;
    assign in2722_1 = {pp72[32]};
    assign in2722_2 = {pp73[31]};
    Full_Adder FA_2722(s2722, c2722, in2722_1, in2722_2, pp71[33]);
    wire[0:0] s2723, in2723_1, in2723_2;
    wire c2723;
    assign in2723_1 = {pp75[29]};
    assign in2723_2 = {pp76[28]};
    Full_Adder FA_2723(s2723, c2723, in2723_1, in2723_2, pp74[30]);
    wire[0:0] s2724, in2724_1, in2724_2;
    wire c2724;
    assign in2724_1 = {pp78[26]};
    assign in2724_2 = {pp79[25]};
    Full_Adder FA_2724(s2724, c2724, in2724_1, in2724_2, pp77[27]);
    wire[0:0] s2725, in2725_1, in2725_2;
    wire c2725;
    assign in2725_1 = {pp81[23]};
    assign in2725_2 = {pp82[22]};
    Full_Adder FA_2725(s2725, c2725, in2725_1, in2725_2, pp80[24]);
    wire[0:0] s2726, in2726_1, in2726_2;
    wire c2726;
    assign in2726_1 = {pp84[20]};
    assign in2726_2 = {pp85[19]};
    Full_Adder FA_2726(s2726, c2726, in2726_1, in2726_2, pp83[21]);
    wire[0:0] s2727, in2727_1, in2727_2;
    wire c2727;
    assign in2727_1 = {pp87[17]};
    assign in2727_2 = {pp88[16]};
    Full_Adder FA_2727(s2727, c2727, in2727_1, in2727_2, pp86[18]);
    wire[0:0] s2728, in2728_1, in2728_2;
    wire c2728;
    assign in2728_1 = {pp90[14]};
    assign in2728_2 = {pp91[13]};
    Full_Adder FA_2728(s2728, c2728, in2728_1, in2728_2, pp89[15]);
    wire[0:0] s2729, in2729_1, in2729_2;
    wire c2729;
    assign in2729_1 = {pp93[11]};
    assign in2729_2 = {pp94[10]};
    Full_Adder FA_2729(s2729, c2729, in2729_1, in2729_2, pp92[12]);
    wire[0:0] s2730, in2730_1, in2730_2;
    wire c2730;
    assign in2730_1 = {pp96[8]};
    assign in2730_2 = {pp97[7]};
    Full_Adder FA_2730(s2730, c2730, in2730_1, in2730_2, pp95[9]);
    wire[0:0] s2731, in2731_1, in2731_2;
    wire c2731;
    assign in2731_1 = {pp99[5]};
    assign in2731_2 = {pp100[4]};
    Full_Adder FA_2731(s2731, c2731, in2731_1, in2731_2, pp98[6]);
    wire[0:0] s2732, in2732_1, in2732_2;
    wire c2732;
    assign in2732_1 = {pp102[2]};
    assign in2732_2 = {pp103[1]};
    Full_Adder FA_2732(s2732, c2732, in2732_1, in2732_2, pp101[3]);
    wire[0:0] s2733, in2733_1, in2733_2;
    wire c2733;
    assign in2733_1 = {c154};
    assign in2733_2 = {c155};
    Full_Adder FA_2733(s2733, c2733, in2733_1, in2733_2, pp104[0]);
    wire[0:0] s2734, in2734_1, in2734_2;
    wire c2734;
    assign in2734_1 = {c157};
    assign in2734_2 = {c158};
    Full_Adder FA_2734(s2734, c2734, in2734_1, in2734_2, c156);
    wire[0:0] s2735, in2735_1, in2735_2;
    wire c2735;
    assign in2735_1 = {c160};
    assign in2735_2 = {c161};
    Full_Adder FA_2735(s2735, c2735, in2735_1, in2735_2, c159);
    wire[0:0] s2736, in2736_1, in2736_2;
    wire c2736;
    assign in2736_1 = {c163};
    assign in2736_2 = {c164};
    Full_Adder FA_2736(s2736, c2736, in2736_1, in2736_2, c162);
    wire[0:0] s2737, in2737_1, in2737_2;
    wire c2737;
    assign in2737_1 = {c166};
    assign in2737_2 = {c167};
    Full_Adder FA_2737(s2737, c2737, in2737_1, in2737_2, c165);
    wire[0:0] s2738, in2738_1, in2738_2;
    wire c2738;
    assign in2738_1 = {c169};
    assign in2738_2 = {c170};
    Full_Adder FA_2738(s2738, c2738, in2738_1, in2738_2, c168);
    wire[0:0] s2739, in2739_1, in2739_2;
    wire c2739;
    assign in2739_1 = {s172[0]};
    assign in2739_2 = {s173[0]};
    Full_Adder FA_2739(s2739, c2739, in2739_1, in2739_2, c171);
    wire[0:0] s2740, in2740_1, in2740_2;
    wire c2740;
    assign in2740_1 = {s175[0]};
    assign in2740_2 = {s176[0]};
    Full_Adder FA_2740(s2740, c2740, in2740_1, in2740_2, s174[0]);
    wire[0:0] s2741, in2741_1, in2741_2;
    wire c2741;
    assign in2741_1 = {s178[0]};
    assign in2741_2 = {s179[0]};
    Full_Adder FA_2741(s2741, c2741, in2741_1, in2741_2, s177[0]);
    wire[0:0] s2742, in2742_1, in2742_2;
    wire c2742;
    assign in2742_1 = {s181[0]};
    assign in2742_2 = {s182[0]};
    Full_Adder FA_2742(s2742, c2742, in2742_1, in2742_2, s180[0]);
    wire[0:0] s2743, in2743_1, in2743_2;
    wire c2743;
    assign in2743_1 = {s184[0]};
    assign in2743_2 = {s185[0]};
    Full_Adder FA_2743(s2743, c2743, in2743_1, in2743_2, s183[0]);
    wire[0:0] s2744, in2744_1, in2744_2;
    wire c2744;
    assign in2744_1 = {s187[0]};
    assign in2744_2 = {s188[0]};
    Full_Adder FA_2744(s2744, c2744, in2744_1, in2744_2, s186[0]);
    wire[0:0] s2745, in2745_1, in2745_2;
    wire c2745;
    assign in2745_1 = {pp60[45]};
    assign in2745_2 = {pp61[44]};
    Full_Adder FA_2745(s2745, c2745, in2745_1, in2745_2, pp59[46]);
    wire[0:0] s2746, in2746_1, in2746_2;
    wire c2746;
    assign in2746_1 = {pp63[42]};
    assign in2746_2 = {pp64[41]};
    Full_Adder FA_2746(s2746, c2746, in2746_1, in2746_2, pp62[43]);
    wire[0:0] s2747, in2747_1, in2747_2;
    wire c2747;
    assign in2747_1 = {pp66[39]};
    assign in2747_2 = {pp67[38]};
    Full_Adder FA_2747(s2747, c2747, in2747_1, in2747_2, pp65[40]);
    wire[0:0] s2748, in2748_1, in2748_2;
    wire c2748;
    assign in2748_1 = {pp69[36]};
    assign in2748_2 = {pp70[35]};
    Full_Adder FA_2748(s2748, c2748, in2748_1, in2748_2, pp68[37]);
    wire[0:0] s2749, in2749_1, in2749_2;
    wire c2749;
    assign in2749_1 = {pp72[33]};
    assign in2749_2 = {pp73[32]};
    Full_Adder FA_2749(s2749, c2749, in2749_1, in2749_2, pp71[34]);
    wire[0:0] s2750, in2750_1, in2750_2;
    wire c2750;
    assign in2750_1 = {pp75[30]};
    assign in2750_2 = {pp76[29]};
    Full_Adder FA_2750(s2750, c2750, in2750_1, in2750_2, pp74[31]);
    wire[0:0] s2751, in2751_1, in2751_2;
    wire c2751;
    assign in2751_1 = {pp78[27]};
    assign in2751_2 = {pp79[26]};
    Full_Adder FA_2751(s2751, c2751, in2751_1, in2751_2, pp77[28]);
    wire[0:0] s2752, in2752_1, in2752_2;
    wire c2752;
    assign in2752_1 = {pp81[24]};
    assign in2752_2 = {pp82[23]};
    Full_Adder FA_2752(s2752, c2752, in2752_1, in2752_2, pp80[25]);
    wire[0:0] s2753, in2753_1, in2753_2;
    wire c2753;
    assign in2753_1 = {pp84[21]};
    assign in2753_2 = {pp85[20]};
    Full_Adder FA_2753(s2753, c2753, in2753_1, in2753_2, pp83[22]);
    wire[0:0] s2754, in2754_1, in2754_2;
    wire c2754;
    assign in2754_1 = {pp87[18]};
    assign in2754_2 = {pp88[17]};
    Full_Adder FA_2754(s2754, c2754, in2754_1, in2754_2, pp86[19]);
    wire[0:0] s2755, in2755_1, in2755_2;
    wire c2755;
    assign in2755_1 = {pp90[15]};
    assign in2755_2 = {pp91[14]};
    Full_Adder FA_2755(s2755, c2755, in2755_1, in2755_2, pp89[16]);
    wire[0:0] s2756, in2756_1, in2756_2;
    wire c2756;
    assign in2756_1 = {pp93[12]};
    assign in2756_2 = {pp94[11]};
    Full_Adder FA_2756(s2756, c2756, in2756_1, in2756_2, pp92[13]);
    wire[0:0] s2757, in2757_1, in2757_2;
    wire c2757;
    assign in2757_1 = {pp96[9]};
    assign in2757_2 = {pp97[8]};
    Full_Adder FA_2757(s2757, c2757, in2757_1, in2757_2, pp95[10]);
    wire[0:0] s2758, in2758_1, in2758_2;
    wire c2758;
    assign in2758_1 = {pp99[6]};
    assign in2758_2 = {pp100[5]};
    Full_Adder FA_2758(s2758, c2758, in2758_1, in2758_2, pp98[7]);
    wire[0:0] s2759, in2759_1, in2759_2;
    wire c2759;
    assign in2759_1 = {pp102[3]};
    assign in2759_2 = {pp103[2]};
    Full_Adder FA_2759(s2759, c2759, in2759_1, in2759_2, pp101[4]);
    wire[0:0] s2760, in2760_1, in2760_2;
    wire c2760;
    assign in2760_1 = {pp105[0]};
    assign in2760_2 = {c172};
    Full_Adder FA_2760(s2760, c2760, in2760_1, in2760_2, pp104[1]);
    wire[0:0] s2761, in2761_1, in2761_2;
    wire c2761;
    assign in2761_1 = {c174};
    assign in2761_2 = {c175};
    Full_Adder FA_2761(s2761, c2761, in2761_1, in2761_2, c173);
    wire[0:0] s2762, in2762_1, in2762_2;
    wire c2762;
    assign in2762_1 = {c177};
    assign in2762_2 = {c178};
    Full_Adder FA_2762(s2762, c2762, in2762_1, in2762_2, c176);
    wire[0:0] s2763, in2763_1, in2763_2;
    wire c2763;
    assign in2763_1 = {c180};
    assign in2763_2 = {c181};
    Full_Adder FA_2763(s2763, c2763, in2763_1, in2763_2, c179);
    wire[0:0] s2764, in2764_1, in2764_2;
    wire c2764;
    assign in2764_1 = {c183};
    assign in2764_2 = {c184};
    Full_Adder FA_2764(s2764, c2764, in2764_1, in2764_2, c182);
    wire[0:0] s2765, in2765_1, in2765_2;
    wire c2765;
    assign in2765_1 = {c186};
    assign in2765_2 = {c187};
    Full_Adder FA_2765(s2765, c2765, in2765_1, in2765_2, c185);
    wire[0:0] s2766, in2766_1, in2766_2;
    wire c2766;
    assign in2766_1 = {c189};
    assign in2766_2 = {c190};
    Full_Adder FA_2766(s2766, c2766, in2766_1, in2766_2, c188);
    wire[0:0] s2767, in2767_1, in2767_2;
    wire c2767;
    assign in2767_1 = {s192[0]};
    assign in2767_2 = {s193[0]};
    Full_Adder FA_2767(s2767, c2767, in2767_1, in2767_2, s191[0]);
    wire[0:0] s2768, in2768_1, in2768_2;
    wire c2768;
    assign in2768_1 = {s195[0]};
    assign in2768_2 = {s196[0]};
    Full_Adder FA_2768(s2768, c2768, in2768_1, in2768_2, s194[0]);
    wire[0:0] s2769, in2769_1, in2769_2;
    wire c2769;
    assign in2769_1 = {s198[0]};
    assign in2769_2 = {s199[0]};
    Full_Adder FA_2769(s2769, c2769, in2769_1, in2769_2, s197[0]);
    wire[0:0] s2770, in2770_1, in2770_2;
    wire c2770;
    assign in2770_1 = {s201[0]};
    assign in2770_2 = {s202[0]};
    Full_Adder FA_2770(s2770, c2770, in2770_1, in2770_2, s200[0]);
    wire[0:0] s2771, in2771_1, in2771_2;
    wire c2771;
    assign in2771_1 = {s204[0]};
    assign in2771_2 = {s205[0]};
    Full_Adder FA_2771(s2771, c2771, in2771_1, in2771_2, s203[0]);
    wire[0:0] s2772, in2772_1, in2772_2;
    wire c2772;
    assign in2772_1 = {s207[0]};
    assign in2772_2 = {s208[0]};
    Full_Adder FA_2772(s2772, c2772, in2772_1, in2772_2, s206[0]);
    wire[0:0] s2773, in2773_1, in2773_2;
    wire c2773;
    assign in2773_1 = {pp63[43]};
    assign in2773_2 = {pp64[42]};
    Full_Adder FA_2773(s2773, c2773, in2773_1, in2773_2, pp62[44]);
    wire[0:0] s2774, in2774_1, in2774_2;
    wire c2774;
    assign in2774_1 = {pp66[40]};
    assign in2774_2 = {pp67[39]};
    Full_Adder FA_2774(s2774, c2774, in2774_1, in2774_2, pp65[41]);
    wire[0:0] s2775, in2775_1, in2775_2;
    wire c2775;
    assign in2775_1 = {pp69[37]};
    assign in2775_2 = {pp70[36]};
    Full_Adder FA_2775(s2775, c2775, in2775_1, in2775_2, pp68[38]);
    wire[0:0] s2776, in2776_1, in2776_2;
    wire c2776;
    assign in2776_1 = {pp72[34]};
    assign in2776_2 = {pp73[33]};
    Full_Adder FA_2776(s2776, c2776, in2776_1, in2776_2, pp71[35]);
    wire[0:0] s2777, in2777_1, in2777_2;
    wire c2777;
    assign in2777_1 = {pp75[31]};
    assign in2777_2 = {pp76[30]};
    Full_Adder FA_2777(s2777, c2777, in2777_1, in2777_2, pp74[32]);
    wire[0:0] s2778, in2778_1, in2778_2;
    wire c2778;
    assign in2778_1 = {pp78[28]};
    assign in2778_2 = {pp79[27]};
    Full_Adder FA_2778(s2778, c2778, in2778_1, in2778_2, pp77[29]);
    wire[0:0] s2779, in2779_1, in2779_2;
    wire c2779;
    assign in2779_1 = {pp81[25]};
    assign in2779_2 = {pp82[24]};
    Full_Adder FA_2779(s2779, c2779, in2779_1, in2779_2, pp80[26]);
    wire[0:0] s2780, in2780_1, in2780_2;
    wire c2780;
    assign in2780_1 = {pp84[22]};
    assign in2780_2 = {pp85[21]};
    Full_Adder FA_2780(s2780, c2780, in2780_1, in2780_2, pp83[23]);
    wire[0:0] s2781, in2781_1, in2781_2;
    wire c2781;
    assign in2781_1 = {pp87[19]};
    assign in2781_2 = {pp88[18]};
    Full_Adder FA_2781(s2781, c2781, in2781_1, in2781_2, pp86[20]);
    wire[0:0] s2782, in2782_1, in2782_2;
    wire c2782;
    assign in2782_1 = {pp90[16]};
    assign in2782_2 = {pp91[15]};
    Full_Adder FA_2782(s2782, c2782, in2782_1, in2782_2, pp89[17]);
    wire[0:0] s2783, in2783_1, in2783_2;
    wire c2783;
    assign in2783_1 = {pp93[13]};
    assign in2783_2 = {pp94[12]};
    Full_Adder FA_2783(s2783, c2783, in2783_1, in2783_2, pp92[14]);
    wire[0:0] s2784, in2784_1, in2784_2;
    wire c2784;
    assign in2784_1 = {pp96[10]};
    assign in2784_2 = {pp97[9]};
    Full_Adder FA_2784(s2784, c2784, in2784_1, in2784_2, pp95[11]);
    wire[0:0] s2785, in2785_1, in2785_2;
    wire c2785;
    assign in2785_1 = {pp99[7]};
    assign in2785_2 = {pp100[6]};
    Full_Adder FA_2785(s2785, c2785, in2785_1, in2785_2, pp98[8]);
    wire[0:0] s2786, in2786_1, in2786_2;
    wire c2786;
    assign in2786_1 = {pp102[4]};
    assign in2786_2 = {pp103[3]};
    Full_Adder FA_2786(s2786, c2786, in2786_1, in2786_2, pp101[5]);
    wire[0:0] s2787, in2787_1, in2787_2;
    wire c2787;
    assign in2787_1 = {pp105[1]};
    assign in2787_2 = {pp106[0]};
    Full_Adder FA_2787(s2787, c2787, in2787_1, in2787_2, pp104[2]);
    wire[0:0] s2788, in2788_1, in2788_2;
    wire c2788;
    assign in2788_1 = {c192};
    assign in2788_2 = {c193};
    Full_Adder FA_2788(s2788, c2788, in2788_1, in2788_2, c191);
    wire[0:0] s2789, in2789_1, in2789_2;
    wire c2789;
    assign in2789_1 = {c195};
    assign in2789_2 = {c196};
    Full_Adder FA_2789(s2789, c2789, in2789_1, in2789_2, c194);
    wire[0:0] s2790, in2790_1, in2790_2;
    wire c2790;
    assign in2790_1 = {c198};
    assign in2790_2 = {c199};
    Full_Adder FA_2790(s2790, c2790, in2790_1, in2790_2, c197);
    wire[0:0] s2791, in2791_1, in2791_2;
    wire c2791;
    assign in2791_1 = {c201};
    assign in2791_2 = {c202};
    Full_Adder FA_2791(s2791, c2791, in2791_1, in2791_2, c200);
    wire[0:0] s2792, in2792_1, in2792_2;
    wire c2792;
    assign in2792_1 = {c204};
    assign in2792_2 = {c205};
    Full_Adder FA_2792(s2792, c2792, in2792_1, in2792_2, c203);
    wire[0:0] s2793, in2793_1, in2793_2;
    wire c2793;
    assign in2793_1 = {c207};
    assign in2793_2 = {c208};
    Full_Adder FA_2793(s2793, c2793, in2793_1, in2793_2, c206);
    wire[0:0] s2794, in2794_1, in2794_2;
    wire c2794;
    assign in2794_1 = {c210};
    assign in2794_2 = {s211[0]};
    Full_Adder FA_2794(s2794, c2794, in2794_1, in2794_2, c209);
    wire[0:0] s2795, in2795_1, in2795_2;
    wire c2795;
    assign in2795_1 = {s213[0]};
    assign in2795_2 = {s214[0]};
    Full_Adder FA_2795(s2795, c2795, in2795_1, in2795_2, s212[0]);
    wire[0:0] s2796, in2796_1, in2796_2;
    wire c2796;
    assign in2796_1 = {s216[0]};
    assign in2796_2 = {s217[0]};
    Full_Adder FA_2796(s2796, c2796, in2796_1, in2796_2, s215[0]);
    wire[0:0] s2797, in2797_1, in2797_2;
    wire c2797;
    assign in2797_1 = {s219[0]};
    assign in2797_2 = {s220[0]};
    Full_Adder FA_2797(s2797, c2797, in2797_1, in2797_2, s218[0]);
    wire[0:0] s2798, in2798_1, in2798_2;
    wire c2798;
    assign in2798_1 = {s222[0]};
    assign in2798_2 = {s223[0]};
    Full_Adder FA_2798(s2798, c2798, in2798_1, in2798_2, s221[0]);
    wire[0:0] s2799, in2799_1, in2799_2;
    wire c2799;
    assign in2799_1 = {s225[0]};
    assign in2799_2 = {s226[0]};
    Full_Adder FA_2799(s2799, c2799, in2799_1, in2799_2, s224[0]);
    wire[0:0] s2800, in2800_1, in2800_2;
    wire c2800;
    assign in2800_1 = {s228[0]};
    assign in2800_2 = {s229[0]};
    Full_Adder FA_2800(s2800, c2800, in2800_1, in2800_2, s227[0]);
    wire[0:0] s2801, in2801_1, in2801_2;
    wire c2801;
    assign in2801_1 = {pp66[41]};
    assign in2801_2 = {pp67[40]};
    Full_Adder FA_2801(s2801, c2801, in2801_1, in2801_2, pp65[42]);
    wire[0:0] s2802, in2802_1, in2802_2;
    wire c2802;
    assign in2802_1 = {pp69[38]};
    assign in2802_2 = {pp70[37]};
    Full_Adder FA_2802(s2802, c2802, in2802_1, in2802_2, pp68[39]);
    wire[0:0] s2803, in2803_1, in2803_2;
    wire c2803;
    assign in2803_1 = {pp72[35]};
    assign in2803_2 = {pp73[34]};
    Full_Adder FA_2803(s2803, c2803, in2803_1, in2803_2, pp71[36]);
    wire[0:0] s2804, in2804_1, in2804_2;
    wire c2804;
    assign in2804_1 = {pp75[32]};
    assign in2804_2 = {pp76[31]};
    Full_Adder FA_2804(s2804, c2804, in2804_1, in2804_2, pp74[33]);
    wire[0:0] s2805, in2805_1, in2805_2;
    wire c2805;
    assign in2805_1 = {pp78[29]};
    assign in2805_2 = {pp79[28]};
    Full_Adder FA_2805(s2805, c2805, in2805_1, in2805_2, pp77[30]);
    wire[0:0] s2806, in2806_1, in2806_2;
    wire c2806;
    assign in2806_1 = {pp81[26]};
    assign in2806_2 = {pp82[25]};
    Full_Adder FA_2806(s2806, c2806, in2806_1, in2806_2, pp80[27]);
    wire[0:0] s2807, in2807_1, in2807_2;
    wire c2807;
    assign in2807_1 = {pp84[23]};
    assign in2807_2 = {pp85[22]};
    Full_Adder FA_2807(s2807, c2807, in2807_1, in2807_2, pp83[24]);
    wire[0:0] s2808, in2808_1, in2808_2;
    wire c2808;
    assign in2808_1 = {pp87[20]};
    assign in2808_2 = {pp88[19]};
    Full_Adder FA_2808(s2808, c2808, in2808_1, in2808_2, pp86[21]);
    wire[0:0] s2809, in2809_1, in2809_2;
    wire c2809;
    assign in2809_1 = {pp90[17]};
    assign in2809_2 = {pp91[16]};
    Full_Adder FA_2809(s2809, c2809, in2809_1, in2809_2, pp89[18]);
    wire[0:0] s2810, in2810_1, in2810_2;
    wire c2810;
    assign in2810_1 = {pp93[14]};
    assign in2810_2 = {pp94[13]};
    Full_Adder FA_2810(s2810, c2810, in2810_1, in2810_2, pp92[15]);
    wire[0:0] s2811, in2811_1, in2811_2;
    wire c2811;
    assign in2811_1 = {pp96[11]};
    assign in2811_2 = {pp97[10]};
    Full_Adder FA_2811(s2811, c2811, in2811_1, in2811_2, pp95[12]);
    wire[0:0] s2812, in2812_1, in2812_2;
    wire c2812;
    assign in2812_1 = {pp99[8]};
    assign in2812_2 = {pp100[7]};
    Full_Adder FA_2812(s2812, c2812, in2812_1, in2812_2, pp98[9]);
    wire[0:0] s2813, in2813_1, in2813_2;
    wire c2813;
    assign in2813_1 = {pp102[5]};
    assign in2813_2 = {pp103[4]};
    Full_Adder FA_2813(s2813, c2813, in2813_1, in2813_2, pp101[6]);
    wire[0:0] s2814, in2814_1, in2814_2;
    wire c2814;
    assign in2814_1 = {pp105[2]};
    assign in2814_2 = {pp106[1]};
    Full_Adder FA_2814(s2814, c2814, in2814_1, in2814_2, pp104[3]);
    wire[0:0] s2815, in2815_1, in2815_2;
    wire c2815;
    assign in2815_1 = {c211};
    assign in2815_2 = {c212};
    Full_Adder FA_2815(s2815, c2815, in2815_1, in2815_2, pp107[0]);
    wire[0:0] s2816, in2816_1, in2816_2;
    wire c2816;
    assign in2816_1 = {c214};
    assign in2816_2 = {c215};
    Full_Adder FA_2816(s2816, c2816, in2816_1, in2816_2, c213);
    wire[0:0] s2817, in2817_1, in2817_2;
    wire c2817;
    assign in2817_1 = {c217};
    assign in2817_2 = {c218};
    Full_Adder FA_2817(s2817, c2817, in2817_1, in2817_2, c216);
    wire[0:0] s2818, in2818_1, in2818_2;
    wire c2818;
    assign in2818_1 = {c220};
    assign in2818_2 = {c221};
    Full_Adder FA_2818(s2818, c2818, in2818_1, in2818_2, c219);
    wire[0:0] s2819, in2819_1, in2819_2;
    wire c2819;
    assign in2819_1 = {c223};
    assign in2819_2 = {c224};
    Full_Adder FA_2819(s2819, c2819, in2819_1, in2819_2, c222);
    wire[0:0] s2820, in2820_1, in2820_2;
    wire c2820;
    assign in2820_1 = {c226};
    assign in2820_2 = {c227};
    Full_Adder FA_2820(s2820, c2820, in2820_1, in2820_2, c225);
    wire[0:0] s2821, in2821_1, in2821_2;
    wire c2821;
    assign in2821_1 = {c229};
    assign in2821_2 = {c230};
    Full_Adder FA_2821(s2821, c2821, in2821_1, in2821_2, c228);
    wire[0:0] s2822, in2822_1, in2822_2;
    wire c2822;
    assign in2822_1 = {s232[0]};
    assign in2822_2 = {s233[0]};
    Full_Adder FA_2822(s2822, c2822, in2822_1, in2822_2, c231);
    wire[0:0] s2823, in2823_1, in2823_2;
    wire c2823;
    assign in2823_1 = {s235[0]};
    assign in2823_2 = {s236[0]};
    Full_Adder FA_2823(s2823, c2823, in2823_1, in2823_2, s234[0]);
    wire[0:0] s2824, in2824_1, in2824_2;
    wire c2824;
    assign in2824_1 = {s238[0]};
    assign in2824_2 = {s239[0]};
    Full_Adder FA_2824(s2824, c2824, in2824_1, in2824_2, s237[0]);
    wire[0:0] s2825, in2825_1, in2825_2;
    wire c2825;
    assign in2825_1 = {s241[0]};
    assign in2825_2 = {s242[0]};
    Full_Adder FA_2825(s2825, c2825, in2825_1, in2825_2, s240[0]);
    wire[0:0] s2826, in2826_1, in2826_2;
    wire c2826;
    assign in2826_1 = {s244[0]};
    assign in2826_2 = {s245[0]};
    Full_Adder FA_2826(s2826, c2826, in2826_1, in2826_2, s243[0]);
    wire[0:0] s2827, in2827_1, in2827_2;
    wire c2827;
    assign in2827_1 = {s247[0]};
    assign in2827_2 = {s248[0]};
    Full_Adder FA_2827(s2827, c2827, in2827_1, in2827_2, s246[0]);
    wire[0:0] s2828, in2828_1, in2828_2;
    wire c2828;
    assign in2828_1 = {s250[0]};
    assign in2828_2 = {s251[0]};
    Full_Adder FA_2828(s2828, c2828, in2828_1, in2828_2, s249[0]);
    wire[0:0] s2829, in2829_1, in2829_2;
    wire c2829;
    assign in2829_1 = {pp69[39]};
    assign in2829_2 = {pp70[38]};
    Full_Adder FA_2829(s2829, c2829, in2829_1, in2829_2, pp68[40]);
    wire[0:0] s2830, in2830_1, in2830_2;
    wire c2830;
    assign in2830_1 = {pp72[36]};
    assign in2830_2 = {pp73[35]};
    Full_Adder FA_2830(s2830, c2830, in2830_1, in2830_2, pp71[37]);
    wire[0:0] s2831, in2831_1, in2831_2;
    wire c2831;
    assign in2831_1 = {pp75[33]};
    assign in2831_2 = {pp76[32]};
    Full_Adder FA_2831(s2831, c2831, in2831_1, in2831_2, pp74[34]);
    wire[0:0] s2832, in2832_1, in2832_2;
    wire c2832;
    assign in2832_1 = {pp78[30]};
    assign in2832_2 = {pp79[29]};
    Full_Adder FA_2832(s2832, c2832, in2832_1, in2832_2, pp77[31]);
    wire[0:0] s2833, in2833_1, in2833_2;
    wire c2833;
    assign in2833_1 = {pp81[27]};
    assign in2833_2 = {pp82[26]};
    Full_Adder FA_2833(s2833, c2833, in2833_1, in2833_2, pp80[28]);
    wire[0:0] s2834, in2834_1, in2834_2;
    wire c2834;
    assign in2834_1 = {pp84[24]};
    assign in2834_2 = {pp85[23]};
    Full_Adder FA_2834(s2834, c2834, in2834_1, in2834_2, pp83[25]);
    wire[0:0] s2835, in2835_1, in2835_2;
    wire c2835;
    assign in2835_1 = {pp87[21]};
    assign in2835_2 = {pp88[20]};
    Full_Adder FA_2835(s2835, c2835, in2835_1, in2835_2, pp86[22]);
    wire[0:0] s2836, in2836_1, in2836_2;
    wire c2836;
    assign in2836_1 = {pp90[18]};
    assign in2836_2 = {pp91[17]};
    Full_Adder FA_2836(s2836, c2836, in2836_1, in2836_2, pp89[19]);
    wire[0:0] s2837, in2837_1, in2837_2;
    wire c2837;
    assign in2837_1 = {pp93[15]};
    assign in2837_2 = {pp94[14]};
    Full_Adder FA_2837(s2837, c2837, in2837_1, in2837_2, pp92[16]);
    wire[0:0] s2838, in2838_1, in2838_2;
    wire c2838;
    assign in2838_1 = {pp96[12]};
    assign in2838_2 = {pp97[11]};
    Full_Adder FA_2838(s2838, c2838, in2838_1, in2838_2, pp95[13]);
    wire[0:0] s2839, in2839_1, in2839_2;
    wire c2839;
    assign in2839_1 = {pp99[9]};
    assign in2839_2 = {pp100[8]};
    Full_Adder FA_2839(s2839, c2839, in2839_1, in2839_2, pp98[10]);
    wire[0:0] s2840, in2840_1, in2840_2;
    wire c2840;
    assign in2840_1 = {pp102[6]};
    assign in2840_2 = {pp103[5]};
    Full_Adder FA_2840(s2840, c2840, in2840_1, in2840_2, pp101[7]);
    wire[0:0] s2841, in2841_1, in2841_2;
    wire c2841;
    assign in2841_1 = {pp105[3]};
    assign in2841_2 = {pp106[2]};
    Full_Adder FA_2841(s2841, c2841, in2841_1, in2841_2, pp104[4]);
    wire[0:0] s2842, in2842_1, in2842_2;
    wire c2842;
    assign in2842_1 = {pp108[0]};
    assign in2842_2 = {c232};
    Full_Adder FA_2842(s2842, c2842, in2842_1, in2842_2, pp107[1]);
    wire[0:0] s2843, in2843_1, in2843_2;
    wire c2843;
    assign in2843_1 = {c234};
    assign in2843_2 = {c235};
    Full_Adder FA_2843(s2843, c2843, in2843_1, in2843_2, c233);
    wire[0:0] s2844, in2844_1, in2844_2;
    wire c2844;
    assign in2844_1 = {c237};
    assign in2844_2 = {c238};
    Full_Adder FA_2844(s2844, c2844, in2844_1, in2844_2, c236);
    wire[0:0] s2845, in2845_1, in2845_2;
    wire c2845;
    assign in2845_1 = {c240};
    assign in2845_2 = {c241};
    Full_Adder FA_2845(s2845, c2845, in2845_1, in2845_2, c239);
    wire[0:0] s2846, in2846_1, in2846_2;
    wire c2846;
    assign in2846_1 = {c243};
    assign in2846_2 = {c244};
    Full_Adder FA_2846(s2846, c2846, in2846_1, in2846_2, c242);
    wire[0:0] s2847, in2847_1, in2847_2;
    wire c2847;
    assign in2847_1 = {c246};
    assign in2847_2 = {c247};
    Full_Adder FA_2847(s2847, c2847, in2847_1, in2847_2, c245);
    wire[0:0] s2848, in2848_1, in2848_2;
    wire c2848;
    assign in2848_1 = {c249};
    assign in2848_2 = {c250};
    Full_Adder FA_2848(s2848, c2848, in2848_1, in2848_2, c248);
    wire[0:0] s2849, in2849_1, in2849_2;
    wire c2849;
    assign in2849_1 = {c252};
    assign in2849_2 = {c253};
    Full_Adder FA_2849(s2849, c2849, in2849_1, in2849_2, c251);
    wire[0:0] s2850, in2850_1, in2850_2;
    wire c2850;
    assign in2850_1 = {s255[0]};
    assign in2850_2 = {s256[0]};
    Full_Adder FA_2850(s2850, c2850, in2850_1, in2850_2, s254[0]);
    wire[0:0] s2851, in2851_1, in2851_2;
    wire c2851;
    assign in2851_1 = {s258[0]};
    assign in2851_2 = {s259[0]};
    Full_Adder FA_2851(s2851, c2851, in2851_1, in2851_2, s257[0]);
    wire[0:0] s2852, in2852_1, in2852_2;
    wire c2852;
    assign in2852_1 = {s261[0]};
    assign in2852_2 = {s262[0]};
    Full_Adder FA_2852(s2852, c2852, in2852_1, in2852_2, s260[0]);
    wire[0:0] s2853, in2853_1, in2853_2;
    wire c2853;
    assign in2853_1 = {s264[0]};
    assign in2853_2 = {s265[0]};
    Full_Adder FA_2853(s2853, c2853, in2853_1, in2853_2, s263[0]);
    wire[0:0] s2854, in2854_1, in2854_2;
    wire c2854;
    assign in2854_1 = {s267[0]};
    assign in2854_2 = {s268[0]};
    Full_Adder FA_2854(s2854, c2854, in2854_1, in2854_2, s266[0]);
    wire[0:0] s2855, in2855_1, in2855_2;
    wire c2855;
    assign in2855_1 = {s270[0]};
    assign in2855_2 = {s271[0]};
    Full_Adder FA_2855(s2855, c2855, in2855_1, in2855_2, s269[0]);
    wire[0:0] s2856, in2856_1, in2856_2;
    wire c2856;
    assign in2856_1 = {s273[0]};
    assign in2856_2 = {s274[0]};
    Full_Adder FA_2856(s2856, c2856, in2856_1, in2856_2, s272[0]);
    wire[0:0] s2857, in2857_1, in2857_2;
    wire c2857;
    assign in2857_1 = {pp72[37]};
    assign in2857_2 = {pp73[36]};
    Full_Adder FA_2857(s2857, c2857, in2857_1, in2857_2, pp71[38]);
    wire[0:0] s2858, in2858_1, in2858_2;
    wire c2858;
    assign in2858_1 = {pp75[34]};
    assign in2858_2 = {pp76[33]};
    Full_Adder FA_2858(s2858, c2858, in2858_1, in2858_2, pp74[35]);
    wire[0:0] s2859, in2859_1, in2859_2;
    wire c2859;
    assign in2859_1 = {pp78[31]};
    assign in2859_2 = {pp79[30]};
    Full_Adder FA_2859(s2859, c2859, in2859_1, in2859_2, pp77[32]);
    wire[0:0] s2860, in2860_1, in2860_2;
    wire c2860;
    assign in2860_1 = {pp81[28]};
    assign in2860_2 = {pp82[27]};
    Full_Adder FA_2860(s2860, c2860, in2860_1, in2860_2, pp80[29]);
    wire[0:0] s2861, in2861_1, in2861_2;
    wire c2861;
    assign in2861_1 = {pp84[25]};
    assign in2861_2 = {pp85[24]};
    Full_Adder FA_2861(s2861, c2861, in2861_1, in2861_2, pp83[26]);
    wire[0:0] s2862, in2862_1, in2862_2;
    wire c2862;
    assign in2862_1 = {pp87[22]};
    assign in2862_2 = {pp88[21]};
    Full_Adder FA_2862(s2862, c2862, in2862_1, in2862_2, pp86[23]);
    wire[0:0] s2863, in2863_1, in2863_2;
    wire c2863;
    assign in2863_1 = {pp90[19]};
    assign in2863_2 = {pp91[18]};
    Full_Adder FA_2863(s2863, c2863, in2863_1, in2863_2, pp89[20]);
    wire[0:0] s2864, in2864_1, in2864_2;
    wire c2864;
    assign in2864_1 = {pp93[16]};
    assign in2864_2 = {pp94[15]};
    Full_Adder FA_2864(s2864, c2864, in2864_1, in2864_2, pp92[17]);
    wire[0:0] s2865, in2865_1, in2865_2;
    wire c2865;
    assign in2865_1 = {pp96[13]};
    assign in2865_2 = {pp97[12]};
    Full_Adder FA_2865(s2865, c2865, in2865_1, in2865_2, pp95[14]);
    wire[0:0] s2866, in2866_1, in2866_2;
    wire c2866;
    assign in2866_1 = {pp99[10]};
    assign in2866_2 = {pp100[9]};
    Full_Adder FA_2866(s2866, c2866, in2866_1, in2866_2, pp98[11]);
    wire[0:0] s2867, in2867_1, in2867_2;
    wire c2867;
    assign in2867_1 = {pp102[7]};
    assign in2867_2 = {pp103[6]};
    Full_Adder FA_2867(s2867, c2867, in2867_1, in2867_2, pp101[8]);
    wire[0:0] s2868, in2868_1, in2868_2;
    wire c2868;
    assign in2868_1 = {pp105[4]};
    assign in2868_2 = {pp106[3]};
    Full_Adder FA_2868(s2868, c2868, in2868_1, in2868_2, pp104[5]);
    wire[0:0] s2869, in2869_1, in2869_2;
    wire c2869;
    assign in2869_1 = {pp108[1]};
    assign in2869_2 = {pp109[0]};
    Full_Adder FA_2869(s2869, c2869, in2869_1, in2869_2, pp107[2]);
    wire[0:0] s2870, in2870_1, in2870_2;
    wire c2870;
    assign in2870_1 = {c255};
    assign in2870_2 = {c256};
    Full_Adder FA_2870(s2870, c2870, in2870_1, in2870_2, c254);
    wire[0:0] s2871, in2871_1, in2871_2;
    wire c2871;
    assign in2871_1 = {c258};
    assign in2871_2 = {c259};
    Full_Adder FA_2871(s2871, c2871, in2871_1, in2871_2, c257);
    wire[0:0] s2872, in2872_1, in2872_2;
    wire c2872;
    assign in2872_1 = {c261};
    assign in2872_2 = {c262};
    Full_Adder FA_2872(s2872, c2872, in2872_1, in2872_2, c260);
    wire[0:0] s2873, in2873_1, in2873_2;
    wire c2873;
    assign in2873_1 = {c264};
    assign in2873_2 = {c265};
    Full_Adder FA_2873(s2873, c2873, in2873_1, in2873_2, c263);
    wire[0:0] s2874, in2874_1, in2874_2;
    wire c2874;
    assign in2874_1 = {c267};
    assign in2874_2 = {c268};
    Full_Adder FA_2874(s2874, c2874, in2874_1, in2874_2, c266);
    wire[0:0] s2875, in2875_1, in2875_2;
    wire c2875;
    assign in2875_1 = {c270};
    assign in2875_2 = {c271};
    Full_Adder FA_2875(s2875, c2875, in2875_1, in2875_2, c269);
    wire[0:0] s2876, in2876_1, in2876_2;
    wire c2876;
    assign in2876_1 = {c273};
    assign in2876_2 = {c274};
    Full_Adder FA_2876(s2876, c2876, in2876_1, in2876_2, c272);
    wire[0:0] s2877, in2877_1, in2877_2;
    wire c2877;
    assign in2877_1 = {c276};
    assign in2877_2 = {s277[0]};
    Full_Adder FA_2877(s2877, c2877, in2877_1, in2877_2, c275);
    wire[0:0] s2878, in2878_1, in2878_2;
    wire c2878;
    assign in2878_1 = {s279[0]};
    assign in2878_2 = {s280[0]};
    Full_Adder FA_2878(s2878, c2878, in2878_1, in2878_2, s278[0]);
    wire[0:0] s2879, in2879_1, in2879_2;
    wire c2879;
    assign in2879_1 = {s282[0]};
    assign in2879_2 = {s283[0]};
    Full_Adder FA_2879(s2879, c2879, in2879_1, in2879_2, s281[0]);
    wire[0:0] s2880, in2880_1, in2880_2;
    wire c2880;
    assign in2880_1 = {s285[0]};
    assign in2880_2 = {s286[0]};
    Full_Adder FA_2880(s2880, c2880, in2880_1, in2880_2, s284[0]);
    wire[0:0] s2881, in2881_1, in2881_2;
    wire c2881;
    assign in2881_1 = {s288[0]};
    assign in2881_2 = {s289[0]};
    Full_Adder FA_2881(s2881, c2881, in2881_1, in2881_2, s287[0]);
    wire[0:0] s2882, in2882_1, in2882_2;
    wire c2882;
    assign in2882_1 = {s291[0]};
    assign in2882_2 = {s292[0]};
    Full_Adder FA_2882(s2882, c2882, in2882_1, in2882_2, s290[0]);
    wire[0:0] s2883, in2883_1, in2883_2;
    wire c2883;
    assign in2883_1 = {s294[0]};
    assign in2883_2 = {s295[0]};
    Full_Adder FA_2883(s2883, c2883, in2883_1, in2883_2, s293[0]);
    wire[0:0] s2884, in2884_1, in2884_2;
    wire c2884;
    assign in2884_1 = {s297[0]};
    assign in2884_2 = {s298[0]};
    Full_Adder FA_2884(s2884, c2884, in2884_1, in2884_2, s296[0]);
    wire[0:0] s2885, in2885_1, in2885_2;
    wire c2885;
    assign in2885_1 = {pp75[35]};
    assign in2885_2 = {pp76[34]};
    Full_Adder FA_2885(s2885, c2885, in2885_1, in2885_2, pp74[36]);
    wire[0:0] s2886, in2886_1, in2886_2;
    wire c2886;
    assign in2886_1 = {pp78[32]};
    assign in2886_2 = {pp79[31]};
    Full_Adder FA_2886(s2886, c2886, in2886_1, in2886_2, pp77[33]);
    wire[0:0] s2887, in2887_1, in2887_2;
    wire c2887;
    assign in2887_1 = {pp81[29]};
    assign in2887_2 = {pp82[28]};
    Full_Adder FA_2887(s2887, c2887, in2887_1, in2887_2, pp80[30]);
    wire[0:0] s2888, in2888_1, in2888_2;
    wire c2888;
    assign in2888_1 = {pp84[26]};
    assign in2888_2 = {pp85[25]};
    Full_Adder FA_2888(s2888, c2888, in2888_1, in2888_2, pp83[27]);
    wire[0:0] s2889, in2889_1, in2889_2;
    wire c2889;
    assign in2889_1 = {pp87[23]};
    assign in2889_2 = {pp88[22]};
    Full_Adder FA_2889(s2889, c2889, in2889_1, in2889_2, pp86[24]);
    wire[0:0] s2890, in2890_1, in2890_2;
    wire c2890;
    assign in2890_1 = {pp90[20]};
    assign in2890_2 = {pp91[19]};
    Full_Adder FA_2890(s2890, c2890, in2890_1, in2890_2, pp89[21]);
    wire[0:0] s2891, in2891_1, in2891_2;
    wire c2891;
    assign in2891_1 = {pp93[17]};
    assign in2891_2 = {pp94[16]};
    Full_Adder FA_2891(s2891, c2891, in2891_1, in2891_2, pp92[18]);
    wire[0:0] s2892, in2892_1, in2892_2;
    wire c2892;
    assign in2892_1 = {pp96[14]};
    assign in2892_2 = {pp97[13]};
    Full_Adder FA_2892(s2892, c2892, in2892_1, in2892_2, pp95[15]);
    wire[0:0] s2893, in2893_1, in2893_2;
    wire c2893;
    assign in2893_1 = {pp99[11]};
    assign in2893_2 = {pp100[10]};
    Full_Adder FA_2893(s2893, c2893, in2893_1, in2893_2, pp98[12]);
    wire[0:0] s2894, in2894_1, in2894_2;
    wire c2894;
    assign in2894_1 = {pp102[8]};
    assign in2894_2 = {pp103[7]};
    Full_Adder FA_2894(s2894, c2894, in2894_1, in2894_2, pp101[9]);
    wire[0:0] s2895, in2895_1, in2895_2;
    wire c2895;
    assign in2895_1 = {pp105[5]};
    assign in2895_2 = {pp106[4]};
    Full_Adder FA_2895(s2895, c2895, in2895_1, in2895_2, pp104[6]);
    wire[0:0] s2896, in2896_1, in2896_2;
    wire c2896;
    assign in2896_1 = {pp108[2]};
    assign in2896_2 = {pp109[1]};
    Full_Adder FA_2896(s2896, c2896, in2896_1, in2896_2, pp107[3]);
    wire[0:0] s2897, in2897_1, in2897_2;
    wire c2897;
    assign in2897_1 = {c277};
    assign in2897_2 = {c278};
    Full_Adder FA_2897(s2897, c2897, in2897_1, in2897_2, pp110[0]);
    wire[0:0] s2898, in2898_1, in2898_2;
    wire c2898;
    assign in2898_1 = {c280};
    assign in2898_2 = {c281};
    Full_Adder FA_2898(s2898, c2898, in2898_1, in2898_2, c279);
    wire[0:0] s2899, in2899_1, in2899_2;
    wire c2899;
    assign in2899_1 = {c283};
    assign in2899_2 = {c284};
    Full_Adder FA_2899(s2899, c2899, in2899_1, in2899_2, c282);
    wire[0:0] s2900, in2900_1, in2900_2;
    wire c2900;
    assign in2900_1 = {c286};
    assign in2900_2 = {c287};
    Full_Adder FA_2900(s2900, c2900, in2900_1, in2900_2, c285);
    wire[0:0] s2901, in2901_1, in2901_2;
    wire c2901;
    assign in2901_1 = {c289};
    assign in2901_2 = {c290};
    Full_Adder FA_2901(s2901, c2901, in2901_1, in2901_2, c288);
    wire[0:0] s2902, in2902_1, in2902_2;
    wire c2902;
    assign in2902_1 = {c292};
    assign in2902_2 = {c293};
    Full_Adder FA_2902(s2902, c2902, in2902_1, in2902_2, c291);
    wire[0:0] s2903, in2903_1, in2903_2;
    wire c2903;
    assign in2903_1 = {c295};
    assign in2903_2 = {c296};
    Full_Adder FA_2903(s2903, c2903, in2903_1, in2903_2, c294);
    wire[0:0] s2904, in2904_1, in2904_2;
    wire c2904;
    assign in2904_1 = {c298};
    assign in2904_2 = {c299};
    Full_Adder FA_2904(s2904, c2904, in2904_1, in2904_2, c297);
    wire[0:0] s2905, in2905_1, in2905_2;
    wire c2905;
    assign in2905_1 = {s301[0]};
    assign in2905_2 = {s302[0]};
    Full_Adder FA_2905(s2905, c2905, in2905_1, in2905_2, c300);
    wire[0:0] s2906, in2906_1, in2906_2;
    wire c2906;
    assign in2906_1 = {s304[0]};
    assign in2906_2 = {s305[0]};
    Full_Adder FA_2906(s2906, c2906, in2906_1, in2906_2, s303[0]);
    wire[0:0] s2907, in2907_1, in2907_2;
    wire c2907;
    assign in2907_1 = {s307[0]};
    assign in2907_2 = {s308[0]};
    Full_Adder FA_2907(s2907, c2907, in2907_1, in2907_2, s306[0]);
    wire[0:0] s2908, in2908_1, in2908_2;
    wire c2908;
    assign in2908_1 = {s310[0]};
    assign in2908_2 = {s311[0]};
    Full_Adder FA_2908(s2908, c2908, in2908_1, in2908_2, s309[0]);
    wire[0:0] s2909, in2909_1, in2909_2;
    wire c2909;
    assign in2909_1 = {s313[0]};
    assign in2909_2 = {s314[0]};
    Full_Adder FA_2909(s2909, c2909, in2909_1, in2909_2, s312[0]);
    wire[0:0] s2910, in2910_1, in2910_2;
    wire c2910;
    assign in2910_1 = {s316[0]};
    assign in2910_2 = {s317[0]};
    Full_Adder FA_2910(s2910, c2910, in2910_1, in2910_2, s315[0]);
    wire[0:0] s2911, in2911_1, in2911_2;
    wire c2911;
    assign in2911_1 = {s319[0]};
    assign in2911_2 = {s320[0]};
    Full_Adder FA_2911(s2911, c2911, in2911_1, in2911_2, s318[0]);
    wire[0:0] s2912, in2912_1, in2912_2;
    wire c2912;
    assign in2912_1 = {s322[0]};
    assign in2912_2 = {s323[0]};
    Full_Adder FA_2912(s2912, c2912, in2912_1, in2912_2, s321[0]);
    wire[0:0] s2913, in2913_1, in2913_2;
    wire c2913;
    assign in2913_1 = {pp78[33]};
    assign in2913_2 = {pp79[32]};
    Full_Adder FA_2913(s2913, c2913, in2913_1, in2913_2, pp77[34]);
    wire[0:0] s2914, in2914_1, in2914_2;
    wire c2914;
    assign in2914_1 = {pp81[30]};
    assign in2914_2 = {pp82[29]};
    Full_Adder FA_2914(s2914, c2914, in2914_1, in2914_2, pp80[31]);
    wire[0:0] s2915, in2915_1, in2915_2;
    wire c2915;
    assign in2915_1 = {pp84[27]};
    assign in2915_2 = {pp85[26]};
    Full_Adder FA_2915(s2915, c2915, in2915_1, in2915_2, pp83[28]);
    wire[0:0] s2916, in2916_1, in2916_2;
    wire c2916;
    assign in2916_1 = {pp87[24]};
    assign in2916_2 = {pp88[23]};
    Full_Adder FA_2916(s2916, c2916, in2916_1, in2916_2, pp86[25]);
    wire[0:0] s2917, in2917_1, in2917_2;
    wire c2917;
    assign in2917_1 = {pp90[21]};
    assign in2917_2 = {pp91[20]};
    Full_Adder FA_2917(s2917, c2917, in2917_1, in2917_2, pp89[22]);
    wire[0:0] s2918, in2918_1, in2918_2;
    wire c2918;
    assign in2918_1 = {pp93[18]};
    assign in2918_2 = {pp94[17]};
    Full_Adder FA_2918(s2918, c2918, in2918_1, in2918_2, pp92[19]);
    wire[0:0] s2919, in2919_1, in2919_2;
    wire c2919;
    assign in2919_1 = {pp96[15]};
    assign in2919_2 = {pp97[14]};
    Full_Adder FA_2919(s2919, c2919, in2919_1, in2919_2, pp95[16]);
    wire[0:0] s2920, in2920_1, in2920_2;
    wire c2920;
    assign in2920_1 = {pp99[12]};
    assign in2920_2 = {pp100[11]};
    Full_Adder FA_2920(s2920, c2920, in2920_1, in2920_2, pp98[13]);
    wire[0:0] s2921, in2921_1, in2921_2;
    wire c2921;
    assign in2921_1 = {pp102[9]};
    assign in2921_2 = {pp103[8]};
    Full_Adder FA_2921(s2921, c2921, in2921_1, in2921_2, pp101[10]);
    wire[0:0] s2922, in2922_1, in2922_2;
    wire c2922;
    assign in2922_1 = {pp105[6]};
    assign in2922_2 = {pp106[5]};
    Full_Adder FA_2922(s2922, c2922, in2922_1, in2922_2, pp104[7]);
    wire[0:0] s2923, in2923_1, in2923_2;
    wire c2923;
    assign in2923_1 = {pp108[3]};
    assign in2923_2 = {pp109[2]};
    Full_Adder FA_2923(s2923, c2923, in2923_1, in2923_2, pp107[4]);
    wire[0:0] s2924, in2924_1, in2924_2;
    wire c2924;
    assign in2924_1 = {pp111[0]};
    assign in2924_2 = {c301};
    Full_Adder FA_2924(s2924, c2924, in2924_1, in2924_2, pp110[1]);
    wire[0:0] s2925, in2925_1, in2925_2;
    wire c2925;
    assign in2925_1 = {c303};
    assign in2925_2 = {c304};
    Full_Adder FA_2925(s2925, c2925, in2925_1, in2925_2, c302);
    wire[0:0] s2926, in2926_1, in2926_2;
    wire c2926;
    assign in2926_1 = {c306};
    assign in2926_2 = {c307};
    Full_Adder FA_2926(s2926, c2926, in2926_1, in2926_2, c305);
    wire[0:0] s2927, in2927_1, in2927_2;
    wire c2927;
    assign in2927_1 = {c309};
    assign in2927_2 = {c310};
    Full_Adder FA_2927(s2927, c2927, in2927_1, in2927_2, c308);
    wire[0:0] s2928, in2928_1, in2928_2;
    wire c2928;
    assign in2928_1 = {c312};
    assign in2928_2 = {c313};
    Full_Adder FA_2928(s2928, c2928, in2928_1, in2928_2, c311);
    wire[0:0] s2929, in2929_1, in2929_2;
    wire c2929;
    assign in2929_1 = {c315};
    assign in2929_2 = {c316};
    Full_Adder FA_2929(s2929, c2929, in2929_1, in2929_2, c314);
    wire[0:0] s2930, in2930_1, in2930_2;
    wire c2930;
    assign in2930_1 = {c318};
    assign in2930_2 = {c319};
    Full_Adder FA_2930(s2930, c2930, in2930_1, in2930_2, c317);
    wire[0:0] s2931, in2931_1, in2931_2;
    wire c2931;
    assign in2931_1 = {c321};
    assign in2931_2 = {c322};
    Full_Adder FA_2931(s2931, c2931, in2931_1, in2931_2, c320);
    wire[0:0] s2932, in2932_1, in2932_2;
    wire c2932;
    assign in2932_1 = {c324};
    assign in2932_2 = {c325};
    Full_Adder FA_2932(s2932, c2932, in2932_1, in2932_2, c323);
    wire[0:0] s2933, in2933_1, in2933_2;
    wire c2933;
    assign in2933_1 = {s327[0]};
    assign in2933_2 = {s328[0]};
    Full_Adder FA_2933(s2933, c2933, in2933_1, in2933_2, s326[0]);
    wire[0:0] s2934, in2934_1, in2934_2;
    wire c2934;
    assign in2934_1 = {s330[0]};
    assign in2934_2 = {s331[0]};
    Full_Adder FA_2934(s2934, c2934, in2934_1, in2934_2, s329[0]);
    wire[0:0] s2935, in2935_1, in2935_2;
    wire c2935;
    assign in2935_1 = {s333[0]};
    assign in2935_2 = {s334[0]};
    Full_Adder FA_2935(s2935, c2935, in2935_1, in2935_2, s332[0]);
    wire[0:0] s2936, in2936_1, in2936_2;
    wire c2936;
    assign in2936_1 = {s336[0]};
    assign in2936_2 = {s337[0]};
    Full_Adder FA_2936(s2936, c2936, in2936_1, in2936_2, s335[0]);
    wire[0:0] s2937, in2937_1, in2937_2;
    wire c2937;
    assign in2937_1 = {s339[0]};
    assign in2937_2 = {s340[0]};
    Full_Adder FA_2937(s2937, c2937, in2937_1, in2937_2, s338[0]);
    wire[0:0] s2938, in2938_1, in2938_2;
    wire c2938;
    assign in2938_1 = {s342[0]};
    assign in2938_2 = {s343[0]};
    Full_Adder FA_2938(s2938, c2938, in2938_1, in2938_2, s341[0]);
    wire[0:0] s2939, in2939_1, in2939_2;
    wire c2939;
    assign in2939_1 = {s345[0]};
    assign in2939_2 = {s346[0]};
    Full_Adder FA_2939(s2939, c2939, in2939_1, in2939_2, s344[0]);
    wire[0:0] s2940, in2940_1, in2940_2;
    wire c2940;
    assign in2940_1 = {s348[0]};
    assign in2940_2 = {s349[0]};
    Full_Adder FA_2940(s2940, c2940, in2940_1, in2940_2, s347[0]);
    wire[0:0] s2941, in2941_1, in2941_2;
    wire c2941;
    assign in2941_1 = {pp81[31]};
    assign in2941_2 = {pp82[30]};
    Full_Adder FA_2941(s2941, c2941, in2941_1, in2941_2, pp80[32]);
    wire[0:0] s2942, in2942_1, in2942_2;
    wire c2942;
    assign in2942_1 = {pp84[28]};
    assign in2942_2 = {pp85[27]};
    Full_Adder FA_2942(s2942, c2942, in2942_1, in2942_2, pp83[29]);
    wire[0:0] s2943, in2943_1, in2943_2;
    wire c2943;
    assign in2943_1 = {pp87[25]};
    assign in2943_2 = {pp88[24]};
    Full_Adder FA_2943(s2943, c2943, in2943_1, in2943_2, pp86[26]);
    wire[0:0] s2944, in2944_1, in2944_2;
    wire c2944;
    assign in2944_1 = {pp90[22]};
    assign in2944_2 = {pp91[21]};
    Full_Adder FA_2944(s2944, c2944, in2944_1, in2944_2, pp89[23]);
    wire[0:0] s2945, in2945_1, in2945_2;
    wire c2945;
    assign in2945_1 = {pp93[19]};
    assign in2945_2 = {pp94[18]};
    Full_Adder FA_2945(s2945, c2945, in2945_1, in2945_2, pp92[20]);
    wire[0:0] s2946, in2946_1, in2946_2;
    wire c2946;
    assign in2946_1 = {pp96[16]};
    assign in2946_2 = {pp97[15]};
    Full_Adder FA_2946(s2946, c2946, in2946_1, in2946_2, pp95[17]);
    wire[0:0] s2947, in2947_1, in2947_2;
    wire c2947;
    assign in2947_1 = {pp99[13]};
    assign in2947_2 = {pp100[12]};
    Full_Adder FA_2947(s2947, c2947, in2947_1, in2947_2, pp98[14]);
    wire[0:0] s2948, in2948_1, in2948_2;
    wire c2948;
    assign in2948_1 = {pp102[10]};
    assign in2948_2 = {pp103[9]};
    Full_Adder FA_2948(s2948, c2948, in2948_1, in2948_2, pp101[11]);
    wire[0:0] s2949, in2949_1, in2949_2;
    wire c2949;
    assign in2949_1 = {pp105[7]};
    assign in2949_2 = {pp106[6]};
    Full_Adder FA_2949(s2949, c2949, in2949_1, in2949_2, pp104[8]);
    wire[0:0] s2950, in2950_1, in2950_2;
    wire c2950;
    assign in2950_1 = {pp108[4]};
    assign in2950_2 = {pp109[3]};
    Full_Adder FA_2950(s2950, c2950, in2950_1, in2950_2, pp107[5]);
    wire[0:0] s2951, in2951_1, in2951_2;
    wire c2951;
    assign in2951_1 = {pp111[1]};
    assign in2951_2 = {pp112[0]};
    Full_Adder FA_2951(s2951, c2951, in2951_1, in2951_2, pp110[2]);
    wire[0:0] s2952, in2952_1, in2952_2;
    wire c2952;
    assign in2952_1 = {c327};
    assign in2952_2 = {c328};
    Full_Adder FA_2952(s2952, c2952, in2952_1, in2952_2, c326);
    wire[0:0] s2953, in2953_1, in2953_2;
    wire c2953;
    assign in2953_1 = {c330};
    assign in2953_2 = {c331};
    Full_Adder FA_2953(s2953, c2953, in2953_1, in2953_2, c329);
    wire[0:0] s2954, in2954_1, in2954_2;
    wire c2954;
    assign in2954_1 = {c333};
    assign in2954_2 = {c334};
    Full_Adder FA_2954(s2954, c2954, in2954_1, in2954_2, c332);
    wire[0:0] s2955, in2955_1, in2955_2;
    wire c2955;
    assign in2955_1 = {c336};
    assign in2955_2 = {c337};
    Full_Adder FA_2955(s2955, c2955, in2955_1, in2955_2, c335);
    wire[0:0] s2956, in2956_1, in2956_2;
    wire c2956;
    assign in2956_1 = {c339};
    assign in2956_2 = {c340};
    Full_Adder FA_2956(s2956, c2956, in2956_1, in2956_2, c338);
    wire[0:0] s2957, in2957_1, in2957_2;
    wire c2957;
    assign in2957_1 = {c342};
    assign in2957_2 = {c343};
    Full_Adder FA_2957(s2957, c2957, in2957_1, in2957_2, c341);
    wire[0:0] s2958, in2958_1, in2958_2;
    wire c2958;
    assign in2958_1 = {c345};
    assign in2958_2 = {c346};
    Full_Adder FA_2958(s2958, c2958, in2958_1, in2958_2, c344);
    wire[0:0] s2959, in2959_1, in2959_2;
    wire c2959;
    assign in2959_1 = {c348};
    assign in2959_2 = {c349};
    Full_Adder FA_2959(s2959, c2959, in2959_1, in2959_2, c347);
    wire[0:0] s2960, in2960_1, in2960_2;
    wire c2960;
    assign in2960_1 = {c351};
    assign in2960_2 = {s352[0]};
    Full_Adder FA_2960(s2960, c2960, in2960_1, in2960_2, c350);
    wire[0:0] s2961, in2961_1, in2961_2;
    wire c2961;
    assign in2961_1 = {s354[0]};
    assign in2961_2 = {s355[0]};
    Full_Adder FA_2961(s2961, c2961, in2961_1, in2961_2, s353[0]);
    wire[0:0] s2962, in2962_1, in2962_2;
    wire c2962;
    assign in2962_1 = {s357[0]};
    assign in2962_2 = {s358[0]};
    Full_Adder FA_2962(s2962, c2962, in2962_1, in2962_2, s356[0]);
    wire[0:0] s2963, in2963_1, in2963_2;
    wire c2963;
    assign in2963_1 = {s360[0]};
    assign in2963_2 = {s361[0]};
    Full_Adder FA_2963(s2963, c2963, in2963_1, in2963_2, s359[0]);
    wire[0:0] s2964, in2964_1, in2964_2;
    wire c2964;
    assign in2964_1 = {s363[0]};
    assign in2964_2 = {s364[0]};
    Full_Adder FA_2964(s2964, c2964, in2964_1, in2964_2, s362[0]);
    wire[0:0] s2965, in2965_1, in2965_2;
    wire c2965;
    assign in2965_1 = {s366[0]};
    assign in2965_2 = {s367[0]};
    Full_Adder FA_2965(s2965, c2965, in2965_1, in2965_2, s365[0]);
    wire[0:0] s2966, in2966_1, in2966_2;
    wire c2966;
    assign in2966_1 = {s369[0]};
    assign in2966_2 = {s370[0]};
    Full_Adder FA_2966(s2966, c2966, in2966_1, in2966_2, s368[0]);
    wire[0:0] s2967, in2967_1, in2967_2;
    wire c2967;
    assign in2967_1 = {s372[0]};
    assign in2967_2 = {s373[0]};
    Full_Adder FA_2967(s2967, c2967, in2967_1, in2967_2, s371[0]);
    wire[0:0] s2968, in2968_1, in2968_2;
    wire c2968;
    assign in2968_1 = {s375[0]};
    assign in2968_2 = {s376[0]};
    Full_Adder FA_2968(s2968, c2968, in2968_1, in2968_2, s374[0]);
    wire[0:0] s2969, in2969_1, in2969_2;
    wire c2969;
    assign in2969_1 = {pp84[29]};
    assign in2969_2 = {pp85[28]};
    Full_Adder FA_2969(s2969, c2969, in2969_1, in2969_2, pp83[30]);
    wire[0:0] s2970, in2970_1, in2970_2;
    wire c2970;
    assign in2970_1 = {pp87[26]};
    assign in2970_2 = {pp88[25]};
    Full_Adder FA_2970(s2970, c2970, in2970_1, in2970_2, pp86[27]);
    wire[0:0] s2971, in2971_1, in2971_2;
    wire c2971;
    assign in2971_1 = {pp90[23]};
    assign in2971_2 = {pp91[22]};
    Full_Adder FA_2971(s2971, c2971, in2971_1, in2971_2, pp89[24]);
    wire[0:0] s2972, in2972_1, in2972_2;
    wire c2972;
    assign in2972_1 = {pp93[20]};
    assign in2972_2 = {pp94[19]};
    Full_Adder FA_2972(s2972, c2972, in2972_1, in2972_2, pp92[21]);
    wire[0:0] s2973, in2973_1, in2973_2;
    wire c2973;
    assign in2973_1 = {pp96[17]};
    assign in2973_2 = {pp97[16]};
    Full_Adder FA_2973(s2973, c2973, in2973_1, in2973_2, pp95[18]);
    wire[0:0] s2974, in2974_1, in2974_2;
    wire c2974;
    assign in2974_1 = {pp99[14]};
    assign in2974_2 = {pp100[13]};
    Full_Adder FA_2974(s2974, c2974, in2974_1, in2974_2, pp98[15]);
    wire[0:0] s2975, in2975_1, in2975_2;
    wire c2975;
    assign in2975_1 = {pp102[11]};
    assign in2975_2 = {pp103[10]};
    Full_Adder FA_2975(s2975, c2975, in2975_1, in2975_2, pp101[12]);
    wire[0:0] s2976, in2976_1, in2976_2;
    wire c2976;
    assign in2976_1 = {pp105[8]};
    assign in2976_2 = {pp106[7]};
    Full_Adder FA_2976(s2976, c2976, in2976_1, in2976_2, pp104[9]);
    wire[0:0] s2977, in2977_1, in2977_2;
    wire c2977;
    assign in2977_1 = {pp108[5]};
    assign in2977_2 = {pp109[4]};
    Full_Adder FA_2977(s2977, c2977, in2977_1, in2977_2, pp107[6]);
    wire[0:0] s2978, in2978_1, in2978_2;
    wire c2978;
    assign in2978_1 = {pp111[2]};
    assign in2978_2 = {pp112[1]};
    Full_Adder FA_2978(s2978, c2978, in2978_1, in2978_2, pp110[3]);
    wire[0:0] s2979, in2979_1, in2979_2;
    wire c2979;
    assign in2979_1 = {c352};
    assign in2979_2 = {c353};
    Full_Adder FA_2979(s2979, c2979, in2979_1, in2979_2, pp113[0]);
    wire[0:0] s2980, in2980_1, in2980_2;
    wire c2980;
    assign in2980_1 = {c355};
    assign in2980_2 = {c356};
    Full_Adder FA_2980(s2980, c2980, in2980_1, in2980_2, c354);
    wire[0:0] s2981, in2981_1, in2981_2;
    wire c2981;
    assign in2981_1 = {c358};
    assign in2981_2 = {c359};
    Full_Adder FA_2981(s2981, c2981, in2981_1, in2981_2, c357);
    wire[0:0] s2982, in2982_1, in2982_2;
    wire c2982;
    assign in2982_1 = {c361};
    assign in2982_2 = {c362};
    Full_Adder FA_2982(s2982, c2982, in2982_1, in2982_2, c360);
    wire[0:0] s2983, in2983_1, in2983_2;
    wire c2983;
    assign in2983_1 = {c364};
    assign in2983_2 = {c365};
    Full_Adder FA_2983(s2983, c2983, in2983_1, in2983_2, c363);
    wire[0:0] s2984, in2984_1, in2984_2;
    wire c2984;
    assign in2984_1 = {c367};
    assign in2984_2 = {c368};
    Full_Adder FA_2984(s2984, c2984, in2984_1, in2984_2, c366);
    wire[0:0] s2985, in2985_1, in2985_2;
    wire c2985;
    assign in2985_1 = {c370};
    assign in2985_2 = {c371};
    Full_Adder FA_2985(s2985, c2985, in2985_1, in2985_2, c369);
    wire[0:0] s2986, in2986_1, in2986_2;
    wire c2986;
    assign in2986_1 = {c373};
    assign in2986_2 = {c374};
    Full_Adder FA_2986(s2986, c2986, in2986_1, in2986_2, c372);
    wire[0:0] s2987, in2987_1, in2987_2;
    wire c2987;
    assign in2987_1 = {c376};
    assign in2987_2 = {c377};
    Full_Adder FA_2987(s2987, c2987, in2987_1, in2987_2, c375);
    wire[0:0] s2988, in2988_1, in2988_2;
    wire c2988;
    assign in2988_1 = {s379[0]};
    assign in2988_2 = {s380[0]};
    Full_Adder FA_2988(s2988, c2988, in2988_1, in2988_2, c378);
    wire[0:0] s2989, in2989_1, in2989_2;
    wire c2989;
    assign in2989_1 = {s382[0]};
    assign in2989_2 = {s383[0]};
    Full_Adder FA_2989(s2989, c2989, in2989_1, in2989_2, s381[0]);
    wire[0:0] s2990, in2990_1, in2990_2;
    wire c2990;
    assign in2990_1 = {s385[0]};
    assign in2990_2 = {s386[0]};
    Full_Adder FA_2990(s2990, c2990, in2990_1, in2990_2, s384[0]);
    wire[0:0] s2991, in2991_1, in2991_2;
    wire c2991;
    assign in2991_1 = {s388[0]};
    assign in2991_2 = {s389[0]};
    Full_Adder FA_2991(s2991, c2991, in2991_1, in2991_2, s387[0]);
    wire[0:0] s2992, in2992_1, in2992_2;
    wire c2992;
    assign in2992_1 = {s391[0]};
    assign in2992_2 = {s392[0]};
    Full_Adder FA_2992(s2992, c2992, in2992_1, in2992_2, s390[0]);
    wire[0:0] s2993, in2993_1, in2993_2;
    wire c2993;
    assign in2993_1 = {s394[0]};
    assign in2993_2 = {s395[0]};
    Full_Adder FA_2993(s2993, c2993, in2993_1, in2993_2, s393[0]);
    wire[0:0] s2994, in2994_1, in2994_2;
    wire c2994;
    assign in2994_1 = {s397[0]};
    assign in2994_2 = {s398[0]};
    Full_Adder FA_2994(s2994, c2994, in2994_1, in2994_2, s396[0]);
    wire[0:0] s2995, in2995_1, in2995_2;
    wire c2995;
    assign in2995_1 = {s400[0]};
    assign in2995_2 = {s401[0]};
    Full_Adder FA_2995(s2995, c2995, in2995_1, in2995_2, s399[0]);
    wire[0:0] s2996, in2996_1, in2996_2;
    wire c2996;
    assign in2996_1 = {s403[0]};
    assign in2996_2 = {s404[0]};
    Full_Adder FA_2996(s2996, c2996, in2996_1, in2996_2, s402[0]);
    wire[0:0] s2997, in2997_1, in2997_2;
    wire c2997;
    assign in2997_1 = {pp87[27]};
    assign in2997_2 = {pp88[26]};
    Full_Adder FA_2997(s2997, c2997, in2997_1, in2997_2, pp86[28]);
    wire[0:0] s2998, in2998_1, in2998_2;
    wire c2998;
    assign in2998_1 = {pp90[24]};
    assign in2998_2 = {pp91[23]};
    Full_Adder FA_2998(s2998, c2998, in2998_1, in2998_2, pp89[25]);
    wire[0:0] s2999, in2999_1, in2999_2;
    wire c2999;
    assign in2999_1 = {pp93[21]};
    assign in2999_2 = {pp94[20]};
    Full_Adder FA_2999(s2999, c2999, in2999_1, in2999_2, pp92[22]);
    wire[0:0] s3000, in3000_1, in3000_2;
    wire c3000;
    assign in3000_1 = {pp96[18]};
    assign in3000_2 = {pp97[17]};
    Full_Adder FA_3000(s3000, c3000, in3000_1, in3000_2, pp95[19]);
    wire[0:0] s3001, in3001_1, in3001_2;
    wire c3001;
    assign in3001_1 = {pp99[15]};
    assign in3001_2 = {pp100[14]};
    Full_Adder FA_3001(s3001, c3001, in3001_1, in3001_2, pp98[16]);
    wire[0:0] s3002, in3002_1, in3002_2;
    wire c3002;
    assign in3002_1 = {pp102[12]};
    assign in3002_2 = {pp103[11]};
    Full_Adder FA_3002(s3002, c3002, in3002_1, in3002_2, pp101[13]);
    wire[0:0] s3003, in3003_1, in3003_2;
    wire c3003;
    assign in3003_1 = {pp105[9]};
    assign in3003_2 = {pp106[8]};
    Full_Adder FA_3003(s3003, c3003, in3003_1, in3003_2, pp104[10]);
    wire[0:0] s3004, in3004_1, in3004_2;
    wire c3004;
    assign in3004_1 = {pp108[6]};
    assign in3004_2 = {pp109[5]};
    Full_Adder FA_3004(s3004, c3004, in3004_1, in3004_2, pp107[7]);
    wire[0:0] s3005, in3005_1, in3005_2;
    wire c3005;
    assign in3005_1 = {pp111[3]};
    assign in3005_2 = {pp112[2]};
    Full_Adder FA_3005(s3005, c3005, in3005_1, in3005_2, pp110[4]);
    wire[0:0] s3006, in3006_1, in3006_2;
    wire c3006;
    assign in3006_1 = {pp114[0]};
    assign in3006_2 = {c379};
    Full_Adder FA_3006(s3006, c3006, in3006_1, in3006_2, pp113[1]);
    wire[0:0] s3007, in3007_1, in3007_2;
    wire c3007;
    assign in3007_1 = {c381};
    assign in3007_2 = {c382};
    Full_Adder FA_3007(s3007, c3007, in3007_1, in3007_2, c380);
    wire[0:0] s3008, in3008_1, in3008_2;
    wire c3008;
    assign in3008_1 = {c384};
    assign in3008_2 = {c385};
    Full_Adder FA_3008(s3008, c3008, in3008_1, in3008_2, c383);
    wire[0:0] s3009, in3009_1, in3009_2;
    wire c3009;
    assign in3009_1 = {c387};
    assign in3009_2 = {c388};
    Full_Adder FA_3009(s3009, c3009, in3009_1, in3009_2, c386);
    wire[0:0] s3010, in3010_1, in3010_2;
    wire c3010;
    assign in3010_1 = {c390};
    assign in3010_2 = {c391};
    Full_Adder FA_3010(s3010, c3010, in3010_1, in3010_2, c389);
    wire[0:0] s3011, in3011_1, in3011_2;
    wire c3011;
    assign in3011_1 = {c393};
    assign in3011_2 = {c394};
    Full_Adder FA_3011(s3011, c3011, in3011_1, in3011_2, c392);
    wire[0:0] s3012, in3012_1, in3012_2;
    wire c3012;
    assign in3012_1 = {c396};
    assign in3012_2 = {c397};
    Full_Adder FA_3012(s3012, c3012, in3012_1, in3012_2, c395);
    wire[0:0] s3013, in3013_1, in3013_2;
    wire c3013;
    assign in3013_1 = {c399};
    assign in3013_2 = {c400};
    Full_Adder FA_3013(s3013, c3013, in3013_1, in3013_2, c398);
    wire[0:0] s3014, in3014_1, in3014_2;
    wire c3014;
    assign in3014_1 = {c402};
    assign in3014_2 = {c403};
    Full_Adder FA_3014(s3014, c3014, in3014_1, in3014_2, c401);
    wire[0:0] s3015, in3015_1, in3015_2;
    wire c3015;
    assign in3015_1 = {c405};
    assign in3015_2 = {c406};
    Full_Adder FA_3015(s3015, c3015, in3015_1, in3015_2, c404);
    wire[0:0] s3016, in3016_1, in3016_2;
    wire c3016;
    assign in3016_1 = {s408[0]};
    assign in3016_2 = {s409[0]};
    Full_Adder FA_3016(s3016, c3016, in3016_1, in3016_2, s407[0]);
    wire[0:0] s3017, in3017_1, in3017_2;
    wire c3017;
    assign in3017_1 = {s411[0]};
    assign in3017_2 = {s412[0]};
    Full_Adder FA_3017(s3017, c3017, in3017_1, in3017_2, s410[0]);
    wire[0:0] s3018, in3018_1, in3018_2;
    wire c3018;
    assign in3018_1 = {s414[0]};
    assign in3018_2 = {s415[0]};
    Full_Adder FA_3018(s3018, c3018, in3018_1, in3018_2, s413[0]);
    wire[0:0] s3019, in3019_1, in3019_2;
    wire c3019;
    assign in3019_1 = {s417[0]};
    assign in3019_2 = {s418[0]};
    Full_Adder FA_3019(s3019, c3019, in3019_1, in3019_2, s416[0]);
    wire[0:0] s3020, in3020_1, in3020_2;
    wire c3020;
    assign in3020_1 = {s420[0]};
    assign in3020_2 = {s421[0]};
    Full_Adder FA_3020(s3020, c3020, in3020_1, in3020_2, s419[0]);
    wire[0:0] s3021, in3021_1, in3021_2;
    wire c3021;
    assign in3021_1 = {s423[0]};
    assign in3021_2 = {s424[0]};
    Full_Adder FA_3021(s3021, c3021, in3021_1, in3021_2, s422[0]);
    wire[0:0] s3022, in3022_1, in3022_2;
    wire c3022;
    assign in3022_1 = {s426[0]};
    assign in3022_2 = {s427[0]};
    Full_Adder FA_3022(s3022, c3022, in3022_1, in3022_2, s425[0]);
    wire[0:0] s3023, in3023_1, in3023_2;
    wire c3023;
    assign in3023_1 = {s429[0]};
    assign in3023_2 = {s430[0]};
    Full_Adder FA_3023(s3023, c3023, in3023_1, in3023_2, s428[0]);
    wire[0:0] s3024, in3024_1, in3024_2;
    wire c3024;
    assign in3024_1 = {s432[0]};
    assign in3024_2 = {s433[0]};
    Full_Adder FA_3024(s3024, c3024, in3024_1, in3024_2, s431[0]);
    wire[0:0] s3025, in3025_1, in3025_2;
    wire c3025;
    assign in3025_1 = {pp90[25]};
    assign in3025_2 = {pp91[24]};
    Full_Adder FA_3025(s3025, c3025, in3025_1, in3025_2, pp89[26]);
    wire[0:0] s3026, in3026_1, in3026_2;
    wire c3026;
    assign in3026_1 = {pp93[22]};
    assign in3026_2 = {pp94[21]};
    Full_Adder FA_3026(s3026, c3026, in3026_1, in3026_2, pp92[23]);
    wire[0:0] s3027, in3027_1, in3027_2;
    wire c3027;
    assign in3027_1 = {pp96[19]};
    assign in3027_2 = {pp97[18]};
    Full_Adder FA_3027(s3027, c3027, in3027_1, in3027_2, pp95[20]);
    wire[0:0] s3028, in3028_1, in3028_2;
    wire c3028;
    assign in3028_1 = {pp99[16]};
    assign in3028_2 = {pp100[15]};
    Full_Adder FA_3028(s3028, c3028, in3028_1, in3028_2, pp98[17]);
    wire[0:0] s3029, in3029_1, in3029_2;
    wire c3029;
    assign in3029_1 = {pp102[13]};
    assign in3029_2 = {pp103[12]};
    Full_Adder FA_3029(s3029, c3029, in3029_1, in3029_2, pp101[14]);
    wire[0:0] s3030, in3030_1, in3030_2;
    wire c3030;
    assign in3030_1 = {pp105[10]};
    assign in3030_2 = {pp106[9]};
    Full_Adder FA_3030(s3030, c3030, in3030_1, in3030_2, pp104[11]);
    wire[0:0] s3031, in3031_1, in3031_2;
    wire c3031;
    assign in3031_1 = {pp108[7]};
    assign in3031_2 = {pp109[6]};
    Full_Adder FA_3031(s3031, c3031, in3031_1, in3031_2, pp107[8]);
    wire[0:0] s3032, in3032_1, in3032_2;
    wire c3032;
    assign in3032_1 = {pp111[4]};
    assign in3032_2 = {pp112[3]};
    Full_Adder FA_3032(s3032, c3032, in3032_1, in3032_2, pp110[5]);
    wire[0:0] s3033, in3033_1, in3033_2;
    wire c3033;
    assign in3033_1 = {pp114[1]};
    assign in3033_2 = {pp115[0]};
    Full_Adder FA_3033(s3033, c3033, in3033_1, in3033_2, pp113[2]);
    wire[0:0] s3034, in3034_1, in3034_2;
    wire c3034;
    assign in3034_1 = {c408};
    assign in3034_2 = {c409};
    Full_Adder FA_3034(s3034, c3034, in3034_1, in3034_2, c407);
    wire[0:0] s3035, in3035_1, in3035_2;
    wire c3035;
    assign in3035_1 = {c411};
    assign in3035_2 = {c412};
    Full_Adder FA_3035(s3035, c3035, in3035_1, in3035_2, c410);
    wire[0:0] s3036, in3036_1, in3036_2;
    wire c3036;
    assign in3036_1 = {c414};
    assign in3036_2 = {c415};
    Full_Adder FA_3036(s3036, c3036, in3036_1, in3036_2, c413);
    wire[0:0] s3037, in3037_1, in3037_2;
    wire c3037;
    assign in3037_1 = {c417};
    assign in3037_2 = {c418};
    Full_Adder FA_3037(s3037, c3037, in3037_1, in3037_2, c416);
    wire[0:0] s3038, in3038_1, in3038_2;
    wire c3038;
    assign in3038_1 = {c420};
    assign in3038_2 = {c421};
    Full_Adder FA_3038(s3038, c3038, in3038_1, in3038_2, c419);
    wire[0:0] s3039, in3039_1, in3039_2;
    wire c3039;
    assign in3039_1 = {c423};
    assign in3039_2 = {c424};
    Full_Adder FA_3039(s3039, c3039, in3039_1, in3039_2, c422);
    wire[0:0] s3040, in3040_1, in3040_2;
    wire c3040;
    assign in3040_1 = {c426};
    assign in3040_2 = {c427};
    Full_Adder FA_3040(s3040, c3040, in3040_1, in3040_2, c425);
    wire[0:0] s3041, in3041_1, in3041_2;
    wire c3041;
    assign in3041_1 = {c429};
    assign in3041_2 = {c430};
    Full_Adder FA_3041(s3041, c3041, in3041_1, in3041_2, c428);
    wire[0:0] s3042, in3042_1, in3042_2;
    wire c3042;
    assign in3042_1 = {c432};
    assign in3042_2 = {c433};
    Full_Adder FA_3042(s3042, c3042, in3042_1, in3042_2, c431);
    wire[0:0] s3043, in3043_1, in3043_2;
    wire c3043;
    assign in3043_1 = {c435};
    assign in3043_2 = {s436[0]};
    Full_Adder FA_3043(s3043, c3043, in3043_1, in3043_2, c434);
    wire[0:0] s3044, in3044_1, in3044_2;
    wire c3044;
    assign in3044_1 = {s438[0]};
    assign in3044_2 = {s439[0]};
    Full_Adder FA_3044(s3044, c3044, in3044_1, in3044_2, s437[0]);
    wire[0:0] s3045, in3045_1, in3045_2;
    wire c3045;
    assign in3045_1 = {s441[0]};
    assign in3045_2 = {s442[0]};
    Full_Adder FA_3045(s3045, c3045, in3045_1, in3045_2, s440[0]);
    wire[0:0] s3046, in3046_1, in3046_2;
    wire c3046;
    assign in3046_1 = {s444[0]};
    assign in3046_2 = {s445[0]};
    Full_Adder FA_3046(s3046, c3046, in3046_1, in3046_2, s443[0]);
    wire[0:0] s3047, in3047_1, in3047_2;
    wire c3047;
    assign in3047_1 = {s447[0]};
    assign in3047_2 = {s448[0]};
    Full_Adder FA_3047(s3047, c3047, in3047_1, in3047_2, s446[0]);
    wire[0:0] s3048, in3048_1, in3048_2;
    wire c3048;
    assign in3048_1 = {s450[0]};
    assign in3048_2 = {s451[0]};
    Full_Adder FA_3048(s3048, c3048, in3048_1, in3048_2, s449[0]);
    wire[0:0] s3049, in3049_1, in3049_2;
    wire c3049;
    assign in3049_1 = {s453[0]};
    assign in3049_2 = {s454[0]};
    Full_Adder FA_3049(s3049, c3049, in3049_1, in3049_2, s452[0]);
    wire[0:0] s3050, in3050_1, in3050_2;
    wire c3050;
    assign in3050_1 = {s456[0]};
    assign in3050_2 = {s457[0]};
    Full_Adder FA_3050(s3050, c3050, in3050_1, in3050_2, s455[0]);
    wire[0:0] s3051, in3051_1, in3051_2;
    wire c3051;
    assign in3051_1 = {s459[0]};
    assign in3051_2 = {s460[0]};
    Full_Adder FA_3051(s3051, c3051, in3051_1, in3051_2, s458[0]);
    wire[0:0] s3052, in3052_1, in3052_2;
    wire c3052;
    assign in3052_1 = {s462[0]};
    assign in3052_2 = {s463[0]};
    Full_Adder FA_3052(s3052, c3052, in3052_1, in3052_2, s461[0]);
    wire[0:0] s3053, in3053_1, in3053_2;
    wire c3053;
    assign in3053_1 = {pp93[23]};
    assign in3053_2 = {pp94[22]};
    Full_Adder FA_3053(s3053, c3053, in3053_1, in3053_2, pp92[24]);
    wire[0:0] s3054, in3054_1, in3054_2;
    wire c3054;
    assign in3054_1 = {pp96[20]};
    assign in3054_2 = {pp97[19]};
    Full_Adder FA_3054(s3054, c3054, in3054_1, in3054_2, pp95[21]);
    wire[0:0] s3055, in3055_1, in3055_2;
    wire c3055;
    assign in3055_1 = {pp99[17]};
    assign in3055_2 = {pp100[16]};
    Full_Adder FA_3055(s3055, c3055, in3055_1, in3055_2, pp98[18]);
    wire[0:0] s3056, in3056_1, in3056_2;
    wire c3056;
    assign in3056_1 = {pp102[14]};
    assign in3056_2 = {pp103[13]};
    Full_Adder FA_3056(s3056, c3056, in3056_1, in3056_2, pp101[15]);
    wire[0:0] s3057, in3057_1, in3057_2;
    wire c3057;
    assign in3057_1 = {pp105[11]};
    assign in3057_2 = {pp106[10]};
    Full_Adder FA_3057(s3057, c3057, in3057_1, in3057_2, pp104[12]);
    wire[0:0] s3058, in3058_1, in3058_2;
    wire c3058;
    assign in3058_1 = {pp108[8]};
    assign in3058_2 = {pp109[7]};
    Full_Adder FA_3058(s3058, c3058, in3058_1, in3058_2, pp107[9]);
    wire[0:0] s3059, in3059_1, in3059_2;
    wire c3059;
    assign in3059_1 = {pp111[5]};
    assign in3059_2 = {pp112[4]};
    Full_Adder FA_3059(s3059, c3059, in3059_1, in3059_2, pp110[6]);
    wire[0:0] s3060, in3060_1, in3060_2;
    wire c3060;
    assign in3060_1 = {pp114[2]};
    assign in3060_2 = {pp115[1]};
    Full_Adder FA_3060(s3060, c3060, in3060_1, in3060_2, pp113[3]);
    wire[0:0] s3061, in3061_1, in3061_2;
    wire c3061;
    assign in3061_1 = {c436};
    assign in3061_2 = {c437};
    Full_Adder FA_3061(s3061, c3061, in3061_1, in3061_2, pp116[0]);
    wire[0:0] s3062, in3062_1, in3062_2;
    wire c3062;
    assign in3062_1 = {c439};
    assign in3062_2 = {c440};
    Full_Adder FA_3062(s3062, c3062, in3062_1, in3062_2, c438);
    wire[0:0] s3063, in3063_1, in3063_2;
    wire c3063;
    assign in3063_1 = {c442};
    assign in3063_2 = {c443};
    Full_Adder FA_3063(s3063, c3063, in3063_1, in3063_2, c441);
    wire[0:0] s3064, in3064_1, in3064_2;
    wire c3064;
    assign in3064_1 = {c445};
    assign in3064_2 = {c446};
    Full_Adder FA_3064(s3064, c3064, in3064_1, in3064_2, c444);
    wire[0:0] s3065, in3065_1, in3065_2;
    wire c3065;
    assign in3065_1 = {c448};
    assign in3065_2 = {c449};
    Full_Adder FA_3065(s3065, c3065, in3065_1, in3065_2, c447);
    wire[0:0] s3066, in3066_1, in3066_2;
    wire c3066;
    assign in3066_1 = {c451};
    assign in3066_2 = {c452};
    Full_Adder FA_3066(s3066, c3066, in3066_1, in3066_2, c450);
    wire[0:0] s3067, in3067_1, in3067_2;
    wire c3067;
    assign in3067_1 = {c454};
    assign in3067_2 = {c455};
    Full_Adder FA_3067(s3067, c3067, in3067_1, in3067_2, c453);
    wire[0:0] s3068, in3068_1, in3068_2;
    wire c3068;
    assign in3068_1 = {c457};
    assign in3068_2 = {c458};
    Full_Adder FA_3068(s3068, c3068, in3068_1, in3068_2, c456);
    wire[0:0] s3069, in3069_1, in3069_2;
    wire c3069;
    assign in3069_1 = {c460};
    assign in3069_2 = {c461};
    Full_Adder FA_3069(s3069, c3069, in3069_1, in3069_2, c459);
    wire[0:0] s3070, in3070_1, in3070_2;
    wire c3070;
    assign in3070_1 = {c463};
    assign in3070_2 = {c464};
    Full_Adder FA_3070(s3070, c3070, in3070_1, in3070_2, c462);
    wire[0:0] s3071, in3071_1, in3071_2;
    wire c3071;
    assign in3071_1 = {s466[0]};
    assign in3071_2 = {s467[0]};
    Full_Adder FA_3071(s3071, c3071, in3071_1, in3071_2, c465);
    wire[0:0] s3072, in3072_1, in3072_2;
    wire c3072;
    assign in3072_1 = {s469[0]};
    assign in3072_2 = {s470[0]};
    Full_Adder FA_3072(s3072, c3072, in3072_1, in3072_2, s468[0]);
    wire[0:0] s3073, in3073_1, in3073_2;
    wire c3073;
    assign in3073_1 = {s472[0]};
    assign in3073_2 = {s473[0]};
    Full_Adder FA_3073(s3073, c3073, in3073_1, in3073_2, s471[0]);
    wire[0:0] s3074, in3074_1, in3074_2;
    wire c3074;
    assign in3074_1 = {s475[0]};
    assign in3074_2 = {s476[0]};
    Full_Adder FA_3074(s3074, c3074, in3074_1, in3074_2, s474[0]);
    wire[0:0] s3075, in3075_1, in3075_2;
    wire c3075;
    assign in3075_1 = {s478[0]};
    assign in3075_2 = {s479[0]};
    Full_Adder FA_3075(s3075, c3075, in3075_1, in3075_2, s477[0]);
    wire[0:0] s3076, in3076_1, in3076_2;
    wire c3076;
    assign in3076_1 = {s481[0]};
    assign in3076_2 = {s482[0]};
    Full_Adder FA_3076(s3076, c3076, in3076_1, in3076_2, s480[0]);
    wire[0:0] s3077, in3077_1, in3077_2;
    wire c3077;
    assign in3077_1 = {s484[0]};
    assign in3077_2 = {s485[0]};
    Full_Adder FA_3077(s3077, c3077, in3077_1, in3077_2, s483[0]);
    wire[0:0] s3078, in3078_1, in3078_2;
    wire c3078;
    assign in3078_1 = {s487[0]};
    assign in3078_2 = {s488[0]};
    Full_Adder FA_3078(s3078, c3078, in3078_1, in3078_2, s486[0]);
    wire[0:0] s3079, in3079_1, in3079_2;
    wire c3079;
    assign in3079_1 = {s490[0]};
    assign in3079_2 = {s491[0]};
    Full_Adder FA_3079(s3079, c3079, in3079_1, in3079_2, s489[0]);
    wire[0:0] s3080, in3080_1, in3080_2;
    wire c3080;
    assign in3080_1 = {s493[0]};
    assign in3080_2 = {s494[0]};
    Full_Adder FA_3080(s3080, c3080, in3080_1, in3080_2, s492[0]);
    wire[0:0] s3081, in3081_1, in3081_2;
    wire c3081;
    assign in3081_1 = {pp96[21]};
    assign in3081_2 = {pp97[20]};
    Full_Adder FA_3081(s3081, c3081, in3081_1, in3081_2, pp95[22]);
    wire[0:0] s3082, in3082_1, in3082_2;
    wire c3082;
    assign in3082_1 = {pp99[18]};
    assign in3082_2 = {pp100[17]};
    Full_Adder FA_3082(s3082, c3082, in3082_1, in3082_2, pp98[19]);
    wire[0:0] s3083, in3083_1, in3083_2;
    wire c3083;
    assign in3083_1 = {pp102[15]};
    assign in3083_2 = {pp103[14]};
    Full_Adder FA_3083(s3083, c3083, in3083_1, in3083_2, pp101[16]);
    wire[0:0] s3084, in3084_1, in3084_2;
    wire c3084;
    assign in3084_1 = {pp105[12]};
    assign in3084_2 = {pp106[11]};
    Full_Adder FA_3084(s3084, c3084, in3084_1, in3084_2, pp104[13]);
    wire[0:0] s3085, in3085_1, in3085_2;
    wire c3085;
    assign in3085_1 = {pp108[9]};
    assign in3085_2 = {pp109[8]};
    Full_Adder FA_3085(s3085, c3085, in3085_1, in3085_2, pp107[10]);
    wire[0:0] s3086, in3086_1, in3086_2;
    wire c3086;
    assign in3086_1 = {pp111[6]};
    assign in3086_2 = {pp112[5]};
    Full_Adder FA_3086(s3086, c3086, in3086_1, in3086_2, pp110[7]);
    wire[0:0] s3087, in3087_1, in3087_2;
    wire c3087;
    assign in3087_1 = {pp114[3]};
    assign in3087_2 = {pp115[2]};
    Full_Adder FA_3087(s3087, c3087, in3087_1, in3087_2, pp113[4]);
    wire[0:0] s3088, in3088_1, in3088_2;
    wire c3088;
    assign in3088_1 = {pp117[0]};
    assign in3088_2 = {c466};
    Full_Adder FA_3088(s3088, c3088, in3088_1, in3088_2, pp116[1]);
    wire[0:0] s3089, in3089_1, in3089_2;
    wire c3089;
    assign in3089_1 = {c468};
    assign in3089_2 = {c469};
    Full_Adder FA_3089(s3089, c3089, in3089_1, in3089_2, c467);
    wire[0:0] s3090, in3090_1, in3090_2;
    wire c3090;
    assign in3090_1 = {c471};
    assign in3090_2 = {c472};
    Full_Adder FA_3090(s3090, c3090, in3090_1, in3090_2, c470);
    wire[0:0] s3091, in3091_1, in3091_2;
    wire c3091;
    assign in3091_1 = {c474};
    assign in3091_2 = {c475};
    Full_Adder FA_3091(s3091, c3091, in3091_1, in3091_2, c473);
    wire[0:0] s3092, in3092_1, in3092_2;
    wire c3092;
    assign in3092_1 = {c477};
    assign in3092_2 = {c478};
    Full_Adder FA_3092(s3092, c3092, in3092_1, in3092_2, c476);
    wire[0:0] s3093, in3093_1, in3093_2;
    wire c3093;
    assign in3093_1 = {c480};
    assign in3093_2 = {c481};
    Full_Adder FA_3093(s3093, c3093, in3093_1, in3093_2, c479);
    wire[0:0] s3094, in3094_1, in3094_2;
    wire c3094;
    assign in3094_1 = {c483};
    assign in3094_2 = {c484};
    Full_Adder FA_3094(s3094, c3094, in3094_1, in3094_2, c482);
    wire[0:0] s3095, in3095_1, in3095_2;
    wire c3095;
    assign in3095_1 = {c486};
    assign in3095_2 = {c487};
    Full_Adder FA_3095(s3095, c3095, in3095_1, in3095_2, c485);
    wire[0:0] s3096, in3096_1, in3096_2;
    wire c3096;
    assign in3096_1 = {c489};
    assign in3096_2 = {c490};
    Full_Adder FA_3096(s3096, c3096, in3096_1, in3096_2, c488);
    wire[0:0] s3097, in3097_1, in3097_2;
    wire c3097;
    assign in3097_1 = {c492};
    assign in3097_2 = {c493};
    Full_Adder FA_3097(s3097, c3097, in3097_1, in3097_2, c491);
    wire[0:0] s3098, in3098_1, in3098_2;
    wire c3098;
    assign in3098_1 = {c495};
    assign in3098_2 = {c496};
    Full_Adder FA_3098(s3098, c3098, in3098_1, in3098_2, c494);
    wire[0:0] s3099, in3099_1, in3099_2;
    wire c3099;
    assign in3099_1 = {s498[0]};
    assign in3099_2 = {s499[0]};
    Full_Adder FA_3099(s3099, c3099, in3099_1, in3099_2, s497[0]);
    wire[0:0] s3100, in3100_1, in3100_2;
    wire c3100;
    assign in3100_1 = {s501[0]};
    assign in3100_2 = {s502[0]};
    Full_Adder FA_3100(s3100, c3100, in3100_1, in3100_2, s500[0]);
    wire[0:0] s3101, in3101_1, in3101_2;
    wire c3101;
    assign in3101_1 = {s504[0]};
    assign in3101_2 = {s505[0]};
    Full_Adder FA_3101(s3101, c3101, in3101_1, in3101_2, s503[0]);
    wire[0:0] s3102, in3102_1, in3102_2;
    wire c3102;
    assign in3102_1 = {s507[0]};
    assign in3102_2 = {s508[0]};
    Full_Adder FA_3102(s3102, c3102, in3102_1, in3102_2, s506[0]);
    wire[0:0] s3103, in3103_1, in3103_2;
    wire c3103;
    assign in3103_1 = {s510[0]};
    assign in3103_2 = {s511[0]};
    Full_Adder FA_3103(s3103, c3103, in3103_1, in3103_2, s509[0]);
    wire[0:0] s3104, in3104_1, in3104_2;
    wire c3104;
    assign in3104_1 = {s513[0]};
    assign in3104_2 = {s514[0]};
    Full_Adder FA_3104(s3104, c3104, in3104_1, in3104_2, s512[0]);
    wire[0:0] s3105, in3105_1, in3105_2;
    wire c3105;
    assign in3105_1 = {s516[0]};
    assign in3105_2 = {s517[0]};
    Full_Adder FA_3105(s3105, c3105, in3105_1, in3105_2, s515[0]);
    wire[0:0] s3106, in3106_1, in3106_2;
    wire c3106;
    assign in3106_1 = {s519[0]};
    assign in3106_2 = {s520[0]};
    Full_Adder FA_3106(s3106, c3106, in3106_1, in3106_2, s518[0]);
    wire[0:0] s3107, in3107_1, in3107_2;
    wire c3107;
    assign in3107_1 = {s522[0]};
    assign in3107_2 = {s523[0]};
    Full_Adder FA_3107(s3107, c3107, in3107_1, in3107_2, s521[0]);
    wire[0:0] s3108, in3108_1, in3108_2;
    wire c3108;
    assign in3108_1 = {s525[0]};
    assign in3108_2 = {s526[0]};
    Full_Adder FA_3108(s3108, c3108, in3108_1, in3108_2, s524[0]);
    wire[0:0] s3109, in3109_1, in3109_2;
    wire c3109;
    assign in3109_1 = {pp99[19]};
    assign in3109_2 = {pp100[18]};
    Full_Adder FA_3109(s3109, c3109, in3109_1, in3109_2, pp98[20]);
    wire[0:0] s3110, in3110_1, in3110_2;
    wire c3110;
    assign in3110_1 = {pp102[16]};
    assign in3110_2 = {pp103[15]};
    Full_Adder FA_3110(s3110, c3110, in3110_1, in3110_2, pp101[17]);
    wire[0:0] s3111, in3111_1, in3111_2;
    wire c3111;
    assign in3111_1 = {pp105[13]};
    assign in3111_2 = {pp106[12]};
    Full_Adder FA_3111(s3111, c3111, in3111_1, in3111_2, pp104[14]);
    wire[0:0] s3112, in3112_1, in3112_2;
    wire c3112;
    assign in3112_1 = {pp108[10]};
    assign in3112_2 = {pp109[9]};
    Full_Adder FA_3112(s3112, c3112, in3112_1, in3112_2, pp107[11]);
    wire[0:0] s3113, in3113_1, in3113_2;
    wire c3113;
    assign in3113_1 = {pp111[7]};
    assign in3113_2 = {pp112[6]};
    Full_Adder FA_3113(s3113, c3113, in3113_1, in3113_2, pp110[8]);
    wire[0:0] s3114, in3114_1, in3114_2;
    wire c3114;
    assign in3114_1 = {pp114[4]};
    assign in3114_2 = {pp115[3]};
    Full_Adder FA_3114(s3114, c3114, in3114_1, in3114_2, pp113[5]);
    wire[0:0] s3115, in3115_1, in3115_2;
    wire c3115;
    assign in3115_1 = {pp117[1]};
    assign in3115_2 = {pp118[0]};
    Full_Adder FA_3115(s3115, c3115, in3115_1, in3115_2, pp116[2]);
    wire[0:0] s3116, in3116_1, in3116_2;
    wire c3116;
    assign in3116_1 = {c498};
    assign in3116_2 = {c499};
    Full_Adder FA_3116(s3116, c3116, in3116_1, in3116_2, c497);
    wire[0:0] s3117, in3117_1, in3117_2;
    wire c3117;
    assign in3117_1 = {c501};
    assign in3117_2 = {c502};
    Full_Adder FA_3117(s3117, c3117, in3117_1, in3117_2, c500);
    wire[0:0] s3118, in3118_1, in3118_2;
    wire c3118;
    assign in3118_1 = {c504};
    assign in3118_2 = {c505};
    Full_Adder FA_3118(s3118, c3118, in3118_1, in3118_2, c503);
    wire[0:0] s3119, in3119_1, in3119_2;
    wire c3119;
    assign in3119_1 = {c507};
    assign in3119_2 = {c508};
    Full_Adder FA_3119(s3119, c3119, in3119_1, in3119_2, c506);
    wire[0:0] s3120, in3120_1, in3120_2;
    wire c3120;
    assign in3120_1 = {c510};
    assign in3120_2 = {c511};
    Full_Adder FA_3120(s3120, c3120, in3120_1, in3120_2, c509);
    wire[0:0] s3121, in3121_1, in3121_2;
    wire c3121;
    assign in3121_1 = {c513};
    assign in3121_2 = {c514};
    Full_Adder FA_3121(s3121, c3121, in3121_1, in3121_2, c512);
    wire[0:0] s3122, in3122_1, in3122_2;
    wire c3122;
    assign in3122_1 = {c516};
    assign in3122_2 = {c517};
    Full_Adder FA_3122(s3122, c3122, in3122_1, in3122_2, c515);
    wire[0:0] s3123, in3123_1, in3123_2;
    wire c3123;
    assign in3123_1 = {c519};
    assign in3123_2 = {c520};
    Full_Adder FA_3123(s3123, c3123, in3123_1, in3123_2, c518);
    wire[0:0] s3124, in3124_1, in3124_2;
    wire c3124;
    assign in3124_1 = {c522};
    assign in3124_2 = {c523};
    Full_Adder FA_3124(s3124, c3124, in3124_1, in3124_2, c521);
    wire[0:0] s3125, in3125_1, in3125_2;
    wire c3125;
    assign in3125_1 = {c525};
    assign in3125_2 = {c526};
    Full_Adder FA_3125(s3125, c3125, in3125_1, in3125_2, c524);
    wire[0:0] s3126, in3126_1, in3126_2;
    wire c3126;
    assign in3126_1 = {c528};
    assign in3126_2 = {s529[0]};
    Full_Adder FA_3126(s3126, c3126, in3126_1, in3126_2, c527);
    wire[0:0] s3127, in3127_1, in3127_2;
    wire c3127;
    assign in3127_1 = {s531[0]};
    assign in3127_2 = {s532[0]};
    Full_Adder FA_3127(s3127, c3127, in3127_1, in3127_2, s530[0]);
    wire[0:0] s3128, in3128_1, in3128_2;
    wire c3128;
    assign in3128_1 = {s534[0]};
    assign in3128_2 = {s535[0]};
    Full_Adder FA_3128(s3128, c3128, in3128_1, in3128_2, s533[0]);
    wire[0:0] s3129, in3129_1, in3129_2;
    wire c3129;
    assign in3129_1 = {s537[0]};
    assign in3129_2 = {s538[0]};
    Full_Adder FA_3129(s3129, c3129, in3129_1, in3129_2, s536[0]);
    wire[0:0] s3130, in3130_1, in3130_2;
    wire c3130;
    assign in3130_1 = {s540[0]};
    assign in3130_2 = {s541[0]};
    Full_Adder FA_3130(s3130, c3130, in3130_1, in3130_2, s539[0]);
    wire[0:0] s3131, in3131_1, in3131_2;
    wire c3131;
    assign in3131_1 = {s543[0]};
    assign in3131_2 = {s544[0]};
    Full_Adder FA_3131(s3131, c3131, in3131_1, in3131_2, s542[0]);
    wire[0:0] s3132, in3132_1, in3132_2;
    wire c3132;
    assign in3132_1 = {s546[0]};
    assign in3132_2 = {s547[0]};
    Full_Adder FA_3132(s3132, c3132, in3132_1, in3132_2, s545[0]);
    wire[0:0] s3133, in3133_1, in3133_2;
    wire c3133;
    assign in3133_1 = {s549[0]};
    assign in3133_2 = {s550[0]};
    Full_Adder FA_3133(s3133, c3133, in3133_1, in3133_2, s548[0]);
    wire[0:0] s3134, in3134_1, in3134_2;
    wire c3134;
    assign in3134_1 = {s552[0]};
    assign in3134_2 = {s553[0]};
    Full_Adder FA_3134(s3134, c3134, in3134_1, in3134_2, s551[0]);
    wire[0:0] s3135, in3135_1, in3135_2;
    wire c3135;
    assign in3135_1 = {s555[0]};
    assign in3135_2 = {s556[0]};
    Full_Adder FA_3135(s3135, c3135, in3135_1, in3135_2, s554[0]);
    wire[0:0] s3136, in3136_1, in3136_2;
    wire c3136;
    assign in3136_1 = {s558[0]};
    assign in3136_2 = {s559[0]};
    Full_Adder FA_3136(s3136, c3136, in3136_1, in3136_2, s557[0]);
    wire[0:0] s3137, in3137_1, in3137_2;
    wire c3137;
    assign in3137_1 = {pp102[17]};
    assign in3137_2 = {pp103[16]};
    Full_Adder FA_3137(s3137, c3137, in3137_1, in3137_2, pp101[18]);
    wire[0:0] s3138, in3138_1, in3138_2;
    wire c3138;
    assign in3138_1 = {pp105[14]};
    assign in3138_2 = {pp106[13]};
    Full_Adder FA_3138(s3138, c3138, in3138_1, in3138_2, pp104[15]);
    wire[0:0] s3139, in3139_1, in3139_2;
    wire c3139;
    assign in3139_1 = {pp108[11]};
    assign in3139_2 = {pp109[10]};
    Full_Adder FA_3139(s3139, c3139, in3139_1, in3139_2, pp107[12]);
    wire[0:0] s3140, in3140_1, in3140_2;
    wire c3140;
    assign in3140_1 = {pp111[8]};
    assign in3140_2 = {pp112[7]};
    Full_Adder FA_3140(s3140, c3140, in3140_1, in3140_2, pp110[9]);
    wire[0:0] s3141, in3141_1, in3141_2;
    wire c3141;
    assign in3141_1 = {pp114[5]};
    assign in3141_2 = {pp115[4]};
    Full_Adder FA_3141(s3141, c3141, in3141_1, in3141_2, pp113[6]);
    wire[0:0] s3142, in3142_1, in3142_2;
    wire c3142;
    assign in3142_1 = {pp117[2]};
    assign in3142_2 = {pp118[1]};
    Full_Adder FA_3142(s3142, c3142, in3142_1, in3142_2, pp116[3]);
    wire[0:0] s3143, in3143_1, in3143_2;
    wire c3143;
    assign in3143_1 = {c529};
    assign in3143_2 = {c530};
    Full_Adder FA_3143(s3143, c3143, in3143_1, in3143_2, pp119[0]);
    wire[0:0] s3144, in3144_1, in3144_2;
    wire c3144;
    assign in3144_1 = {c532};
    assign in3144_2 = {c533};
    Full_Adder FA_3144(s3144, c3144, in3144_1, in3144_2, c531);
    wire[0:0] s3145, in3145_1, in3145_2;
    wire c3145;
    assign in3145_1 = {c535};
    assign in3145_2 = {c536};
    Full_Adder FA_3145(s3145, c3145, in3145_1, in3145_2, c534);
    wire[0:0] s3146, in3146_1, in3146_2;
    wire c3146;
    assign in3146_1 = {c538};
    assign in3146_2 = {c539};
    Full_Adder FA_3146(s3146, c3146, in3146_1, in3146_2, c537);
    wire[0:0] s3147, in3147_1, in3147_2;
    wire c3147;
    assign in3147_1 = {c541};
    assign in3147_2 = {c542};
    Full_Adder FA_3147(s3147, c3147, in3147_1, in3147_2, c540);
    wire[0:0] s3148, in3148_1, in3148_2;
    wire c3148;
    assign in3148_1 = {c544};
    assign in3148_2 = {c545};
    Full_Adder FA_3148(s3148, c3148, in3148_1, in3148_2, c543);
    wire[0:0] s3149, in3149_1, in3149_2;
    wire c3149;
    assign in3149_1 = {c547};
    assign in3149_2 = {c548};
    Full_Adder FA_3149(s3149, c3149, in3149_1, in3149_2, c546);
    wire[0:0] s3150, in3150_1, in3150_2;
    wire c3150;
    assign in3150_1 = {c550};
    assign in3150_2 = {c551};
    Full_Adder FA_3150(s3150, c3150, in3150_1, in3150_2, c549);
    wire[0:0] s3151, in3151_1, in3151_2;
    wire c3151;
    assign in3151_1 = {c553};
    assign in3151_2 = {c554};
    Full_Adder FA_3151(s3151, c3151, in3151_1, in3151_2, c552);
    wire[0:0] s3152, in3152_1, in3152_2;
    wire c3152;
    assign in3152_1 = {c556};
    assign in3152_2 = {c557};
    Full_Adder FA_3152(s3152, c3152, in3152_1, in3152_2, c555);
    wire[0:0] s3153, in3153_1, in3153_2;
    wire c3153;
    assign in3153_1 = {c559};
    assign in3153_2 = {c560};
    Full_Adder FA_3153(s3153, c3153, in3153_1, in3153_2, c558);
    wire[0:0] s3154, in3154_1, in3154_2;
    wire c3154;
    assign in3154_1 = {s562[0]};
    assign in3154_2 = {s563[0]};
    Full_Adder FA_3154(s3154, c3154, in3154_1, in3154_2, c561);
    wire[0:0] s3155, in3155_1, in3155_2;
    wire c3155;
    assign in3155_1 = {s565[0]};
    assign in3155_2 = {s566[0]};
    Full_Adder FA_3155(s3155, c3155, in3155_1, in3155_2, s564[0]);
    wire[0:0] s3156, in3156_1, in3156_2;
    wire c3156;
    assign in3156_1 = {s568[0]};
    assign in3156_2 = {s569[0]};
    Full_Adder FA_3156(s3156, c3156, in3156_1, in3156_2, s567[0]);
    wire[0:0] s3157, in3157_1, in3157_2;
    wire c3157;
    assign in3157_1 = {s571[0]};
    assign in3157_2 = {s572[0]};
    Full_Adder FA_3157(s3157, c3157, in3157_1, in3157_2, s570[0]);
    wire[0:0] s3158, in3158_1, in3158_2;
    wire c3158;
    assign in3158_1 = {s574[0]};
    assign in3158_2 = {s575[0]};
    Full_Adder FA_3158(s3158, c3158, in3158_1, in3158_2, s573[0]);
    wire[0:0] s3159, in3159_1, in3159_2;
    wire c3159;
    assign in3159_1 = {s577[0]};
    assign in3159_2 = {s578[0]};
    Full_Adder FA_3159(s3159, c3159, in3159_1, in3159_2, s576[0]);
    wire[0:0] s3160, in3160_1, in3160_2;
    wire c3160;
    assign in3160_1 = {s580[0]};
    assign in3160_2 = {s581[0]};
    Full_Adder FA_3160(s3160, c3160, in3160_1, in3160_2, s579[0]);
    wire[0:0] s3161, in3161_1, in3161_2;
    wire c3161;
    assign in3161_1 = {s583[0]};
    assign in3161_2 = {s584[0]};
    Full_Adder FA_3161(s3161, c3161, in3161_1, in3161_2, s582[0]);
    wire[0:0] s3162, in3162_1, in3162_2;
    wire c3162;
    assign in3162_1 = {s586[0]};
    assign in3162_2 = {s587[0]};
    Full_Adder FA_3162(s3162, c3162, in3162_1, in3162_2, s585[0]);
    wire[0:0] s3163, in3163_1, in3163_2;
    wire c3163;
    assign in3163_1 = {s589[0]};
    assign in3163_2 = {s590[0]};
    Full_Adder FA_3163(s3163, c3163, in3163_1, in3163_2, s588[0]);
    wire[0:0] s3164, in3164_1, in3164_2;
    wire c3164;
    assign in3164_1 = {s592[0]};
    assign in3164_2 = {s593[0]};
    Full_Adder FA_3164(s3164, c3164, in3164_1, in3164_2, s591[0]);
    wire[0:0] s3165, in3165_1, in3165_2;
    wire c3165;
    assign in3165_1 = {pp105[15]};
    assign in3165_2 = {pp106[14]};
    Full_Adder FA_3165(s3165, c3165, in3165_1, in3165_2, pp104[16]);
    wire[0:0] s3166, in3166_1, in3166_2;
    wire c3166;
    assign in3166_1 = {pp108[12]};
    assign in3166_2 = {pp109[11]};
    Full_Adder FA_3166(s3166, c3166, in3166_1, in3166_2, pp107[13]);
    wire[0:0] s3167, in3167_1, in3167_2;
    wire c3167;
    assign in3167_1 = {pp111[9]};
    assign in3167_2 = {pp112[8]};
    Full_Adder FA_3167(s3167, c3167, in3167_1, in3167_2, pp110[10]);
    wire[0:0] s3168, in3168_1, in3168_2;
    wire c3168;
    assign in3168_1 = {pp114[6]};
    assign in3168_2 = {pp115[5]};
    Full_Adder FA_3168(s3168, c3168, in3168_1, in3168_2, pp113[7]);
    wire[0:0] s3169, in3169_1, in3169_2;
    wire c3169;
    assign in3169_1 = {pp117[3]};
    assign in3169_2 = {pp118[2]};
    Full_Adder FA_3169(s3169, c3169, in3169_1, in3169_2, pp116[4]);
    wire[0:0] s3170, in3170_1, in3170_2;
    wire c3170;
    assign in3170_1 = {pp120[0]};
    assign in3170_2 = {c562};
    Full_Adder FA_3170(s3170, c3170, in3170_1, in3170_2, pp119[1]);
    wire[0:0] s3171, in3171_1, in3171_2;
    wire c3171;
    assign in3171_1 = {c564};
    assign in3171_2 = {c565};
    Full_Adder FA_3171(s3171, c3171, in3171_1, in3171_2, c563);
    wire[0:0] s3172, in3172_1, in3172_2;
    wire c3172;
    assign in3172_1 = {c567};
    assign in3172_2 = {c568};
    Full_Adder FA_3172(s3172, c3172, in3172_1, in3172_2, c566);
    wire[0:0] s3173, in3173_1, in3173_2;
    wire c3173;
    assign in3173_1 = {c570};
    assign in3173_2 = {c571};
    Full_Adder FA_3173(s3173, c3173, in3173_1, in3173_2, c569);
    wire[0:0] s3174, in3174_1, in3174_2;
    wire c3174;
    assign in3174_1 = {c573};
    assign in3174_2 = {c574};
    Full_Adder FA_3174(s3174, c3174, in3174_1, in3174_2, c572);
    wire[0:0] s3175, in3175_1, in3175_2;
    wire c3175;
    assign in3175_1 = {c576};
    assign in3175_2 = {c577};
    Full_Adder FA_3175(s3175, c3175, in3175_1, in3175_2, c575);
    wire[0:0] s3176, in3176_1, in3176_2;
    wire c3176;
    assign in3176_1 = {c579};
    assign in3176_2 = {c580};
    Full_Adder FA_3176(s3176, c3176, in3176_1, in3176_2, c578);
    wire[0:0] s3177, in3177_1, in3177_2;
    wire c3177;
    assign in3177_1 = {c582};
    assign in3177_2 = {c583};
    Full_Adder FA_3177(s3177, c3177, in3177_1, in3177_2, c581);
    wire[0:0] s3178, in3178_1, in3178_2;
    wire c3178;
    assign in3178_1 = {c585};
    assign in3178_2 = {c586};
    Full_Adder FA_3178(s3178, c3178, in3178_1, in3178_2, c584);
    wire[0:0] s3179, in3179_1, in3179_2;
    wire c3179;
    assign in3179_1 = {c588};
    assign in3179_2 = {c589};
    Full_Adder FA_3179(s3179, c3179, in3179_1, in3179_2, c587);
    wire[0:0] s3180, in3180_1, in3180_2;
    wire c3180;
    assign in3180_1 = {c591};
    assign in3180_2 = {c592};
    Full_Adder FA_3180(s3180, c3180, in3180_1, in3180_2, c590);
    wire[0:0] s3181, in3181_1, in3181_2;
    wire c3181;
    assign in3181_1 = {c594};
    assign in3181_2 = {c595};
    Full_Adder FA_3181(s3181, c3181, in3181_1, in3181_2, c593);
    wire[0:0] s3182, in3182_1, in3182_2;
    wire c3182;
    assign in3182_1 = {s597[0]};
    assign in3182_2 = {s598[0]};
    Full_Adder FA_3182(s3182, c3182, in3182_1, in3182_2, s596[0]);
    wire[0:0] s3183, in3183_1, in3183_2;
    wire c3183;
    assign in3183_1 = {s600[0]};
    assign in3183_2 = {s601[0]};
    Full_Adder FA_3183(s3183, c3183, in3183_1, in3183_2, s599[0]);
    wire[0:0] s3184, in3184_1, in3184_2;
    wire c3184;
    assign in3184_1 = {s603[0]};
    assign in3184_2 = {s604[0]};
    Full_Adder FA_3184(s3184, c3184, in3184_1, in3184_2, s602[0]);
    wire[0:0] s3185, in3185_1, in3185_2;
    wire c3185;
    assign in3185_1 = {s606[0]};
    assign in3185_2 = {s607[0]};
    Full_Adder FA_3185(s3185, c3185, in3185_1, in3185_2, s605[0]);
    wire[0:0] s3186, in3186_1, in3186_2;
    wire c3186;
    assign in3186_1 = {s609[0]};
    assign in3186_2 = {s610[0]};
    Full_Adder FA_3186(s3186, c3186, in3186_1, in3186_2, s608[0]);
    wire[0:0] s3187, in3187_1, in3187_2;
    wire c3187;
    assign in3187_1 = {s612[0]};
    assign in3187_2 = {s613[0]};
    Full_Adder FA_3187(s3187, c3187, in3187_1, in3187_2, s611[0]);
    wire[0:0] s3188, in3188_1, in3188_2;
    wire c3188;
    assign in3188_1 = {s615[0]};
    assign in3188_2 = {s616[0]};
    Full_Adder FA_3188(s3188, c3188, in3188_1, in3188_2, s614[0]);
    wire[0:0] s3189, in3189_1, in3189_2;
    wire c3189;
    assign in3189_1 = {s618[0]};
    assign in3189_2 = {s619[0]};
    Full_Adder FA_3189(s3189, c3189, in3189_1, in3189_2, s617[0]);
    wire[0:0] s3190, in3190_1, in3190_2;
    wire c3190;
    assign in3190_1 = {s621[0]};
    assign in3190_2 = {s622[0]};
    Full_Adder FA_3190(s3190, c3190, in3190_1, in3190_2, s620[0]);
    wire[0:0] s3191, in3191_1, in3191_2;
    wire c3191;
    assign in3191_1 = {s624[0]};
    assign in3191_2 = {s625[0]};
    Full_Adder FA_3191(s3191, c3191, in3191_1, in3191_2, s623[0]);
    wire[0:0] s3192, in3192_1, in3192_2;
    wire c3192;
    assign in3192_1 = {s627[0]};
    assign in3192_2 = {s628[0]};
    Full_Adder FA_3192(s3192, c3192, in3192_1, in3192_2, s626[0]);
    wire[0:0] s3193, in3193_1, in3193_2;
    wire c3193;
    assign in3193_1 = {pp108[13]};
    assign in3193_2 = {pp109[12]};
    Full_Adder FA_3193(s3193, c3193, in3193_1, in3193_2, pp107[14]);
    wire[0:0] s3194, in3194_1, in3194_2;
    wire c3194;
    assign in3194_1 = {pp111[10]};
    assign in3194_2 = {pp112[9]};
    Full_Adder FA_3194(s3194, c3194, in3194_1, in3194_2, pp110[11]);
    wire[0:0] s3195, in3195_1, in3195_2;
    wire c3195;
    assign in3195_1 = {pp114[7]};
    assign in3195_2 = {pp115[6]};
    Full_Adder FA_3195(s3195, c3195, in3195_1, in3195_2, pp113[8]);
    wire[0:0] s3196, in3196_1, in3196_2;
    wire c3196;
    assign in3196_1 = {pp117[4]};
    assign in3196_2 = {pp118[3]};
    Full_Adder FA_3196(s3196, c3196, in3196_1, in3196_2, pp116[5]);
    wire[0:0] s3197, in3197_1, in3197_2;
    wire c3197;
    assign in3197_1 = {pp120[1]};
    assign in3197_2 = {pp121[0]};
    Full_Adder FA_3197(s3197, c3197, in3197_1, in3197_2, pp119[2]);
    wire[0:0] s3198, in3198_1, in3198_2;
    wire c3198;
    assign in3198_1 = {c597};
    assign in3198_2 = {c598};
    Full_Adder FA_3198(s3198, c3198, in3198_1, in3198_2, c596);
    wire[0:0] s3199, in3199_1, in3199_2;
    wire c3199;
    assign in3199_1 = {c600};
    assign in3199_2 = {c601};
    Full_Adder FA_3199(s3199, c3199, in3199_1, in3199_2, c599);
    wire[0:0] s3200, in3200_1, in3200_2;
    wire c3200;
    assign in3200_1 = {c603};
    assign in3200_2 = {c604};
    Full_Adder FA_3200(s3200, c3200, in3200_1, in3200_2, c602);
    wire[0:0] s3201, in3201_1, in3201_2;
    wire c3201;
    assign in3201_1 = {c606};
    assign in3201_2 = {c607};
    Full_Adder FA_3201(s3201, c3201, in3201_1, in3201_2, c605);
    wire[0:0] s3202, in3202_1, in3202_2;
    wire c3202;
    assign in3202_1 = {c609};
    assign in3202_2 = {c610};
    Full_Adder FA_3202(s3202, c3202, in3202_1, in3202_2, c608);
    wire[0:0] s3203, in3203_1, in3203_2;
    wire c3203;
    assign in3203_1 = {c612};
    assign in3203_2 = {c613};
    Full_Adder FA_3203(s3203, c3203, in3203_1, in3203_2, c611);
    wire[0:0] s3204, in3204_1, in3204_2;
    wire c3204;
    assign in3204_1 = {c615};
    assign in3204_2 = {c616};
    Full_Adder FA_3204(s3204, c3204, in3204_1, in3204_2, c614);
    wire[0:0] s3205, in3205_1, in3205_2;
    wire c3205;
    assign in3205_1 = {c618};
    assign in3205_2 = {c619};
    Full_Adder FA_3205(s3205, c3205, in3205_1, in3205_2, c617);
    wire[0:0] s3206, in3206_1, in3206_2;
    wire c3206;
    assign in3206_1 = {c621};
    assign in3206_2 = {c622};
    Full_Adder FA_3206(s3206, c3206, in3206_1, in3206_2, c620);
    wire[0:0] s3207, in3207_1, in3207_2;
    wire c3207;
    assign in3207_1 = {c624};
    assign in3207_2 = {c625};
    Full_Adder FA_3207(s3207, c3207, in3207_1, in3207_2, c623);
    wire[0:0] s3208, in3208_1, in3208_2;
    wire c3208;
    assign in3208_1 = {c627};
    assign in3208_2 = {c628};
    Full_Adder FA_3208(s3208, c3208, in3208_1, in3208_2, c626);
    wire[0:0] s3209, in3209_1, in3209_2;
    wire c3209;
    assign in3209_1 = {c630};
    assign in3209_2 = {s631[0]};
    Full_Adder FA_3209(s3209, c3209, in3209_1, in3209_2, c629);
    wire[0:0] s3210, in3210_1, in3210_2;
    wire c3210;
    assign in3210_1 = {s633[0]};
    assign in3210_2 = {s634[0]};
    Full_Adder FA_3210(s3210, c3210, in3210_1, in3210_2, s632[0]);
    wire[0:0] s3211, in3211_1, in3211_2;
    wire c3211;
    assign in3211_1 = {s636[0]};
    assign in3211_2 = {s637[0]};
    Full_Adder FA_3211(s3211, c3211, in3211_1, in3211_2, s635[0]);
    wire[0:0] s3212, in3212_1, in3212_2;
    wire c3212;
    assign in3212_1 = {s639[0]};
    assign in3212_2 = {s640[0]};
    Full_Adder FA_3212(s3212, c3212, in3212_1, in3212_2, s638[0]);
    wire[0:0] s3213, in3213_1, in3213_2;
    wire c3213;
    assign in3213_1 = {s642[0]};
    assign in3213_2 = {s643[0]};
    Full_Adder FA_3213(s3213, c3213, in3213_1, in3213_2, s641[0]);
    wire[0:0] s3214, in3214_1, in3214_2;
    wire c3214;
    assign in3214_1 = {s645[0]};
    assign in3214_2 = {s646[0]};
    Full_Adder FA_3214(s3214, c3214, in3214_1, in3214_2, s644[0]);
    wire[0:0] s3215, in3215_1, in3215_2;
    wire c3215;
    assign in3215_1 = {s648[0]};
    assign in3215_2 = {s649[0]};
    Full_Adder FA_3215(s3215, c3215, in3215_1, in3215_2, s647[0]);
    wire[0:0] s3216, in3216_1, in3216_2;
    wire c3216;
    assign in3216_1 = {s651[0]};
    assign in3216_2 = {s652[0]};
    Full_Adder FA_3216(s3216, c3216, in3216_1, in3216_2, s650[0]);
    wire[0:0] s3217, in3217_1, in3217_2;
    wire c3217;
    assign in3217_1 = {s654[0]};
    assign in3217_2 = {s655[0]};
    Full_Adder FA_3217(s3217, c3217, in3217_1, in3217_2, s653[0]);
    wire[0:0] s3218, in3218_1, in3218_2;
    wire c3218;
    assign in3218_1 = {s657[0]};
    assign in3218_2 = {s658[0]};
    Full_Adder FA_3218(s3218, c3218, in3218_1, in3218_2, s656[0]);
    wire[0:0] s3219, in3219_1, in3219_2;
    wire c3219;
    assign in3219_1 = {s660[0]};
    assign in3219_2 = {s661[0]};
    Full_Adder FA_3219(s3219, c3219, in3219_1, in3219_2, s659[0]);
    wire[0:0] s3220, in3220_1, in3220_2;
    wire c3220;
    assign in3220_1 = {s663[0]};
    assign in3220_2 = {s664[0]};
    Full_Adder FA_3220(s3220, c3220, in3220_1, in3220_2, s662[0]);
    wire[0:0] s3221, in3221_1, in3221_2;
    wire c3221;
    assign in3221_1 = {pp111[11]};
    assign in3221_2 = {pp112[10]};
    Full_Adder FA_3221(s3221, c3221, in3221_1, in3221_2, pp110[12]);
    wire[0:0] s3222, in3222_1, in3222_2;
    wire c3222;
    assign in3222_1 = {pp114[8]};
    assign in3222_2 = {pp115[7]};
    Full_Adder FA_3222(s3222, c3222, in3222_1, in3222_2, pp113[9]);
    wire[0:0] s3223, in3223_1, in3223_2;
    wire c3223;
    assign in3223_1 = {pp117[5]};
    assign in3223_2 = {pp118[4]};
    Full_Adder FA_3223(s3223, c3223, in3223_1, in3223_2, pp116[6]);
    wire[0:0] s3224, in3224_1, in3224_2;
    wire c3224;
    assign in3224_1 = {pp120[2]};
    assign in3224_2 = {pp121[1]};
    Full_Adder FA_3224(s3224, c3224, in3224_1, in3224_2, pp119[3]);
    wire[0:0] s3225, in3225_1, in3225_2;
    wire c3225;
    assign in3225_1 = {c631};
    assign in3225_2 = {c632};
    Full_Adder FA_3225(s3225, c3225, in3225_1, in3225_2, pp122[0]);
    wire[0:0] s3226, in3226_1, in3226_2;
    wire c3226;
    assign in3226_1 = {c634};
    assign in3226_2 = {c635};
    Full_Adder FA_3226(s3226, c3226, in3226_1, in3226_2, c633);
    wire[0:0] s3227, in3227_1, in3227_2;
    wire c3227;
    assign in3227_1 = {c637};
    assign in3227_2 = {c638};
    Full_Adder FA_3227(s3227, c3227, in3227_1, in3227_2, c636);
    wire[0:0] s3228, in3228_1, in3228_2;
    wire c3228;
    assign in3228_1 = {c640};
    assign in3228_2 = {c641};
    Full_Adder FA_3228(s3228, c3228, in3228_1, in3228_2, c639);
    wire[0:0] s3229, in3229_1, in3229_2;
    wire c3229;
    assign in3229_1 = {c643};
    assign in3229_2 = {c644};
    Full_Adder FA_3229(s3229, c3229, in3229_1, in3229_2, c642);
    wire[0:0] s3230, in3230_1, in3230_2;
    wire c3230;
    assign in3230_1 = {c646};
    assign in3230_2 = {c647};
    Full_Adder FA_3230(s3230, c3230, in3230_1, in3230_2, c645);
    wire[0:0] s3231, in3231_1, in3231_2;
    wire c3231;
    assign in3231_1 = {c649};
    assign in3231_2 = {c650};
    Full_Adder FA_3231(s3231, c3231, in3231_1, in3231_2, c648);
    wire[0:0] s3232, in3232_1, in3232_2;
    wire c3232;
    assign in3232_1 = {c652};
    assign in3232_2 = {c653};
    Full_Adder FA_3232(s3232, c3232, in3232_1, in3232_2, c651);
    wire[0:0] s3233, in3233_1, in3233_2;
    wire c3233;
    assign in3233_1 = {c655};
    assign in3233_2 = {c656};
    Full_Adder FA_3233(s3233, c3233, in3233_1, in3233_2, c654);
    wire[0:0] s3234, in3234_1, in3234_2;
    wire c3234;
    assign in3234_1 = {c658};
    assign in3234_2 = {c659};
    Full_Adder FA_3234(s3234, c3234, in3234_1, in3234_2, c657);
    wire[0:0] s3235, in3235_1, in3235_2;
    wire c3235;
    assign in3235_1 = {c661};
    assign in3235_2 = {c662};
    Full_Adder FA_3235(s3235, c3235, in3235_1, in3235_2, c660);
    wire[0:0] s3236, in3236_1, in3236_2;
    wire c3236;
    assign in3236_1 = {c664};
    assign in3236_2 = {c665};
    Full_Adder FA_3236(s3236, c3236, in3236_1, in3236_2, c663);
    wire[0:0] s3237, in3237_1, in3237_2;
    wire c3237;
    assign in3237_1 = {s667[0]};
    assign in3237_2 = {s668[0]};
    Full_Adder FA_3237(s3237, c3237, in3237_1, in3237_2, c666);
    wire[0:0] s3238, in3238_1, in3238_2;
    wire c3238;
    assign in3238_1 = {s670[0]};
    assign in3238_2 = {s671[0]};
    Full_Adder FA_3238(s3238, c3238, in3238_1, in3238_2, s669[0]);
    wire[0:0] s3239, in3239_1, in3239_2;
    wire c3239;
    assign in3239_1 = {s673[0]};
    assign in3239_2 = {s674[0]};
    Full_Adder FA_3239(s3239, c3239, in3239_1, in3239_2, s672[0]);
    wire[0:0] s3240, in3240_1, in3240_2;
    wire c3240;
    assign in3240_1 = {s676[0]};
    assign in3240_2 = {s677[0]};
    Full_Adder FA_3240(s3240, c3240, in3240_1, in3240_2, s675[0]);
    wire[0:0] s3241, in3241_1, in3241_2;
    wire c3241;
    assign in3241_1 = {s679[0]};
    assign in3241_2 = {s680[0]};
    Full_Adder FA_3241(s3241, c3241, in3241_1, in3241_2, s678[0]);
    wire[0:0] s3242, in3242_1, in3242_2;
    wire c3242;
    assign in3242_1 = {s682[0]};
    assign in3242_2 = {s683[0]};
    Full_Adder FA_3242(s3242, c3242, in3242_1, in3242_2, s681[0]);
    wire[0:0] s3243, in3243_1, in3243_2;
    wire c3243;
    assign in3243_1 = {s685[0]};
    assign in3243_2 = {s686[0]};
    Full_Adder FA_3243(s3243, c3243, in3243_1, in3243_2, s684[0]);
    wire[0:0] s3244, in3244_1, in3244_2;
    wire c3244;
    assign in3244_1 = {s688[0]};
    assign in3244_2 = {s689[0]};
    Full_Adder FA_3244(s3244, c3244, in3244_1, in3244_2, s687[0]);
    wire[0:0] s3245, in3245_1, in3245_2;
    wire c3245;
    assign in3245_1 = {s691[0]};
    assign in3245_2 = {s692[0]};
    Full_Adder FA_3245(s3245, c3245, in3245_1, in3245_2, s690[0]);
    wire[0:0] s3246, in3246_1, in3246_2;
    wire c3246;
    assign in3246_1 = {s694[0]};
    assign in3246_2 = {s695[0]};
    Full_Adder FA_3246(s3246, c3246, in3246_1, in3246_2, s693[0]);
    wire[0:0] s3247, in3247_1, in3247_2;
    wire c3247;
    assign in3247_1 = {s697[0]};
    assign in3247_2 = {s698[0]};
    Full_Adder FA_3247(s3247, c3247, in3247_1, in3247_2, s696[0]);
    wire[0:0] s3248, in3248_1, in3248_2;
    wire c3248;
    assign in3248_1 = {s700[0]};
    assign in3248_2 = {s701[0]};
    Full_Adder FA_3248(s3248, c3248, in3248_1, in3248_2, s699[0]);
    wire[0:0] s3249, in3249_1, in3249_2;
    wire c3249;
    assign in3249_1 = {pp114[9]};
    assign in3249_2 = {pp115[8]};
    Full_Adder FA_3249(s3249, c3249, in3249_1, in3249_2, pp113[10]);
    wire[0:0] s3250, in3250_1, in3250_2;
    wire c3250;
    assign in3250_1 = {pp117[6]};
    assign in3250_2 = {pp118[5]};
    Full_Adder FA_3250(s3250, c3250, in3250_1, in3250_2, pp116[7]);
    wire[0:0] s3251, in3251_1, in3251_2;
    wire c3251;
    assign in3251_1 = {pp120[3]};
    assign in3251_2 = {pp121[2]};
    Full_Adder FA_3251(s3251, c3251, in3251_1, in3251_2, pp119[4]);
    wire[0:0] s3252, in3252_1, in3252_2;
    wire c3252;
    assign in3252_1 = {pp123[0]};
    assign in3252_2 = {c667};
    Full_Adder FA_3252(s3252, c3252, in3252_1, in3252_2, pp122[1]);
    wire[0:0] s3253, in3253_1, in3253_2;
    wire c3253;
    assign in3253_1 = {c669};
    assign in3253_2 = {c670};
    Full_Adder FA_3253(s3253, c3253, in3253_1, in3253_2, c668);
    wire[0:0] s3254, in3254_1, in3254_2;
    wire c3254;
    assign in3254_1 = {c672};
    assign in3254_2 = {c673};
    Full_Adder FA_3254(s3254, c3254, in3254_1, in3254_2, c671);
    wire[0:0] s3255, in3255_1, in3255_2;
    wire c3255;
    assign in3255_1 = {c675};
    assign in3255_2 = {c676};
    Full_Adder FA_3255(s3255, c3255, in3255_1, in3255_2, c674);
    wire[0:0] s3256, in3256_1, in3256_2;
    wire c3256;
    assign in3256_1 = {c678};
    assign in3256_2 = {c679};
    Full_Adder FA_3256(s3256, c3256, in3256_1, in3256_2, c677);
    wire[0:0] s3257, in3257_1, in3257_2;
    wire c3257;
    assign in3257_1 = {c681};
    assign in3257_2 = {c682};
    Full_Adder FA_3257(s3257, c3257, in3257_1, in3257_2, c680);
    wire[0:0] s3258, in3258_1, in3258_2;
    wire c3258;
    assign in3258_1 = {c684};
    assign in3258_2 = {c685};
    Full_Adder FA_3258(s3258, c3258, in3258_1, in3258_2, c683);
    wire[0:0] s3259, in3259_1, in3259_2;
    wire c3259;
    assign in3259_1 = {c687};
    assign in3259_2 = {c688};
    Full_Adder FA_3259(s3259, c3259, in3259_1, in3259_2, c686);
    wire[0:0] s3260, in3260_1, in3260_2;
    wire c3260;
    assign in3260_1 = {c690};
    assign in3260_2 = {c691};
    Full_Adder FA_3260(s3260, c3260, in3260_1, in3260_2, c689);
    wire[0:0] s3261, in3261_1, in3261_2;
    wire c3261;
    assign in3261_1 = {c693};
    assign in3261_2 = {c694};
    Full_Adder FA_3261(s3261, c3261, in3261_1, in3261_2, c692);
    wire[0:0] s3262, in3262_1, in3262_2;
    wire c3262;
    assign in3262_1 = {c696};
    assign in3262_2 = {c697};
    Full_Adder FA_3262(s3262, c3262, in3262_1, in3262_2, c695);
    wire[0:0] s3263, in3263_1, in3263_2;
    wire c3263;
    assign in3263_1 = {c699};
    assign in3263_2 = {c700};
    Full_Adder FA_3263(s3263, c3263, in3263_1, in3263_2, c698);
    wire[0:0] s3264, in3264_1, in3264_2;
    wire c3264;
    assign in3264_1 = {c702};
    assign in3264_2 = {c703};
    Full_Adder FA_3264(s3264, c3264, in3264_1, in3264_2, c701);
    wire[0:0] s3265, in3265_1, in3265_2;
    wire c3265;
    assign in3265_1 = {s705[0]};
    assign in3265_2 = {s706[0]};
    Full_Adder FA_3265(s3265, c3265, in3265_1, in3265_2, s704[0]);
    wire[0:0] s3266, in3266_1, in3266_2;
    wire c3266;
    assign in3266_1 = {s708[0]};
    assign in3266_2 = {s709[0]};
    Full_Adder FA_3266(s3266, c3266, in3266_1, in3266_2, s707[0]);
    wire[0:0] s3267, in3267_1, in3267_2;
    wire c3267;
    assign in3267_1 = {s711[0]};
    assign in3267_2 = {s712[0]};
    Full_Adder FA_3267(s3267, c3267, in3267_1, in3267_2, s710[0]);
    wire[0:0] s3268, in3268_1, in3268_2;
    wire c3268;
    assign in3268_1 = {s714[0]};
    assign in3268_2 = {s715[0]};
    Full_Adder FA_3268(s3268, c3268, in3268_1, in3268_2, s713[0]);
    wire[0:0] s3269, in3269_1, in3269_2;
    wire c3269;
    assign in3269_1 = {s717[0]};
    assign in3269_2 = {s718[0]};
    Full_Adder FA_3269(s3269, c3269, in3269_1, in3269_2, s716[0]);
    wire[0:0] s3270, in3270_1, in3270_2;
    wire c3270;
    assign in3270_1 = {s720[0]};
    assign in3270_2 = {s721[0]};
    Full_Adder FA_3270(s3270, c3270, in3270_1, in3270_2, s719[0]);
    wire[0:0] s3271, in3271_1, in3271_2;
    wire c3271;
    assign in3271_1 = {s723[0]};
    assign in3271_2 = {s724[0]};
    Full_Adder FA_3271(s3271, c3271, in3271_1, in3271_2, s722[0]);
    wire[0:0] s3272, in3272_1, in3272_2;
    wire c3272;
    assign in3272_1 = {s726[0]};
    assign in3272_2 = {s727[0]};
    Full_Adder FA_3272(s3272, c3272, in3272_1, in3272_2, s725[0]);
    wire[0:0] s3273, in3273_1, in3273_2;
    wire c3273;
    assign in3273_1 = {s729[0]};
    assign in3273_2 = {s730[0]};
    Full_Adder FA_3273(s3273, c3273, in3273_1, in3273_2, s728[0]);
    wire[0:0] s3274, in3274_1, in3274_2;
    wire c3274;
    assign in3274_1 = {s732[0]};
    assign in3274_2 = {s733[0]};
    Full_Adder FA_3274(s3274, c3274, in3274_1, in3274_2, s731[0]);
    wire[0:0] s3275, in3275_1, in3275_2;
    wire c3275;
    assign in3275_1 = {s735[0]};
    assign in3275_2 = {s736[0]};
    Full_Adder FA_3275(s3275, c3275, in3275_1, in3275_2, s734[0]);
    wire[0:0] s3276, in3276_1, in3276_2;
    wire c3276;
    assign in3276_1 = {s738[0]};
    assign in3276_2 = {s739[0]};
    Full_Adder FA_3276(s3276, c3276, in3276_1, in3276_2, s737[0]);
    wire[0:0] s3277, in3277_1, in3277_2;
    wire c3277;
    assign in3277_1 = {pp117[7]};
    assign in3277_2 = {pp118[6]};
    Full_Adder FA_3277(s3277, c3277, in3277_1, in3277_2, pp116[8]);
    wire[0:0] s3278, in3278_1, in3278_2;
    wire c3278;
    assign in3278_1 = {pp120[4]};
    assign in3278_2 = {pp121[3]};
    Full_Adder FA_3278(s3278, c3278, in3278_1, in3278_2, pp119[5]);
    wire[0:0] s3279, in3279_1, in3279_2;
    wire c3279;
    assign in3279_1 = {pp123[1]};
    assign in3279_2 = {pp124[0]};
    Full_Adder FA_3279(s3279, c3279, in3279_1, in3279_2, pp122[2]);
    wire[0:0] s3280, in3280_1, in3280_2;
    wire c3280;
    assign in3280_1 = {c705};
    assign in3280_2 = {c706};
    Full_Adder FA_3280(s3280, c3280, in3280_1, in3280_2, c704);
    wire[0:0] s3281, in3281_1, in3281_2;
    wire c3281;
    assign in3281_1 = {c708};
    assign in3281_2 = {c709};
    Full_Adder FA_3281(s3281, c3281, in3281_1, in3281_2, c707);
    wire[0:0] s3282, in3282_1, in3282_2;
    wire c3282;
    assign in3282_1 = {c711};
    assign in3282_2 = {c712};
    Full_Adder FA_3282(s3282, c3282, in3282_1, in3282_2, c710);
    wire[0:0] s3283, in3283_1, in3283_2;
    wire c3283;
    assign in3283_1 = {c714};
    assign in3283_2 = {c715};
    Full_Adder FA_3283(s3283, c3283, in3283_1, in3283_2, c713);
    wire[0:0] s3284, in3284_1, in3284_2;
    wire c3284;
    assign in3284_1 = {c717};
    assign in3284_2 = {c718};
    Full_Adder FA_3284(s3284, c3284, in3284_1, in3284_2, c716);
    wire[0:0] s3285, in3285_1, in3285_2;
    wire c3285;
    assign in3285_1 = {c720};
    assign in3285_2 = {c721};
    Full_Adder FA_3285(s3285, c3285, in3285_1, in3285_2, c719);
    wire[0:0] s3286, in3286_1, in3286_2;
    wire c3286;
    assign in3286_1 = {c723};
    assign in3286_2 = {c724};
    Full_Adder FA_3286(s3286, c3286, in3286_1, in3286_2, c722);
    wire[0:0] s3287, in3287_1, in3287_2;
    wire c3287;
    assign in3287_1 = {c726};
    assign in3287_2 = {c727};
    Full_Adder FA_3287(s3287, c3287, in3287_1, in3287_2, c725);
    wire[0:0] s3288, in3288_1, in3288_2;
    wire c3288;
    assign in3288_1 = {c729};
    assign in3288_2 = {c730};
    Full_Adder FA_3288(s3288, c3288, in3288_1, in3288_2, c728);
    wire[0:0] s3289, in3289_1, in3289_2;
    wire c3289;
    assign in3289_1 = {c732};
    assign in3289_2 = {c733};
    Full_Adder FA_3289(s3289, c3289, in3289_1, in3289_2, c731);
    wire[0:0] s3290, in3290_1, in3290_2;
    wire c3290;
    assign in3290_1 = {c735};
    assign in3290_2 = {c736};
    Full_Adder FA_3290(s3290, c3290, in3290_1, in3290_2, c734);
    wire[0:0] s3291, in3291_1, in3291_2;
    wire c3291;
    assign in3291_1 = {c738};
    assign in3291_2 = {c739};
    Full_Adder FA_3291(s3291, c3291, in3291_1, in3291_2, c737);
    wire[0:0] s3292, in3292_1, in3292_2;
    wire c3292;
    assign in3292_1 = {c741};
    assign in3292_2 = {s742[0]};
    Full_Adder FA_3292(s3292, c3292, in3292_1, in3292_2, c740);
    wire[0:0] s3293, in3293_1, in3293_2;
    wire c3293;
    assign in3293_1 = {s744[0]};
    assign in3293_2 = {s745[0]};
    Full_Adder FA_3293(s3293, c3293, in3293_1, in3293_2, s743[0]);
    wire[0:0] s3294, in3294_1, in3294_2;
    wire c3294;
    assign in3294_1 = {s747[0]};
    assign in3294_2 = {s748[0]};
    Full_Adder FA_3294(s3294, c3294, in3294_1, in3294_2, s746[0]);
    wire[0:0] s3295, in3295_1, in3295_2;
    wire c3295;
    assign in3295_1 = {s750[0]};
    assign in3295_2 = {s751[0]};
    Full_Adder FA_3295(s3295, c3295, in3295_1, in3295_2, s749[0]);
    wire[0:0] s3296, in3296_1, in3296_2;
    wire c3296;
    assign in3296_1 = {s753[0]};
    assign in3296_2 = {s754[0]};
    Full_Adder FA_3296(s3296, c3296, in3296_1, in3296_2, s752[0]);
    wire[0:0] s3297, in3297_1, in3297_2;
    wire c3297;
    assign in3297_1 = {s756[0]};
    assign in3297_2 = {s757[0]};
    Full_Adder FA_3297(s3297, c3297, in3297_1, in3297_2, s755[0]);
    wire[0:0] s3298, in3298_1, in3298_2;
    wire c3298;
    assign in3298_1 = {s759[0]};
    assign in3298_2 = {s760[0]};
    Full_Adder FA_3298(s3298, c3298, in3298_1, in3298_2, s758[0]);
    wire[0:0] s3299, in3299_1, in3299_2;
    wire c3299;
    assign in3299_1 = {s762[0]};
    assign in3299_2 = {s763[0]};
    Full_Adder FA_3299(s3299, c3299, in3299_1, in3299_2, s761[0]);
    wire[0:0] s3300, in3300_1, in3300_2;
    wire c3300;
    assign in3300_1 = {s765[0]};
    assign in3300_2 = {s766[0]};
    Full_Adder FA_3300(s3300, c3300, in3300_1, in3300_2, s764[0]);
    wire[0:0] s3301, in3301_1, in3301_2;
    wire c3301;
    assign in3301_1 = {s768[0]};
    assign in3301_2 = {s769[0]};
    Full_Adder FA_3301(s3301, c3301, in3301_1, in3301_2, s767[0]);
    wire[0:0] s3302, in3302_1, in3302_2;
    wire c3302;
    assign in3302_1 = {s771[0]};
    assign in3302_2 = {s772[0]};
    Full_Adder FA_3302(s3302, c3302, in3302_1, in3302_2, s770[0]);
    wire[0:0] s3303, in3303_1, in3303_2;
    wire c3303;
    assign in3303_1 = {s774[0]};
    assign in3303_2 = {s775[0]};
    Full_Adder FA_3303(s3303, c3303, in3303_1, in3303_2, s773[0]);
    wire[0:0] s3304, in3304_1, in3304_2;
    wire c3304;
    assign in3304_1 = {s777[0]};
    assign in3304_2 = {s778[0]};
    Full_Adder FA_3304(s3304, c3304, in3304_1, in3304_2, s776[0]);
    wire[0:0] s3305, in3305_1, in3305_2;
    wire c3305;
    assign in3305_1 = {pp120[5]};
    assign in3305_2 = {pp121[4]};
    Full_Adder FA_3305(s3305, c3305, in3305_1, in3305_2, pp119[6]);
    wire[0:0] s3306, in3306_1, in3306_2;
    wire c3306;
    assign in3306_1 = {pp123[2]};
    assign in3306_2 = {pp124[1]};
    Full_Adder FA_3306(s3306, c3306, in3306_1, in3306_2, pp122[3]);
    wire[0:0] s3307, in3307_1, in3307_2;
    wire c3307;
    assign in3307_1 = {c742};
    assign in3307_2 = {c743};
    Full_Adder FA_3307(s3307, c3307, in3307_1, in3307_2, pp125[0]);
    wire[0:0] s3308, in3308_1, in3308_2;
    wire c3308;
    assign in3308_1 = {c745};
    assign in3308_2 = {c746};
    Full_Adder FA_3308(s3308, c3308, in3308_1, in3308_2, c744);
    wire[0:0] s3309, in3309_1, in3309_2;
    wire c3309;
    assign in3309_1 = {c748};
    assign in3309_2 = {c749};
    Full_Adder FA_3309(s3309, c3309, in3309_1, in3309_2, c747);
    wire[0:0] s3310, in3310_1, in3310_2;
    wire c3310;
    assign in3310_1 = {c751};
    assign in3310_2 = {c752};
    Full_Adder FA_3310(s3310, c3310, in3310_1, in3310_2, c750);
    wire[0:0] s3311, in3311_1, in3311_2;
    wire c3311;
    assign in3311_1 = {c754};
    assign in3311_2 = {c755};
    Full_Adder FA_3311(s3311, c3311, in3311_1, in3311_2, c753);
    wire[0:0] s3312, in3312_1, in3312_2;
    wire c3312;
    assign in3312_1 = {c757};
    assign in3312_2 = {c758};
    Full_Adder FA_3312(s3312, c3312, in3312_1, in3312_2, c756);
    wire[0:0] s3313, in3313_1, in3313_2;
    wire c3313;
    assign in3313_1 = {c760};
    assign in3313_2 = {c761};
    Full_Adder FA_3313(s3313, c3313, in3313_1, in3313_2, c759);
    wire[0:0] s3314, in3314_1, in3314_2;
    wire c3314;
    assign in3314_1 = {c763};
    assign in3314_2 = {c764};
    Full_Adder FA_3314(s3314, c3314, in3314_1, in3314_2, c762);
    wire[0:0] s3315, in3315_1, in3315_2;
    wire c3315;
    assign in3315_1 = {c766};
    assign in3315_2 = {c767};
    Full_Adder FA_3315(s3315, c3315, in3315_1, in3315_2, c765);
    wire[0:0] s3316, in3316_1, in3316_2;
    wire c3316;
    assign in3316_1 = {c769};
    assign in3316_2 = {c770};
    Full_Adder FA_3316(s3316, c3316, in3316_1, in3316_2, c768);
    wire[0:0] s3317, in3317_1, in3317_2;
    wire c3317;
    assign in3317_1 = {c772};
    assign in3317_2 = {c773};
    Full_Adder FA_3317(s3317, c3317, in3317_1, in3317_2, c771);
    wire[0:0] s3318, in3318_1, in3318_2;
    wire c3318;
    assign in3318_1 = {c775};
    assign in3318_2 = {c776};
    Full_Adder FA_3318(s3318, c3318, in3318_1, in3318_2, c774);
    wire[0:0] s3319, in3319_1, in3319_2;
    wire c3319;
    assign in3319_1 = {c778};
    assign in3319_2 = {c779};
    Full_Adder FA_3319(s3319, c3319, in3319_1, in3319_2, c777);
    wire[0:0] s3320, in3320_1, in3320_2;
    wire c3320;
    assign in3320_1 = {s781[0]};
    assign in3320_2 = {s782[0]};
    Full_Adder FA_3320(s3320, c3320, in3320_1, in3320_2, c780);
    wire[0:0] s3321, in3321_1, in3321_2;
    wire c3321;
    assign in3321_1 = {s784[0]};
    assign in3321_2 = {s785[0]};
    Full_Adder FA_3321(s3321, c3321, in3321_1, in3321_2, s783[0]);
    wire[0:0] s3322, in3322_1, in3322_2;
    wire c3322;
    assign in3322_1 = {s787[0]};
    assign in3322_2 = {s788[0]};
    Full_Adder FA_3322(s3322, c3322, in3322_1, in3322_2, s786[0]);
    wire[0:0] s3323, in3323_1, in3323_2;
    wire c3323;
    assign in3323_1 = {s790[0]};
    assign in3323_2 = {s791[0]};
    Full_Adder FA_3323(s3323, c3323, in3323_1, in3323_2, s789[0]);
    wire[0:0] s3324, in3324_1, in3324_2;
    wire c3324;
    assign in3324_1 = {s793[0]};
    assign in3324_2 = {s794[0]};
    Full_Adder FA_3324(s3324, c3324, in3324_1, in3324_2, s792[0]);
    wire[0:0] s3325, in3325_1, in3325_2;
    wire c3325;
    assign in3325_1 = {s796[0]};
    assign in3325_2 = {s797[0]};
    Full_Adder FA_3325(s3325, c3325, in3325_1, in3325_2, s795[0]);
    wire[0:0] s3326, in3326_1, in3326_2;
    wire c3326;
    assign in3326_1 = {s799[0]};
    assign in3326_2 = {s800[0]};
    Full_Adder FA_3326(s3326, c3326, in3326_1, in3326_2, s798[0]);
    wire[0:0] s3327, in3327_1, in3327_2;
    wire c3327;
    assign in3327_1 = {s802[0]};
    assign in3327_2 = {s803[0]};
    Full_Adder FA_3327(s3327, c3327, in3327_1, in3327_2, s801[0]);
    wire[0:0] s3328, in3328_1, in3328_2;
    wire c3328;
    assign in3328_1 = {s805[0]};
    assign in3328_2 = {s806[0]};
    Full_Adder FA_3328(s3328, c3328, in3328_1, in3328_2, s804[0]);
    wire[0:0] s3329, in3329_1, in3329_2;
    wire c3329;
    assign in3329_1 = {s808[0]};
    assign in3329_2 = {s809[0]};
    Full_Adder FA_3329(s3329, c3329, in3329_1, in3329_2, s807[0]);
    wire[0:0] s3330, in3330_1, in3330_2;
    wire c3330;
    assign in3330_1 = {s811[0]};
    assign in3330_2 = {s812[0]};
    Full_Adder FA_3330(s3330, c3330, in3330_1, in3330_2, s810[0]);
    wire[0:0] s3331, in3331_1, in3331_2;
    wire c3331;
    assign in3331_1 = {s814[0]};
    assign in3331_2 = {s815[0]};
    Full_Adder FA_3331(s3331, c3331, in3331_1, in3331_2, s813[0]);
    wire[0:0] s3332, in3332_1, in3332_2;
    wire c3332;
    assign in3332_1 = {s817[0]};
    assign in3332_2 = {s818[0]};
    Full_Adder FA_3332(s3332, c3332, in3332_1, in3332_2, s816[0]);
    wire[0:0] s3333, in3333_1, in3333_2;
    wire c3333;
    assign in3333_1 = {pp123[3]};
    assign in3333_2 = {pp124[2]};
    Full_Adder FA_3333(s3333, c3333, in3333_1, in3333_2, pp122[4]);
    wire[0:0] s3334, in3334_1, in3334_2;
    wire c3334;
    assign in3334_1 = {pp126[0]};
    assign in3334_2 = {c781};
    Full_Adder FA_3334(s3334, c3334, in3334_1, in3334_2, pp125[1]);
    wire[0:0] s3335, in3335_1, in3335_2;
    wire c3335;
    assign in3335_1 = {c783};
    assign in3335_2 = {c784};
    Full_Adder FA_3335(s3335, c3335, in3335_1, in3335_2, c782);
    wire[0:0] s3336, in3336_1, in3336_2;
    wire c3336;
    assign in3336_1 = {c786};
    assign in3336_2 = {c787};
    Full_Adder FA_3336(s3336, c3336, in3336_1, in3336_2, c785);
    wire[0:0] s3337, in3337_1, in3337_2;
    wire c3337;
    assign in3337_1 = {c789};
    assign in3337_2 = {c790};
    Full_Adder FA_3337(s3337, c3337, in3337_1, in3337_2, c788);
    wire[0:0] s3338, in3338_1, in3338_2;
    wire c3338;
    assign in3338_1 = {c792};
    assign in3338_2 = {c793};
    Full_Adder FA_3338(s3338, c3338, in3338_1, in3338_2, c791);
    wire[0:0] s3339, in3339_1, in3339_2;
    wire c3339;
    assign in3339_1 = {c795};
    assign in3339_2 = {c796};
    Full_Adder FA_3339(s3339, c3339, in3339_1, in3339_2, c794);
    wire[0:0] s3340, in3340_1, in3340_2;
    wire c3340;
    assign in3340_1 = {c798};
    assign in3340_2 = {c799};
    Full_Adder FA_3340(s3340, c3340, in3340_1, in3340_2, c797);
    wire[0:0] s3341, in3341_1, in3341_2;
    wire c3341;
    assign in3341_1 = {c801};
    assign in3341_2 = {c802};
    Full_Adder FA_3341(s3341, c3341, in3341_1, in3341_2, c800);
    wire[0:0] s3342, in3342_1, in3342_2;
    wire c3342;
    assign in3342_1 = {c804};
    assign in3342_2 = {c805};
    Full_Adder FA_3342(s3342, c3342, in3342_1, in3342_2, c803);
    wire[0:0] s3343, in3343_1, in3343_2;
    wire c3343;
    assign in3343_1 = {c807};
    assign in3343_2 = {c808};
    Full_Adder FA_3343(s3343, c3343, in3343_1, in3343_2, c806);
    wire[0:0] s3344, in3344_1, in3344_2;
    wire c3344;
    assign in3344_1 = {c810};
    assign in3344_2 = {c811};
    Full_Adder FA_3344(s3344, c3344, in3344_1, in3344_2, c809);
    wire[0:0] s3345, in3345_1, in3345_2;
    wire c3345;
    assign in3345_1 = {c813};
    assign in3345_2 = {c814};
    Full_Adder FA_3345(s3345, c3345, in3345_1, in3345_2, c812);
    wire[0:0] s3346, in3346_1, in3346_2;
    wire c3346;
    assign in3346_1 = {c816};
    assign in3346_2 = {c817};
    Full_Adder FA_3346(s3346, c3346, in3346_1, in3346_2, c815);
    wire[0:0] s3347, in3347_1, in3347_2;
    wire c3347;
    assign in3347_1 = {c819};
    assign in3347_2 = {c820};
    Full_Adder FA_3347(s3347, c3347, in3347_1, in3347_2, c818);
    wire[0:0] s3348, in3348_1, in3348_2;
    wire c3348;
    assign in3348_1 = {s822[0]};
    assign in3348_2 = {s823[0]};
    Full_Adder FA_3348(s3348, c3348, in3348_1, in3348_2, s821[0]);
    wire[0:0] s3349, in3349_1, in3349_2;
    wire c3349;
    assign in3349_1 = {s825[0]};
    assign in3349_2 = {s826[0]};
    Full_Adder FA_3349(s3349, c3349, in3349_1, in3349_2, s824[0]);
    wire[0:0] s3350, in3350_1, in3350_2;
    wire c3350;
    assign in3350_1 = {s828[0]};
    assign in3350_2 = {s829[0]};
    Full_Adder FA_3350(s3350, c3350, in3350_1, in3350_2, s827[0]);
    wire[0:0] s3351, in3351_1, in3351_2;
    wire c3351;
    assign in3351_1 = {s831[0]};
    assign in3351_2 = {s832[0]};
    Full_Adder FA_3351(s3351, c3351, in3351_1, in3351_2, s830[0]);
    wire[0:0] s3352, in3352_1, in3352_2;
    wire c3352;
    assign in3352_1 = {s834[0]};
    assign in3352_2 = {s835[0]};
    Full_Adder FA_3352(s3352, c3352, in3352_1, in3352_2, s833[0]);
    wire[0:0] s3353, in3353_1, in3353_2;
    wire c3353;
    assign in3353_1 = {s837[0]};
    assign in3353_2 = {s838[0]};
    Full_Adder FA_3353(s3353, c3353, in3353_1, in3353_2, s836[0]);
    wire[0:0] s3354, in3354_1, in3354_2;
    wire c3354;
    assign in3354_1 = {s840[0]};
    assign in3354_2 = {s841[0]};
    Full_Adder FA_3354(s3354, c3354, in3354_1, in3354_2, s839[0]);
    wire[0:0] s3355, in3355_1, in3355_2;
    wire c3355;
    assign in3355_1 = {s843[0]};
    assign in3355_2 = {s844[0]};
    Full_Adder FA_3355(s3355, c3355, in3355_1, in3355_2, s842[0]);
    wire[0:0] s3356, in3356_1, in3356_2;
    wire c3356;
    assign in3356_1 = {s846[0]};
    assign in3356_2 = {s847[0]};
    Full_Adder FA_3356(s3356, c3356, in3356_1, in3356_2, s845[0]);
    wire[0:0] s3357, in3357_1, in3357_2;
    wire c3357;
    assign in3357_1 = {s849[0]};
    assign in3357_2 = {s850[0]};
    Full_Adder FA_3357(s3357, c3357, in3357_1, in3357_2, s848[0]);
    wire[0:0] s3358, in3358_1, in3358_2;
    wire c3358;
    assign in3358_1 = {s852[0]};
    assign in3358_2 = {s853[0]};
    Full_Adder FA_3358(s3358, c3358, in3358_1, in3358_2, s851[0]);
    wire[0:0] s3359, in3359_1, in3359_2;
    wire c3359;
    assign in3359_1 = {s855[0]};
    assign in3359_2 = {s856[0]};
    Full_Adder FA_3359(s3359, c3359, in3359_1, in3359_2, s854[0]);
    wire[0:0] s3360, in3360_1, in3360_2;
    wire c3360;
    assign in3360_1 = {s858[0]};
    assign in3360_2 = {s859[0]};
    Full_Adder FA_3360(s3360, c3360, in3360_1, in3360_2, s857[0]);
    wire[0:0] s3361, in3361_1, in3361_2;
    wire c3361;
    assign in3361_1 = {pp126[1]};
    assign in3361_2 = {pp127[0]};
    Full_Adder FA_3361(s3361, c3361, in3361_1, in3361_2, pp125[2]);
    wire[0:0] s3362, in3362_1, in3362_2;
    wire c3362;
    assign in3362_1 = {c822};
    assign in3362_2 = {c823};
    Full_Adder FA_3362(s3362, c3362, in3362_1, in3362_2, c821);
    wire[0:0] s3363, in3363_1, in3363_2;
    wire c3363;
    assign in3363_1 = {c825};
    assign in3363_2 = {c826};
    Full_Adder FA_3363(s3363, c3363, in3363_1, in3363_2, c824);
    wire[0:0] s3364, in3364_1, in3364_2;
    wire c3364;
    assign in3364_1 = {c828};
    assign in3364_2 = {c829};
    Full_Adder FA_3364(s3364, c3364, in3364_1, in3364_2, c827);
    wire[0:0] s3365, in3365_1, in3365_2;
    wire c3365;
    assign in3365_1 = {c831};
    assign in3365_2 = {c832};
    Full_Adder FA_3365(s3365, c3365, in3365_1, in3365_2, c830);
    wire[0:0] s3366, in3366_1, in3366_2;
    wire c3366;
    assign in3366_1 = {c834};
    assign in3366_2 = {c835};
    Full_Adder FA_3366(s3366, c3366, in3366_1, in3366_2, c833);
    wire[0:0] s3367, in3367_1, in3367_2;
    wire c3367;
    assign in3367_1 = {c837};
    assign in3367_2 = {c838};
    Full_Adder FA_3367(s3367, c3367, in3367_1, in3367_2, c836);
    wire[0:0] s3368, in3368_1, in3368_2;
    wire c3368;
    assign in3368_1 = {c840};
    assign in3368_2 = {c841};
    Full_Adder FA_3368(s3368, c3368, in3368_1, in3368_2, c839);
    wire[0:0] s3369, in3369_1, in3369_2;
    wire c3369;
    assign in3369_1 = {c843};
    assign in3369_2 = {c844};
    Full_Adder FA_3369(s3369, c3369, in3369_1, in3369_2, c842);
    wire[0:0] s3370, in3370_1, in3370_2;
    wire c3370;
    assign in3370_1 = {c846};
    assign in3370_2 = {c847};
    Full_Adder FA_3370(s3370, c3370, in3370_1, in3370_2, c845);
    wire[0:0] s3371, in3371_1, in3371_2;
    wire c3371;
    assign in3371_1 = {c849};
    assign in3371_2 = {c850};
    Full_Adder FA_3371(s3371, c3371, in3371_1, in3371_2, c848);
    wire[0:0] s3372, in3372_1, in3372_2;
    wire c3372;
    assign in3372_1 = {c852};
    assign in3372_2 = {c853};
    Full_Adder FA_3372(s3372, c3372, in3372_1, in3372_2, c851);
    wire[0:0] s3373, in3373_1, in3373_2;
    wire c3373;
    assign in3373_1 = {c855};
    assign in3373_2 = {c856};
    Full_Adder FA_3373(s3373, c3373, in3373_1, in3373_2, c854);
    wire[0:0] s3374, in3374_1, in3374_2;
    wire c3374;
    assign in3374_1 = {c858};
    assign in3374_2 = {c859};
    Full_Adder FA_3374(s3374, c3374, in3374_1, in3374_2, c857);
    wire[0:0] s3375, in3375_1, in3375_2;
    wire c3375;
    assign in3375_1 = {c861};
    assign in3375_2 = {s862[0]};
    Full_Adder FA_3375(s3375, c3375, in3375_1, in3375_2, c860);
    wire[0:0] s3376, in3376_1, in3376_2;
    wire c3376;
    assign in3376_1 = {s864[0]};
    assign in3376_2 = {s865[0]};
    Full_Adder FA_3376(s3376, c3376, in3376_1, in3376_2, s863[0]);
    wire[0:0] s3377, in3377_1, in3377_2;
    wire c3377;
    assign in3377_1 = {s867[0]};
    assign in3377_2 = {s868[0]};
    Full_Adder FA_3377(s3377, c3377, in3377_1, in3377_2, s866[0]);
    wire[0:0] s3378, in3378_1, in3378_2;
    wire c3378;
    assign in3378_1 = {s870[0]};
    assign in3378_2 = {s871[0]};
    Full_Adder FA_3378(s3378, c3378, in3378_1, in3378_2, s869[0]);
    wire[0:0] s3379, in3379_1, in3379_2;
    wire c3379;
    assign in3379_1 = {s873[0]};
    assign in3379_2 = {s874[0]};
    Full_Adder FA_3379(s3379, c3379, in3379_1, in3379_2, s872[0]);
    wire[0:0] s3380, in3380_1, in3380_2;
    wire c3380;
    assign in3380_1 = {s876[0]};
    assign in3380_2 = {s877[0]};
    Full_Adder FA_3380(s3380, c3380, in3380_1, in3380_2, s875[0]);
    wire[0:0] s3381, in3381_1, in3381_2;
    wire c3381;
    assign in3381_1 = {s879[0]};
    assign in3381_2 = {s880[0]};
    Full_Adder FA_3381(s3381, c3381, in3381_1, in3381_2, s878[0]);
    wire[0:0] s3382, in3382_1, in3382_2;
    wire c3382;
    assign in3382_1 = {s882[0]};
    assign in3382_2 = {s883[0]};
    Full_Adder FA_3382(s3382, c3382, in3382_1, in3382_2, s881[0]);
    wire[0:0] s3383, in3383_1, in3383_2;
    wire c3383;
    assign in3383_1 = {s885[0]};
    assign in3383_2 = {s886[0]};
    Full_Adder FA_3383(s3383, c3383, in3383_1, in3383_2, s884[0]);
    wire[0:0] s3384, in3384_1, in3384_2;
    wire c3384;
    assign in3384_1 = {s888[0]};
    assign in3384_2 = {s889[0]};
    Full_Adder FA_3384(s3384, c3384, in3384_1, in3384_2, s887[0]);
    wire[0:0] s3385, in3385_1, in3385_2;
    wire c3385;
    assign in3385_1 = {s891[0]};
    assign in3385_2 = {s892[0]};
    Full_Adder FA_3385(s3385, c3385, in3385_1, in3385_2, s890[0]);
    wire[0:0] s3386, in3386_1, in3386_2;
    wire c3386;
    assign in3386_1 = {s894[0]};
    assign in3386_2 = {s895[0]};
    Full_Adder FA_3386(s3386, c3386, in3386_1, in3386_2, s893[0]);
    wire[0:0] s3387, in3387_1, in3387_2;
    wire c3387;
    assign in3387_1 = {s897[0]};
    assign in3387_2 = {s898[0]};
    Full_Adder FA_3387(s3387, c3387, in3387_1, in3387_2, s896[0]);
    wire[0:0] s3388, in3388_1, in3388_2;
    wire c3388;
    assign in3388_1 = {s900[0]};
    assign in3388_2 = {s901[0]};
    Full_Adder FA_3388(s3388, c3388, in3388_1, in3388_2, s899[0]);
    wire[0:0] s3389, in3389_1, in3389_2;
    wire c3389;
    assign in3389_1 = {pp127[1]};
    assign in3389_2 = {c862};
    Full_Adder FA_3389(s3389, c3389, in3389_1, in3389_2, pp126[2]);
    wire[0:0] s3390, in3390_1, in3390_2;
    wire c3390;
    assign in3390_1 = {c864};
    assign in3390_2 = {c865};
    Full_Adder FA_3390(s3390, c3390, in3390_1, in3390_2, c863);
    wire[0:0] s3391, in3391_1, in3391_2;
    wire c3391;
    assign in3391_1 = {c867};
    assign in3391_2 = {c868};
    Full_Adder FA_3391(s3391, c3391, in3391_1, in3391_2, c866);
    wire[0:0] s3392, in3392_1, in3392_2;
    wire c3392;
    assign in3392_1 = {c870};
    assign in3392_2 = {c871};
    Full_Adder FA_3392(s3392, c3392, in3392_1, in3392_2, c869);
    wire[0:0] s3393, in3393_1, in3393_2;
    wire c3393;
    assign in3393_1 = {c873};
    assign in3393_2 = {c874};
    Full_Adder FA_3393(s3393, c3393, in3393_1, in3393_2, c872);
    wire[0:0] s3394, in3394_1, in3394_2;
    wire c3394;
    assign in3394_1 = {c876};
    assign in3394_2 = {c877};
    Full_Adder FA_3394(s3394, c3394, in3394_1, in3394_2, c875);
    wire[0:0] s3395, in3395_1, in3395_2;
    wire c3395;
    assign in3395_1 = {c879};
    assign in3395_2 = {c880};
    Full_Adder FA_3395(s3395, c3395, in3395_1, in3395_2, c878);
    wire[0:0] s3396, in3396_1, in3396_2;
    wire c3396;
    assign in3396_1 = {c882};
    assign in3396_2 = {c883};
    Full_Adder FA_3396(s3396, c3396, in3396_1, in3396_2, c881);
    wire[0:0] s3397, in3397_1, in3397_2;
    wire c3397;
    assign in3397_1 = {c885};
    assign in3397_2 = {c886};
    Full_Adder FA_3397(s3397, c3397, in3397_1, in3397_2, c884);
    wire[0:0] s3398, in3398_1, in3398_2;
    wire c3398;
    assign in3398_1 = {c888};
    assign in3398_2 = {c889};
    Full_Adder FA_3398(s3398, c3398, in3398_1, in3398_2, c887);
    wire[0:0] s3399, in3399_1, in3399_2;
    wire c3399;
    assign in3399_1 = {c891};
    assign in3399_2 = {c892};
    Full_Adder FA_3399(s3399, c3399, in3399_1, in3399_2, c890);
    wire[0:0] s3400, in3400_1, in3400_2;
    wire c3400;
    assign in3400_1 = {c894};
    assign in3400_2 = {c895};
    Full_Adder FA_3400(s3400, c3400, in3400_1, in3400_2, c893);
    wire[0:0] s3401, in3401_1, in3401_2;
    wire c3401;
    assign in3401_1 = {c897};
    assign in3401_2 = {c898};
    Full_Adder FA_3401(s3401, c3401, in3401_1, in3401_2, c896);
    wire[0:0] s3402, in3402_1, in3402_2;
    wire c3402;
    assign in3402_1 = {c900};
    assign in3402_2 = {c901};
    Full_Adder FA_3402(s3402, c3402, in3402_1, in3402_2, c899);
    wire[0:0] s3403, in3403_1, in3403_2;
    wire c3403;
    assign in3403_1 = {c903};
    assign in3403_2 = {s904[0]};
    Full_Adder FA_3403(s3403, c3403, in3403_1, in3403_2, c902);
    wire[0:0] s3404, in3404_1, in3404_2;
    wire c3404;
    assign in3404_1 = {s906[0]};
    assign in3404_2 = {s907[0]};
    Full_Adder FA_3404(s3404, c3404, in3404_1, in3404_2, s905[0]);
    wire[0:0] s3405, in3405_1, in3405_2;
    wire c3405;
    assign in3405_1 = {s909[0]};
    assign in3405_2 = {s910[0]};
    Full_Adder FA_3405(s3405, c3405, in3405_1, in3405_2, s908[0]);
    wire[0:0] s3406, in3406_1, in3406_2;
    wire c3406;
    assign in3406_1 = {s912[0]};
    assign in3406_2 = {s913[0]};
    Full_Adder FA_3406(s3406, c3406, in3406_1, in3406_2, s911[0]);
    wire[0:0] s3407, in3407_1, in3407_2;
    wire c3407;
    assign in3407_1 = {s915[0]};
    assign in3407_2 = {s916[0]};
    Full_Adder FA_3407(s3407, c3407, in3407_1, in3407_2, s914[0]);
    wire[0:0] s3408, in3408_1, in3408_2;
    wire c3408;
    assign in3408_1 = {s918[0]};
    assign in3408_2 = {s919[0]};
    Full_Adder FA_3408(s3408, c3408, in3408_1, in3408_2, s917[0]);
    wire[0:0] s3409, in3409_1, in3409_2;
    wire c3409;
    assign in3409_1 = {s921[0]};
    assign in3409_2 = {s922[0]};
    Full_Adder FA_3409(s3409, c3409, in3409_1, in3409_2, s920[0]);
    wire[0:0] s3410, in3410_1, in3410_2;
    wire c3410;
    assign in3410_1 = {s924[0]};
    assign in3410_2 = {s925[0]};
    Full_Adder FA_3410(s3410, c3410, in3410_1, in3410_2, s923[0]);
    wire[0:0] s3411, in3411_1, in3411_2;
    wire c3411;
    assign in3411_1 = {s927[0]};
    assign in3411_2 = {s928[0]};
    Full_Adder FA_3411(s3411, c3411, in3411_1, in3411_2, s926[0]);
    wire[0:0] s3412, in3412_1, in3412_2;
    wire c3412;
    assign in3412_1 = {s930[0]};
    assign in3412_2 = {s931[0]};
    Full_Adder FA_3412(s3412, c3412, in3412_1, in3412_2, s929[0]);
    wire[0:0] s3413, in3413_1, in3413_2;
    wire c3413;
    assign in3413_1 = {s933[0]};
    assign in3413_2 = {s934[0]};
    Full_Adder FA_3413(s3413, c3413, in3413_1, in3413_2, s932[0]);
    wire[0:0] s3414, in3414_1, in3414_2;
    wire c3414;
    assign in3414_1 = {s936[0]};
    assign in3414_2 = {s937[0]};
    Full_Adder FA_3414(s3414, c3414, in3414_1, in3414_2, s935[0]);
    wire[0:0] s3415, in3415_1, in3415_2;
    wire c3415;
    assign in3415_1 = {s939[0]};
    assign in3415_2 = {s940[0]};
    Full_Adder FA_3415(s3415, c3415, in3415_1, in3415_2, s938[0]);
    wire[0:0] s3416, in3416_1, in3416_2;
    wire c3416;
    assign in3416_1 = {s942[0]};
    assign in3416_2 = {s943[0]};
    Full_Adder FA_3416(s3416, c3416, in3416_1, in3416_2, s941[0]);
    wire[0:0] s3417, in3417_1, in3417_2;
    wire c3417;
    assign in3417_1 = {pp126[3]};
    assign in3417_2 = {pp127[2]};
    Full_Adder FA_3417(s3417, c3417, in3417_1, in3417_2, pp125[4]);
    wire[0:0] s3418, in3418_1, in3418_2;
    wire c3418;
    assign in3418_1 = {c905};
    assign in3418_2 = {c906};
    Full_Adder FA_3418(s3418, c3418, in3418_1, in3418_2, c904);
    wire[0:0] s3419, in3419_1, in3419_2;
    wire c3419;
    assign in3419_1 = {c908};
    assign in3419_2 = {c909};
    Full_Adder FA_3419(s3419, c3419, in3419_1, in3419_2, c907);
    wire[0:0] s3420, in3420_1, in3420_2;
    wire c3420;
    assign in3420_1 = {c911};
    assign in3420_2 = {c912};
    Full_Adder FA_3420(s3420, c3420, in3420_1, in3420_2, c910);
    wire[0:0] s3421, in3421_1, in3421_2;
    wire c3421;
    assign in3421_1 = {c914};
    assign in3421_2 = {c915};
    Full_Adder FA_3421(s3421, c3421, in3421_1, in3421_2, c913);
    wire[0:0] s3422, in3422_1, in3422_2;
    wire c3422;
    assign in3422_1 = {c917};
    assign in3422_2 = {c918};
    Full_Adder FA_3422(s3422, c3422, in3422_1, in3422_2, c916);
    wire[0:0] s3423, in3423_1, in3423_2;
    wire c3423;
    assign in3423_1 = {c920};
    assign in3423_2 = {c921};
    Full_Adder FA_3423(s3423, c3423, in3423_1, in3423_2, c919);
    wire[0:0] s3424, in3424_1, in3424_2;
    wire c3424;
    assign in3424_1 = {c923};
    assign in3424_2 = {c924};
    Full_Adder FA_3424(s3424, c3424, in3424_1, in3424_2, c922);
    wire[0:0] s3425, in3425_1, in3425_2;
    wire c3425;
    assign in3425_1 = {c926};
    assign in3425_2 = {c927};
    Full_Adder FA_3425(s3425, c3425, in3425_1, in3425_2, c925);
    wire[0:0] s3426, in3426_1, in3426_2;
    wire c3426;
    assign in3426_1 = {c929};
    assign in3426_2 = {c930};
    Full_Adder FA_3426(s3426, c3426, in3426_1, in3426_2, c928);
    wire[0:0] s3427, in3427_1, in3427_2;
    wire c3427;
    assign in3427_1 = {c932};
    assign in3427_2 = {c933};
    Full_Adder FA_3427(s3427, c3427, in3427_1, in3427_2, c931);
    wire[0:0] s3428, in3428_1, in3428_2;
    wire c3428;
    assign in3428_1 = {c935};
    assign in3428_2 = {c936};
    Full_Adder FA_3428(s3428, c3428, in3428_1, in3428_2, c934);
    wire[0:0] s3429, in3429_1, in3429_2;
    wire c3429;
    assign in3429_1 = {c938};
    assign in3429_2 = {c939};
    Full_Adder FA_3429(s3429, c3429, in3429_1, in3429_2, c937);
    wire[0:0] s3430, in3430_1, in3430_2;
    wire c3430;
    assign in3430_1 = {c941};
    assign in3430_2 = {c942};
    Full_Adder FA_3430(s3430, c3430, in3430_1, in3430_2, c940);
    wire[0:0] s3431, in3431_1, in3431_2;
    wire c3431;
    assign in3431_1 = {c944};
    assign in3431_2 = {c945};
    Full_Adder FA_3431(s3431, c3431, in3431_1, in3431_2, c943);
    wire[0:0] s3432, in3432_1, in3432_2;
    wire c3432;
    assign in3432_1 = {s947[0]};
    assign in3432_2 = {s948[0]};
    Full_Adder FA_3432(s3432, c3432, in3432_1, in3432_2, s946[0]);
    wire[0:0] s3433, in3433_1, in3433_2;
    wire c3433;
    assign in3433_1 = {s950[0]};
    assign in3433_2 = {s951[0]};
    Full_Adder FA_3433(s3433, c3433, in3433_1, in3433_2, s949[0]);
    wire[0:0] s3434, in3434_1, in3434_2;
    wire c3434;
    assign in3434_1 = {s953[0]};
    assign in3434_2 = {s954[0]};
    Full_Adder FA_3434(s3434, c3434, in3434_1, in3434_2, s952[0]);
    wire[0:0] s3435, in3435_1, in3435_2;
    wire c3435;
    assign in3435_1 = {s956[0]};
    assign in3435_2 = {s957[0]};
    Full_Adder FA_3435(s3435, c3435, in3435_1, in3435_2, s955[0]);
    wire[0:0] s3436, in3436_1, in3436_2;
    wire c3436;
    assign in3436_1 = {s959[0]};
    assign in3436_2 = {s960[0]};
    Full_Adder FA_3436(s3436, c3436, in3436_1, in3436_2, s958[0]);
    wire[0:0] s3437, in3437_1, in3437_2;
    wire c3437;
    assign in3437_1 = {s962[0]};
    assign in3437_2 = {s963[0]};
    Full_Adder FA_3437(s3437, c3437, in3437_1, in3437_2, s961[0]);
    wire[0:0] s3438, in3438_1, in3438_2;
    wire c3438;
    assign in3438_1 = {s965[0]};
    assign in3438_2 = {s966[0]};
    Full_Adder FA_3438(s3438, c3438, in3438_1, in3438_2, s964[0]);
    wire[0:0] s3439, in3439_1, in3439_2;
    wire c3439;
    assign in3439_1 = {s968[0]};
    assign in3439_2 = {s969[0]};
    Full_Adder FA_3439(s3439, c3439, in3439_1, in3439_2, s967[0]);
    wire[0:0] s3440, in3440_1, in3440_2;
    wire c3440;
    assign in3440_1 = {s971[0]};
    assign in3440_2 = {s972[0]};
    Full_Adder FA_3440(s3440, c3440, in3440_1, in3440_2, s970[0]);
    wire[0:0] s3441, in3441_1, in3441_2;
    wire c3441;
    assign in3441_1 = {s974[0]};
    assign in3441_2 = {s975[0]};
    Full_Adder FA_3441(s3441, c3441, in3441_1, in3441_2, s973[0]);
    wire[0:0] s3442, in3442_1, in3442_2;
    wire c3442;
    assign in3442_1 = {s977[0]};
    assign in3442_2 = {s978[0]};
    Full_Adder FA_3442(s3442, c3442, in3442_1, in3442_2, s976[0]);
    wire[0:0] s3443, in3443_1, in3443_2;
    wire c3443;
    assign in3443_1 = {s980[0]};
    assign in3443_2 = {s981[0]};
    Full_Adder FA_3443(s3443, c3443, in3443_1, in3443_2, s979[0]);
    wire[0:0] s3444, in3444_1, in3444_2;
    wire c3444;
    assign in3444_1 = {s983[0]};
    assign in3444_2 = {s984[0]};
    Full_Adder FA_3444(s3444, c3444, in3444_1, in3444_2, s982[0]);
    wire[0:0] s3445, in3445_1, in3445_2;
    wire c3445;
    assign in3445_1 = {pp124[6]};
    assign in3445_2 = {pp125[5]};
    Full_Adder FA_3445(s3445, c3445, in3445_1, in3445_2, pp123[7]);
    wire[0:0] s3446, in3446_1, in3446_2;
    wire c3446;
    assign in3446_1 = {pp127[3]};
    assign in3446_2 = {c946};
    Full_Adder FA_3446(s3446, c3446, in3446_1, in3446_2, pp126[4]);
    wire[0:0] s3447, in3447_1, in3447_2;
    wire c3447;
    assign in3447_1 = {c948};
    assign in3447_2 = {c949};
    Full_Adder FA_3447(s3447, c3447, in3447_1, in3447_2, c947);
    wire[0:0] s3448, in3448_1, in3448_2;
    wire c3448;
    assign in3448_1 = {c951};
    assign in3448_2 = {c952};
    Full_Adder FA_3448(s3448, c3448, in3448_1, in3448_2, c950);
    wire[0:0] s3449, in3449_1, in3449_2;
    wire c3449;
    assign in3449_1 = {c954};
    assign in3449_2 = {c955};
    Full_Adder FA_3449(s3449, c3449, in3449_1, in3449_2, c953);
    wire[0:0] s3450, in3450_1, in3450_2;
    wire c3450;
    assign in3450_1 = {c957};
    assign in3450_2 = {c958};
    Full_Adder FA_3450(s3450, c3450, in3450_1, in3450_2, c956);
    wire[0:0] s3451, in3451_1, in3451_2;
    wire c3451;
    assign in3451_1 = {c960};
    assign in3451_2 = {c961};
    Full_Adder FA_3451(s3451, c3451, in3451_1, in3451_2, c959);
    wire[0:0] s3452, in3452_1, in3452_2;
    wire c3452;
    assign in3452_1 = {c963};
    assign in3452_2 = {c964};
    Full_Adder FA_3452(s3452, c3452, in3452_1, in3452_2, c962);
    wire[0:0] s3453, in3453_1, in3453_2;
    wire c3453;
    assign in3453_1 = {c966};
    assign in3453_2 = {c967};
    Full_Adder FA_3453(s3453, c3453, in3453_1, in3453_2, c965);
    wire[0:0] s3454, in3454_1, in3454_2;
    wire c3454;
    assign in3454_1 = {c969};
    assign in3454_2 = {c970};
    Full_Adder FA_3454(s3454, c3454, in3454_1, in3454_2, c968);
    wire[0:0] s3455, in3455_1, in3455_2;
    wire c3455;
    assign in3455_1 = {c972};
    assign in3455_2 = {c973};
    Full_Adder FA_3455(s3455, c3455, in3455_1, in3455_2, c971);
    wire[0:0] s3456, in3456_1, in3456_2;
    wire c3456;
    assign in3456_1 = {c975};
    assign in3456_2 = {c976};
    Full_Adder FA_3456(s3456, c3456, in3456_1, in3456_2, c974);
    wire[0:0] s3457, in3457_1, in3457_2;
    wire c3457;
    assign in3457_1 = {c978};
    assign in3457_2 = {c979};
    Full_Adder FA_3457(s3457, c3457, in3457_1, in3457_2, c977);
    wire[0:0] s3458, in3458_1, in3458_2;
    wire c3458;
    assign in3458_1 = {c981};
    assign in3458_2 = {c982};
    Full_Adder FA_3458(s3458, c3458, in3458_1, in3458_2, c980);
    wire[0:0] s3459, in3459_1, in3459_2;
    wire c3459;
    assign in3459_1 = {c984};
    assign in3459_2 = {c985};
    Full_Adder FA_3459(s3459, c3459, in3459_1, in3459_2, c983);
    wire[0:0] s3460, in3460_1, in3460_2;
    wire c3460;
    assign in3460_1 = {s987[0]};
    assign in3460_2 = {s988[0]};
    Full_Adder FA_3460(s3460, c3460, in3460_1, in3460_2, c986);
    wire[0:0] s3461, in3461_1, in3461_2;
    wire c3461;
    assign in3461_1 = {s990[0]};
    assign in3461_2 = {s991[0]};
    Full_Adder FA_3461(s3461, c3461, in3461_1, in3461_2, s989[0]);
    wire[0:0] s3462, in3462_1, in3462_2;
    wire c3462;
    assign in3462_1 = {s993[0]};
    assign in3462_2 = {s994[0]};
    Full_Adder FA_3462(s3462, c3462, in3462_1, in3462_2, s992[0]);
    wire[0:0] s3463, in3463_1, in3463_2;
    wire c3463;
    assign in3463_1 = {s996[0]};
    assign in3463_2 = {s997[0]};
    Full_Adder FA_3463(s3463, c3463, in3463_1, in3463_2, s995[0]);
    wire[0:0] s3464, in3464_1, in3464_2;
    wire c3464;
    assign in3464_1 = {s999[0]};
    assign in3464_2 = {s1000[0]};
    Full_Adder FA_3464(s3464, c3464, in3464_1, in3464_2, s998[0]);
    wire[0:0] s3465, in3465_1, in3465_2;
    wire c3465;
    assign in3465_1 = {s1002[0]};
    assign in3465_2 = {s1003[0]};
    Full_Adder FA_3465(s3465, c3465, in3465_1, in3465_2, s1001[0]);
    wire[0:0] s3466, in3466_1, in3466_2;
    wire c3466;
    assign in3466_1 = {s1005[0]};
    assign in3466_2 = {s1006[0]};
    Full_Adder FA_3466(s3466, c3466, in3466_1, in3466_2, s1004[0]);
    wire[0:0] s3467, in3467_1, in3467_2;
    wire c3467;
    assign in3467_1 = {s1008[0]};
    assign in3467_2 = {s1009[0]};
    Full_Adder FA_3467(s3467, c3467, in3467_1, in3467_2, s1007[0]);
    wire[0:0] s3468, in3468_1, in3468_2;
    wire c3468;
    assign in3468_1 = {s1011[0]};
    assign in3468_2 = {s1012[0]};
    Full_Adder FA_3468(s3468, c3468, in3468_1, in3468_2, s1010[0]);
    wire[0:0] s3469, in3469_1, in3469_2;
    wire c3469;
    assign in3469_1 = {s1014[0]};
    assign in3469_2 = {s1015[0]};
    Full_Adder FA_3469(s3469, c3469, in3469_1, in3469_2, s1013[0]);
    wire[0:0] s3470, in3470_1, in3470_2;
    wire c3470;
    assign in3470_1 = {s1017[0]};
    assign in3470_2 = {s1018[0]};
    Full_Adder FA_3470(s3470, c3470, in3470_1, in3470_2, s1016[0]);
    wire[0:0] s3471, in3471_1, in3471_2;
    wire c3471;
    assign in3471_1 = {s1020[0]};
    assign in3471_2 = {s1021[0]};
    Full_Adder FA_3471(s3471, c3471, in3471_1, in3471_2, s1019[0]);
    wire[0:0] s3472, in3472_1, in3472_2;
    wire c3472;
    assign in3472_1 = {s1023[0]};
    assign in3472_2 = {s1024[0]};
    Full_Adder FA_3472(s3472, c3472, in3472_1, in3472_2, s1022[0]);
    wire[0:0] s3473, in3473_1, in3473_2;
    wire c3473;
    assign in3473_1 = {pp122[9]};
    assign in3473_2 = {pp123[8]};
    Full_Adder FA_3473(s3473, c3473, in3473_1, in3473_2, pp121[10]);
    wire[0:0] s3474, in3474_1, in3474_2;
    wire c3474;
    assign in3474_1 = {pp125[6]};
    assign in3474_2 = {pp126[5]};
    Full_Adder FA_3474(s3474, c3474, in3474_1, in3474_2, pp124[7]);
    wire[0:0] s3475, in3475_1, in3475_2;
    wire c3475;
    assign in3475_1 = {c987};
    assign in3475_2 = {c988};
    Full_Adder FA_3475(s3475, c3475, in3475_1, in3475_2, pp127[4]);
    wire[0:0] s3476, in3476_1, in3476_2;
    wire c3476;
    assign in3476_1 = {c990};
    assign in3476_2 = {c991};
    Full_Adder FA_3476(s3476, c3476, in3476_1, in3476_2, c989);
    wire[0:0] s3477, in3477_1, in3477_2;
    wire c3477;
    assign in3477_1 = {c993};
    assign in3477_2 = {c994};
    Full_Adder FA_3477(s3477, c3477, in3477_1, in3477_2, c992);
    wire[0:0] s3478, in3478_1, in3478_2;
    wire c3478;
    assign in3478_1 = {c996};
    assign in3478_2 = {c997};
    Full_Adder FA_3478(s3478, c3478, in3478_1, in3478_2, c995);
    wire[0:0] s3479, in3479_1, in3479_2;
    wire c3479;
    assign in3479_1 = {c999};
    assign in3479_2 = {c1000};
    Full_Adder FA_3479(s3479, c3479, in3479_1, in3479_2, c998);
    wire[0:0] s3480, in3480_1, in3480_2;
    wire c3480;
    assign in3480_1 = {c1002};
    assign in3480_2 = {c1003};
    Full_Adder FA_3480(s3480, c3480, in3480_1, in3480_2, c1001);
    wire[0:0] s3481, in3481_1, in3481_2;
    wire c3481;
    assign in3481_1 = {c1005};
    assign in3481_2 = {c1006};
    Full_Adder FA_3481(s3481, c3481, in3481_1, in3481_2, c1004);
    wire[0:0] s3482, in3482_1, in3482_2;
    wire c3482;
    assign in3482_1 = {c1008};
    assign in3482_2 = {c1009};
    Full_Adder FA_3482(s3482, c3482, in3482_1, in3482_2, c1007);
    wire[0:0] s3483, in3483_1, in3483_2;
    wire c3483;
    assign in3483_1 = {c1011};
    assign in3483_2 = {c1012};
    Full_Adder FA_3483(s3483, c3483, in3483_1, in3483_2, c1010);
    wire[0:0] s3484, in3484_1, in3484_2;
    wire c3484;
    assign in3484_1 = {c1014};
    assign in3484_2 = {c1015};
    Full_Adder FA_3484(s3484, c3484, in3484_1, in3484_2, c1013);
    wire[0:0] s3485, in3485_1, in3485_2;
    wire c3485;
    assign in3485_1 = {c1017};
    assign in3485_2 = {c1018};
    Full_Adder FA_3485(s3485, c3485, in3485_1, in3485_2, c1016);
    wire[0:0] s3486, in3486_1, in3486_2;
    wire c3486;
    assign in3486_1 = {c1020};
    assign in3486_2 = {c1021};
    Full_Adder FA_3486(s3486, c3486, in3486_1, in3486_2, c1019);
    wire[0:0] s3487, in3487_1, in3487_2;
    wire c3487;
    assign in3487_1 = {c1023};
    assign in3487_2 = {c1024};
    Full_Adder FA_3487(s3487, c3487, in3487_1, in3487_2, c1022);
    wire[0:0] s3488, in3488_1, in3488_2;
    wire c3488;
    assign in3488_1 = {c1026};
    assign in3488_2 = {s1027[0]};
    Full_Adder FA_3488(s3488, c3488, in3488_1, in3488_2, c1025);
    wire[0:0] s3489, in3489_1, in3489_2;
    wire c3489;
    assign in3489_1 = {s1029[0]};
    assign in3489_2 = {s1030[0]};
    Full_Adder FA_3489(s3489, c3489, in3489_1, in3489_2, s1028[0]);
    wire[0:0] s3490, in3490_1, in3490_2;
    wire c3490;
    assign in3490_1 = {s1032[0]};
    assign in3490_2 = {s1033[0]};
    Full_Adder FA_3490(s3490, c3490, in3490_1, in3490_2, s1031[0]);
    wire[0:0] s3491, in3491_1, in3491_2;
    wire c3491;
    assign in3491_1 = {s1035[0]};
    assign in3491_2 = {s1036[0]};
    Full_Adder FA_3491(s3491, c3491, in3491_1, in3491_2, s1034[0]);
    wire[0:0] s3492, in3492_1, in3492_2;
    wire c3492;
    assign in3492_1 = {s1038[0]};
    assign in3492_2 = {s1039[0]};
    Full_Adder FA_3492(s3492, c3492, in3492_1, in3492_2, s1037[0]);
    wire[0:0] s3493, in3493_1, in3493_2;
    wire c3493;
    assign in3493_1 = {s1041[0]};
    assign in3493_2 = {s1042[0]};
    Full_Adder FA_3493(s3493, c3493, in3493_1, in3493_2, s1040[0]);
    wire[0:0] s3494, in3494_1, in3494_2;
    wire c3494;
    assign in3494_1 = {s1044[0]};
    assign in3494_2 = {s1045[0]};
    Full_Adder FA_3494(s3494, c3494, in3494_1, in3494_2, s1043[0]);
    wire[0:0] s3495, in3495_1, in3495_2;
    wire c3495;
    assign in3495_1 = {s1047[0]};
    assign in3495_2 = {s1048[0]};
    Full_Adder FA_3495(s3495, c3495, in3495_1, in3495_2, s1046[0]);
    wire[0:0] s3496, in3496_1, in3496_2;
    wire c3496;
    assign in3496_1 = {s1050[0]};
    assign in3496_2 = {s1051[0]};
    Full_Adder FA_3496(s3496, c3496, in3496_1, in3496_2, s1049[0]);
    wire[0:0] s3497, in3497_1, in3497_2;
    wire c3497;
    assign in3497_1 = {s1053[0]};
    assign in3497_2 = {s1054[0]};
    Full_Adder FA_3497(s3497, c3497, in3497_1, in3497_2, s1052[0]);
    wire[0:0] s3498, in3498_1, in3498_2;
    wire c3498;
    assign in3498_1 = {s1056[0]};
    assign in3498_2 = {s1057[0]};
    Full_Adder FA_3498(s3498, c3498, in3498_1, in3498_2, s1055[0]);
    wire[0:0] s3499, in3499_1, in3499_2;
    wire c3499;
    assign in3499_1 = {s1059[0]};
    assign in3499_2 = {s1060[0]};
    Full_Adder FA_3499(s3499, c3499, in3499_1, in3499_2, s1058[0]);
    wire[0:0] s3500, in3500_1, in3500_2;
    wire c3500;
    assign in3500_1 = {s1062[0]};
    assign in3500_2 = {s1063[0]};
    Full_Adder FA_3500(s3500, c3500, in3500_1, in3500_2, s1061[0]);
    wire[0:0] s3501, in3501_1, in3501_2;
    wire c3501;
    assign in3501_1 = {pp120[12]};
    assign in3501_2 = {pp121[11]};
    Full_Adder FA_3501(s3501, c3501, in3501_1, in3501_2, pp119[13]);
    wire[0:0] s3502, in3502_1, in3502_2;
    wire c3502;
    assign in3502_1 = {pp123[9]};
    assign in3502_2 = {pp124[8]};
    Full_Adder FA_3502(s3502, c3502, in3502_1, in3502_2, pp122[10]);
    wire[0:0] s3503, in3503_1, in3503_2;
    wire c3503;
    assign in3503_1 = {pp126[6]};
    assign in3503_2 = {pp127[5]};
    Full_Adder FA_3503(s3503, c3503, in3503_1, in3503_2, pp125[7]);
    wire[0:0] s3504, in3504_1, in3504_2;
    wire c3504;
    assign in3504_1 = {c1028};
    assign in3504_2 = {c1029};
    Full_Adder FA_3504(s3504, c3504, in3504_1, in3504_2, c1027);
    wire[0:0] s3505, in3505_1, in3505_2;
    wire c3505;
    assign in3505_1 = {c1031};
    assign in3505_2 = {c1032};
    Full_Adder FA_3505(s3505, c3505, in3505_1, in3505_2, c1030);
    wire[0:0] s3506, in3506_1, in3506_2;
    wire c3506;
    assign in3506_1 = {c1034};
    assign in3506_2 = {c1035};
    Full_Adder FA_3506(s3506, c3506, in3506_1, in3506_2, c1033);
    wire[0:0] s3507, in3507_1, in3507_2;
    wire c3507;
    assign in3507_1 = {c1037};
    assign in3507_2 = {c1038};
    Full_Adder FA_3507(s3507, c3507, in3507_1, in3507_2, c1036);
    wire[0:0] s3508, in3508_1, in3508_2;
    wire c3508;
    assign in3508_1 = {c1040};
    assign in3508_2 = {c1041};
    Full_Adder FA_3508(s3508, c3508, in3508_1, in3508_2, c1039);
    wire[0:0] s3509, in3509_1, in3509_2;
    wire c3509;
    assign in3509_1 = {c1043};
    assign in3509_2 = {c1044};
    Full_Adder FA_3509(s3509, c3509, in3509_1, in3509_2, c1042);
    wire[0:0] s3510, in3510_1, in3510_2;
    wire c3510;
    assign in3510_1 = {c1046};
    assign in3510_2 = {c1047};
    Full_Adder FA_3510(s3510, c3510, in3510_1, in3510_2, c1045);
    wire[0:0] s3511, in3511_1, in3511_2;
    wire c3511;
    assign in3511_1 = {c1049};
    assign in3511_2 = {c1050};
    Full_Adder FA_3511(s3511, c3511, in3511_1, in3511_2, c1048);
    wire[0:0] s3512, in3512_1, in3512_2;
    wire c3512;
    assign in3512_1 = {c1052};
    assign in3512_2 = {c1053};
    Full_Adder FA_3512(s3512, c3512, in3512_1, in3512_2, c1051);
    wire[0:0] s3513, in3513_1, in3513_2;
    wire c3513;
    assign in3513_1 = {c1055};
    assign in3513_2 = {c1056};
    Full_Adder FA_3513(s3513, c3513, in3513_1, in3513_2, c1054);
    wire[0:0] s3514, in3514_1, in3514_2;
    wire c3514;
    assign in3514_1 = {c1058};
    assign in3514_2 = {c1059};
    Full_Adder FA_3514(s3514, c3514, in3514_1, in3514_2, c1057);
    wire[0:0] s3515, in3515_1, in3515_2;
    wire c3515;
    assign in3515_1 = {c1061};
    assign in3515_2 = {c1062};
    Full_Adder FA_3515(s3515, c3515, in3515_1, in3515_2, c1060);
    wire[0:0] s3516, in3516_1, in3516_2;
    wire c3516;
    assign in3516_1 = {c1064};
    assign in3516_2 = {c1065};
    Full_Adder FA_3516(s3516, c3516, in3516_1, in3516_2, c1063);
    wire[0:0] s3517, in3517_1, in3517_2;
    wire c3517;
    assign in3517_1 = {s1067[0]};
    assign in3517_2 = {s1068[0]};
    Full_Adder FA_3517(s3517, c3517, in3517_1, in3517_2, s1066[0]);
    wire[0:0] s3518, in3518_1, in3518_2;
    wire c3518;
    assign in3518_1 = {s1070[0]};
    assign in3518_2 = {s1071[0]};
    Full_Adder FA_3518(s3518, c3518, in3518_1, in3518_2, s1069[0]);
    wire[0:0] s3519, in3519_1, in3519_2;
    wire c3519;
    assign in3519_1 = {s1073[0]};
    assign in3519_2 = {s1074[0]};
    Full_Adder FA_3519(s3519, c3519, in3519_1, in3519_2, s1072[0]);
    wire[0:0] s3520, in3520_1, in3520_2;
    wire c3520;
    assign in3520_1 = {s1076[0]};
    assign in3520_2 = {s1077[0]};
    Full_Adder FA_3520(s3520, c3520, in3520_1, in3520_2, s1075[0]);
    wire[0:0] s3521, in3521_1, in3521_2;
    wire c3521;
    assign in3521_1 = {s1079[0]};
    assign in3521_2 = {s1080[0]};
    Full_Adder FA_3521(s3521, c3521, in3521_1, in3521_2, s1078[0]);
    wire[0:0] s3522, in3522_1, in3522_2;
    wire c3522;
    assign in3522_1 = {s1082[0]};
    assign in3522_2 = {s1083[0]};
    Full_Adder FA_3522(s3522, c3522, in3522_1, in3522_2, s1081[0]);
    wire[0:0] s3523, in3523_1, in3523_2;
    wire c3523;
    assign in3523_1 = {s1085[0]};
    assign in3523_2 = {s1086[0]};
    Full_Adder FA_3523(s3523, c3523, in3523_1, in3523_2, s1084[0]);
    wire[0:0] s3524, in3524_1, in3524_2;
    wire c3524;
    assign in3524_1 = {s1088[0]};
    assign in3524_2 = {s1089[0]};
    Full_Adder FA_3524(s3524, c3524, in3524_1, in3524_2, s1087[0]);
    wire[0:0] s3525, in3525_1, in3525_2;
    wire c3525;
    assign in3525_1 = {s1091[0]};
    assign in3525_2 = {s1092[0]};
    Full_Adder FA_3525(s3525, c3525, in3525_1, in3525_2, s1090[0]);
    wire[0:0] s3526, in3526_1, in3526_2;
    wire c3526;
    assign in3526_1 = {s1094[0]};
    assign in3526_2 = {s1095[0]};
    Full_Adder FA_3526(s3526, c3526, in3526_1, in3526_2, s1093[0]);
    wire[0:0] s3527, in3527_1, in3527_2;
    wire c3527;
    assign in3527_1 = {s1097[0]};
    assign in3527_2 = {s1098[0]};
    Full_Adder FA_3527(s3527, c3527, in3527_1, in3527_2, s1096[0]);
    wire[0:0] s3528, in3528_1, in3528_2;
    wire c3528;
    assign in3528_1 = {s1100[0]};
    assign in3528_2 = {s1101[0]};
    Full_Adder FA_3528(s3528, c3528, in3528_1, in3528_2, s1099[0]);
    wire[0:0] s3529, in3529_1, in3529_2;
    wire c3529;
    assign in3529_1 = {pp118[15]};
    assign in3529_2 = {pp119[14]};
    Full_Adder FA_3529(s3529, c3529, in3529_1, in3529_2, pp117[16]);
    wire[0:0] s3530, in3530_1, in3530_2;
    wire c3530;
    assign in3530_1 = {pp121[12]};
    assign in3530_2 = {pp122[11]};
    Full_Adder FA_3530(s3530, c3530, in3530_1, in3530_2, pp120[13]);
    wire[0:0] s3531, in3531_1, in3531_2;
    wire c3531;
    assign in3531_1 = {pp124[9]};
    assign in3531_2 = {pp125[8]};
    Full_Adder FA_3531(s3531, c3531, in3531_1, in3531_2, pp123[10]);
    wire[0:0] s3532, in3532_1, in3532_2;
    wire c3532;
    assign in3532_1 = {pp127[6]};
    assign in3532_2 = {c1066};
    Full_Adder FA_3532(s3532, c3532, in3532_1, in3532_2, pp126[7]);
    wire[0:0] s3533, in3533_1, in3533_2;
    wire c3533;
    assign in3533_1 = {c1068};
    assign in3533_2 = {c1069};
    Full_Adder FA_3533(s3533, c3533, in3533_1, in3533_2, c1067);
    wire[0:0] s3534, in3534_1, in3534_2;
    wire c3534;
    assign in3534_1 = {c1071};
    assign in3534_2 = {c1072};
    Full_Adder FA_3534(s3534, c3534, in3534_1, in3534_2, c1070);
    wire[0:0] s3535, in3535_1, in3535_2;
    wire c3535;
    assign in3535_1 = {c1074};
    assign in3535_2 = {c1075};
    Full_Adder FA_3535(s3535, c3535, in3535_1, in3535_2, c1073);
    wire[0:0] s3536, in3536_1, in3536_2;
    wire c3536;
    assign in3536_1 = {c1077};
    assign in3536_2 = {c1078};
    Full_Adder FA_3536(s3536, c3536, in3536_1, in3536_2, c1076);
    wire[0:0] s3537, in3537_1, in3537_2;
    wire c3537;
    assign in3537_1 = {c1080};
    assign in3537_2 = {c1081};
    Full_Adder FA_3537(s3537, c3537, in3537_1, in3537_2, c1079);
    wire[0:0] s3538, in3538_1, in3538_2;
    wire c3538;
    assign in3538_1 = {c1083};
    assign in3538_2 = {c1084};
    Full_Adder FA_3538(s3538, c3538, in3538_1, in3538_2, c1082);
    wire[0:0] s3539, in3539_1, in3539_2;
    wire c3539;
    assign in3539_1 = {c1086};
    assign in3539_2 = {c1087};
    Full_Adder FA_3539(s3539, c3539, in3539_1, in3539_2, c1085);
    wire[0:0] s3540, in3540_1, in3540_2;
    wire c3540;
    assign in3540_1 = {c1089};
    assign in3540_2 = {c1090};
    Full_Adder FA_3540(s3540, c3540, in3540_1, in3540_2, c1088);
    wire[0:0] s3541, in3541_1, in3541_2;
    wire c3541;
    assign in3541_1 = {c1092};
    assign in3541_2 = {c1093};
    Full_Adder FA_3541(s3541, c3541, in3541_1, in3541_2, c1091);
    wire[0:0] s3542, in3542_1, in3542_2;
    wire c3542;
    assign in3542_1 = {c1095};
    assign in3542_2 = {c1096};
    Full_Adder FA_3542(s3542, c3542, in3542_1, in3542_2, c1094);
    wire[0:0] s3543, in3543_1, in3543_2;
    wire c3543;
    assign in3543_1 = {c1098};
    assign in3543_2 = {c1099};
    Full_Adder FA_3543(s3543, c3543, in3543_1, in3543_2, c1097);
    wire[0:0] s3544, in3544_1, in3544_2;
    wire c3544;
    assign in3544_1 = {c1101};
    assign in3544_2 = {c1102};
    Full_Adder FA_3544(s3544, c3544, in3544_1, in3544_2, c1100);
    wire[0:0] s3545, in3545_1, in3545_2;
    wire c3545;
    assign in3545_1 = {s1104[0]};
    assign in3545_2 = {s1105[0]};
    Full_Adder FA_3545(s3545, c3545, in3545_1, in3545_2, c1103);
    wire[0:0] s3546, in3546_1, in3546_2;
    wire c3546;
    assign in3546_1 = {s1107[0]};
    assign in3546_2 = {s1108[0]};
    Full_Adder FA_3546(s3546, c3546, in3546_1, in3546_2, s1106[0]);
    wire[0:0] s3547, in3547_1, in3547_2;
    wire c3547;
    assign in3547_1 = {s1110[0]};
    assign in3547_2 = {s1111[0]};
    Full_Adder FA_3547(s3547, c3547, in3547_1, in3547_2, s1109[0]);
    wire[0:0] s3548, in3548_1, in3548_2;
    wire c3548;
    assign in3548_1 = {s1113[0]};
    assign in3548_2 = {s1114[0]};
    Full_Adder FA_3548(s3548, c3548, in3548_1, in3548_2, s1112[0]);
    wire[0:0] s3549, in3549_1, in3549_2;
    wire c3549;
    assign in3549_1 = {s1116[0]};
    assign in3549_2 = {s1117[0]};
    Full_Adder FA_3549(s3549, c3549, in3549_1, in3549_2, s1115[0]);
    wire[0:0] s3550, in3550_1, in3550_2;
    wire c3550;
    assign in3550_1 = {s1119[0]};
    assign in3550_2 = {s1120[0]};
    Full_Adder FA_3550(s3550, c3550, in3550_1, in3550_2, s1118[0]);
    wire[0:0] s3551, in3551_1, in3551_2;
    wire c3551;
    assign in3551_1 = {s1122[0]};
    assign in3551_2 = {s1123[0]};
    Full_Adder FA_3551(s3551, c3551, in3551_1, in3551_2, s1121[0]);
    wire[0:0] s3552, in3552_1, in3552_2;
    wire c3552;
    assign in3552_1 = {s1125[0]};
    assign in3552_2 = {s1126[0]};
    Full_Adder FA_3552(s3552, c3552, in3552_1, in3552_2, s1124[0]);
    wire[0:0] s3553, in3553_1, in3553_2;
    wire c3553;
    assign in3553_1 = {s1128[0]};
    assign in3553_2 = {s1129[0]};
    Full_Adder FA_3553(s3553, c3553, in3553_1, in3553_2, s1127[0]);
    wire[0:0] s3554, in3554_1, in3554_2;
    wire c3554;
    assign in3554_1 = {s1131[0]};
    assign in3554_2 = {s1132[0]};
    Full_Adder FA_3554(s3554, c3554, in3554_1, in3554_2, s1130[0]);
    wire[0:0] s3555, in3555_1, in3555_2;
    wire c3555;
    assign in3555_1 = {s1134[0]};
    assign in3555_2 = {s1135[0]};
    Full_Adder FA_3555(s3555, c3555, in3555_1, in3555_2, s1133[0]);
    wire[0:0] s3556, in3556_1, in3556_2;
    wire c3556;
    assign in3556_1 = {s1137[0]};
    assign in3556_2 = {s1138[0]};
    Full_Adder FA_3556(s3556, c3556, in3556_1, in3556_2, s1136[0]);
    wire[0:0] s3557, in3557_1, in3557_2;
    wire c3557;
    assign in3557_1 = {pp116[18]};
    assign in3557_2 = {pp117[17]};
    Full_Adder FA_3557(s3557, c3557, in3557_1, in3557_2, pp115[19]);
    wire[0:0] s3558, in3558_1, in3558_2;
    wire c3558;
    assign in3558_1 = {pp119[15]};
    assign in3558_2 = {pp120[14]};
    Full_Adder FA_3558(s3558, c3558, in3558_1, in3558_2, pp118[16]);
    wire[0:0] s3559, in3559_1, in3559_2;
    wire c3559;
    assign in3559_1 = {pp122[12]};
    assign in3559_2 = {pp123[11]};
    Full_Adder FA_3559(s3559, c3559, in3559_1, in3559_2, pp121[13]);
    wire[0:0] s3560, in3560_1, in3560_2;
    wire c3560;
    assign in3560_1 = {pp125[9]};
    assign in3560_2 = {pp126[8]};
    Full_Adder FA_3560(s3560, c3560, in3560_1, in3560_2, pp124[10]);
    wire[0:0] s3561, in3561_1, in3561_2;
    wire c3561;
    assign in3561_1 = {c1104};
    assign in3561_2 = {c1105};
    Full_Adder FA_3561(s3561, c3561, in3561_1, in3561_2, pp127[7]);
    wire[0:0] s3562, in3562_1, in3562_2;
    wire c3562;
    assign in3562_1 = {c1107};
    assign in3562_2 = {c1108};
    Full_Adder FA_3562(s3562, c3562, in3562_1, in3562_2, c1106);
    wire[0:0] s3563, in3563_1, in3563_2;
    wire c3563;
    assign in3563_1 = {c1110};
    assign in3563_2 = {c1111};
    Full_Adder FA_3563(s3563, c3563, in3563_1, in3563_2, c1109);
    wire[0:0] s3564, in3564_1, in3564_2;
    wire c3564;
    assign in3564_1 = {c1113};
    assign in3564_2 = {c1114};
    Full_Adder FA_3564(s3564, c3564, in3564_1, in3564_2, c1112);
    wire[0:0] s3565, in3565_1, in3565_2;
    wire c3565;
    assign in3565_1 = {c1116};
    assign in3565_2 = {c1117};
    Full_Adder FA_3565(s3565, c3565, in3565_1, in3565_2, c1115);
    wire[0:0] s3566, in3566_1, in3566_2;
    wire c3566;
    assign in3566_1 = {c1119};
    assign in3566_2 = {c1120};
    Full_Adder FA_3566(s3566, c3566, in3566_1, in3566_2, c1118);
    wire[0:0] s3567, in3567_1, in3567_2;
    wire c3567;
    assign in3567_1 = {c1122};
    assign in3567_2 = {c1123};
    Full_Adder FA_3567(s3567, c3567, in3567_1, in3567_2, c1121);
    wire[0:0] s3568, in3568_1, in3568_2;
    wire c3568;
    assign in3568_1 = {c1125};
    assign in3568_2 = {c1126};
    Full_Adder FA_3568(s3568, c3568, in3568_1, in3568_2, c1124);
    wire[0:0] s3569, in3569_1, in3569_2;
    wire c3569;
    assign in3569_1 = {c1128};
    assign in3569_2 = {c1129};
    Full_Adder FA_3569(s3569, c3569, in3569_1, in3569_2, c1127);
    wire[0:0] s3570, in3570_1, in3570_2;
    wire c3570;
    assign in3570_1 = {c1131};
    assign in3570_2 = {c1132};
    Full_Adder FA_3570(s3570, c3570, in3570_1, in3570_2, c1130);
    wire[0:0] s3571, in3571_1, in3571_2;
    wire c3571;
    assign in3571_1 = {c1134};
    assign in3571_2 = {c1135};
    Full_Adder FA_3571(s3571, c3571, in3571_1, in3571_2, c1133);
    wire[0:0] s3572, in3572_1, in3572_2;
    wire c3572;
    assign in3572_1 = {c1137};
    assign in3572_2 = {c1138};
    Full_Adder FA_3572(s3572, c3572, in3572_1, in3572_2, c1136);
    wire[0:0] s3573, in3573_1, in3573_2;
    wire c3573;
    assign in3573_1 = {c1140};
    assign in3573_2 = {s1141[0]};
    Full_Adder FA_3573(s3573, c3573, in3573_1, in3573_2, c1139);
    wire[0:0] s3574, in3574_1, in3574_2;
    wire c3574;
    assign in3574_1 = {s1143[0]};
    assign in3574_2 = {s1144[0]};
    Full_Adder FA_3574(s3574, c3574, in3574_1, in3574_2, s1142[0]);
    wire[0:0] s3575, in3575_1, in3575_2;
    wire c3575;
    assign in3575_1 = {s1146[0]};
    assign in3575_2 = {s1147[0]};
    Full_Adder FA_3575(s3575, c3575, in3575_1, in3575_2, s1145[0]);
    wire[0:0] s3576, in3576_1, in3576_2;
    wire c3576;
    assign in3576_1 = {s1149[0]};
    assign in3576_2 = {s1150[0]};
    Full_Adder FA_3576(s3576, c3576, in3576_1, in3576_2, s1148[0]);
    wire[0:0] s3577, in3577_1, in3577_2;
    wire c3577;
    assign in3577_1 = {s1152[0]};
    assign in3577_2 = {s1153[0]};
    Full_Adder FA_3577(s3577, c3577, in3577_1, in3577_2, s1151[0]);
    wire[0:0] s3578, in3578_1, in3578_2;
    wire c3578;
    assign in3578_1 = {s1155[0]};
    assign in3578_2 = {s1156[0]};
    Full_Adder FA_3578(s3578, c3578, in3578_1, in3578_2, s1154[0]);
    wire[0:0] s3579, in3579_1, in3579_2;
    wire c3579;
    assign in3579_1 = {s1158[0]};
    assign in3579_2 = {s1159[0]};
    Full_Adder FA_3579(s3579, c3579, in3579_1, in3579_2, s1157[0]);
    wire[0:0] s3580, in3580_1, in3580_2;
    wire c3580;
    assign in3580_1 = {s1161[0]};
    assign in3580_2 = {s1162[0]};
    Full_Adder FA_3580(s3580, c3580, in3580_1, in3580_2, s1160[0]);
    wire[0:0] s3581, in3581_1, in3581_2;
    wire c3581;
    assign in3581_1 = {s1164[0]};
    assign in3581_2 = {s1165[0]};
    Full_Adder FA_3581(s3581, c3581, in3581_1, in3581_2, s1163[0]);
    wire[0:0] s3582, in3582_1, in3582_2;
    wire c3582;
    assign in3582_1 = {s1167[0]};
    assign in3582_2 = {s1168[0]};
    Full_Adder FA_3582(s3582, c3582, in3582_1, in3582_2, s1166[0]);
    wire[0:0] s3583, in3583_1, in3583_2;
    wire c3583;
    assign in3583_1 = {s1170[0]};
    assign in3583_2 = {s1171[0]};
    Full_Adder FA_3583(s3583, c3583, in3583_1, in3583_2, s1169[0]);
    wire[0:0] s3584, in3584_1, in3584_2;
    wire c3584;
    assign in3584_1 = {s1173[0]};
    assign in3584_2 = {s1174[0]};
    Full_Adder FA_3584(s3584, c3584, in3584_1, in3584_2, s1172[0]);
    wire[0:0] s3585, in3585_1, in3585_2;
    wire c3585;
    assign in3585_1 = {pp114[21]};
    assign in3585_2 = {pp115[20]};
    Full_Adder FA_3585(s3585, c3585, in3585_1, in3585_2, pp113[22]);
    wire[0:0] s3586, in3586_1, in3586_2;
    wire c3586;
    assign in3586_1 = {pp117[18]};
    assign in3586_2 = {pp118[17]};
    Full_Adder FA_3586(s3586, c3586, in3586_1, in3586_2, pp116[19]);
    wire[0:0] s3587, in3587_1, in3587_2;
    wire c3587;
    assign in3587_1 = {pp120[15]};
    assign in3587_2 = {pp121[14]};
    Full_Adder FA_3587(s3587, c3587, in3587_1, in3587_2, pp119[16]);
    wire[0:0] s3588, in3588_1, in3588_2;
    wire c3588;
    assign in3588_1 = {pp123[12]};
    assign in3588_2 = {pp124[11]};
    Full_Adder FA_3588(s3588, c3588, in3588_1, in3588_2, pp122[13]);
    wire[0:0] s3589, in3589_1, in3589_2;
    wire c3589;
    assign in3589_1 = {pp126[9]};
    assign in3589_2 = {pp127[8]};
    Full_Adder FA_3589(s3589, c3589, in3589_1, in3589_2, pp125[10]);
    wire[0:0] s3590, in3590_1, in3590_2;
    wire c3590;
    assign in3590_1 = {c1142};
    assign in3590_2 = {c1143};
    Full_Adder FA_3590(s3590, c3590, in3590_1, in3590_2, c1141);
    wire[0:0] s3591, in3591_1, in3591_2;
    wire c3591;
    assign in3591_1 = {c1145};
    assign in3591_2 = {c1146};
    Full_Adder FA_3591(s3591, c3591, in3591_1, in3591_2, c1144);
    wire[0:0] s3592, in3592_1, in3592_2;
    wire c3592;
    assign in3592_1 = {c1148};
    assign in3592_2 = {c1149};
    Full_Adder FA_3592(s3592, c3592, in3592_1, in3592_2, c1147);
    wire[0:0] s3593, in3593_1, in3593_2;
    wire c3593;
    assign in3593_1 = {c1151};
    assign in3593_2 = {c1152};
    Full_Adder FA_3593(s3593, c3593, in3593_1, in3593_2, c1150);
    wire[0:0] s3594, in3594_1, in3594_2;
    wire c3594;
    assign in3594_1 = {c1154};
    assign in3594_2 = {c1155};
    Full_Adder FA_3594(s3594, c3594, in3594_1, in3594_2, c1153);
    wire[0:0] s3595, in3595_1, in3595_2;
    wire c3595;
    assign in3595_1 = {c1157};
    assign in3595_2 = {c1158};
    Full_Adder FA_3595(s3595, c3595, in3595_1, in3595_2, c1156);
    wire[0:0] s3596, in3596_1, in3596_2;
    wire c3596;
    assign in3596_1 = {c1160};
    assign in3596_2 = {c1161};
    Full_Adder FA_3596(s3596, c3596, in3596_1, in3596_2, c1159);
    wire[0:0] s3597, in3597_1, in3597_2;
    wire c3597;
    assign in3597_1 = {c1163};
    assign in3597_2 = {c1164};
    Full_Adder FA_3597(s3597, c3597, in3597_1, in3597_2, c1162);
    wire[0:0] s3598, in3598_1, in3598_2;
    wire c3598;
    assign in3598_1 = {c1166};
    assign in3598_2 = {c1167};
    Full_Adder FA_3598(s3598, c3598, in3598_1, in3598_2, c1165);
    wire[0:0] s3599, in3599_1, in3599_2;
    wire c3599;
    assign in3599_1 = {c1169};
    assign in3599_2 = {c1170};
    Full_Adder FA_3599(s3599, c3599, in3599_1, in3599_2, c1168);
    wire[0:0] s3600, in3600_1, in3600_2;
    wire c3600;
    assign in3600_1 = {c1172};
    assign in3600_2 = {c1173};
    Full_Adder FA_3600(s3600, c3600, in3600_1, in3600_2, c1171);
    wire[0:0] s3601, in3601_1, in3601_2;
    wire c3601;
    assign in3601_1 = {c1175};
    assign in3601_2 = {c1176};
    Full_Adder FA_3601(s3601, c3601, in3601_1, in3601_2, c1174);
    wire[0:0] s3602, in3602_1, in3602_2;
    wire c3602;
    assign in3602_1 = {s1178[0]};
    assign in3602_2 = {s1179[0]};
    Full_Adder FA_3602(s3602, c3602, in3602_1, in3602_2, s1177[0]);
    wire[0:0] s3603, in3603_1, in3603_2;
    wire c3603;
    assign in3603_1 = {s1181[0]};
    assign in3603_2 = {s1182[0]};
    Full_Adder FA_3603(s3603, c3603, in3603_1, in3603_2, s1180[0]);
    wire[0:0] s3604, in3604_1, in3604_2;
    wire c3604;
    assign in3604_1 = {s1184[0]};
    assign in3604_2 = {s1185[0]};
    Full_Adder FA_3604(s3604, c3604, in3604_1, in3604_2, s1183[0]);
    wire[0:0] s3605, in3605_1, in3605_2;
    wire c3605;
    assign in3605_1 = {s1187[0]};
    assign in3605_2 = {s1188[0]};
    Full_Adder FA_3605(s3605, c3605, in3605_1, in3605_2, s1186[0]);
    wire[0:0] s3606, in3606_1, in3606_2;
    wire c3606;
    assign in3606_1 = {s1190[0]};
    assign in3606_2 = {s1191[0]};
    Full_Adder FA_3606(s3606, c3606, in3606_1, in3606_2, s1189[0]);
    wire[0:0] s3607, in3607_1, in3607_2;
    wire c3607;
    assign in3607_1 = {s1193[0]};
    assign in3607_2 = {s1194[0]};
    Full_Adder FA_3607(s3607, c3607, in3607_1, in3607_2, s1192[0]);
    wire[0:0] s3608, in3608_1, in3608_2;
    wire c3608;
    assign in3608_1 = {s1196[0]};
    assign in3608_2 = {s1197[0]};
    Full_Adder FA_3608(s3608, c3608, in3608_1, in3608_2, s1195[0]);
    wire[0:0] s3609, in3609_1, in3609_2;
    wire c3609;
    assign in3609_1 = {s1199[0]};
    assign in3609_2 = {s1200[0]};
    Full_Adder FA_3609(s3609, c3609, in3609_1, in3609_2, s1198[0]);
    wire[0:0] s3610, in3610_1, in3610_2;
    wire c3610;
    assign in3610_1 = {s1202[0]};
    assign in3610_2 = {s1203[0]};
    Full_Adder FA_3610(s3610, c3610, in3610_1, in3610_2, s1201[0]);
    wire[0:0] s3611, in3611_1, in3611_2;
    wire c3611;
    assign in3611_1 = {s1205[0]};
    assign in3611_2 = {s1206[0]};
    Full_Adder FA_3611(s3611, c3611, in3611_1, in3611_2, s1204[0]);
    wire[0:0] s3612, in3612_1, in3612_2;
    wire c3612;
    assign in3612_1 = {s1208[0]};
    assign in3612_2 = {s1209[0]};
    Full_Adder FA_3612(s3612, c3612, in3612_1, in3612_2, s1207[0]);
    wire[0:0] s3613, in3613_1, in3613_2;
    wire c3613;
    assign in3613_1 = {pp112[24]};
    assign in3613_2 = {pp113[23]};
    Full_Adder FA_3613(s3613, c3613, in3613_1, in3613_2, pp111[25]);
    wire[0:0] s3614, in3614_1, in3614_2;
    wire c3614;
    assign in3614_1 = {pp115[21]};
    assign in3614_2 = {pp116[20]};
    Full_Adder FA_3614(s3614, c3614, in3614_1, in3614_2, pp114[22]);
    wire[0:0] s3615, in3615_1, in3615_2;
    wire c3615;
    assign in3615_1 = {pp118[18]};
    assign in3615_2 = {pp119[17]};
    Full_Adder FA_3615(s3615, c3615, in3615_1, in3615_2, pp117[19]);
    wire[0:0] s3616, in3616_1, in3616_2;
    wire c3616;
    assign in3616_1 = {pp121[15]};
    assign in3616_2 = {pp122[14]};
    Full_Adder FA_3616(s3616, c3616, in3616_1, in3616_2, pp120[16]);
    wire[0:0] s3617, in3617_1, in3617_2;
    wire c3617;
    assign in3617_1 = {pp124[12]};
    assign in3617_2 = {pp125[11]};
    Full_Adder FA_3617(s3617, c3617, in3617_1, in3617_2, pp123[13]);
    wire[0:0] s3618, in3618_1, in3618_2;
    wire c3618;
    assign in3618_1 = {pp127[9]};
    assign in3618_2 = {c1177};
    Full_Adder FA_3618(s3618, c3618, in3618_1, in3618_2, pp126[10]);
    wire[0:0] s3619, in3619_1, in3619_2;
    wire c3619;
    assign in3619_1 = {c1179};
    assign in3619_2 = {c1180};
    Full_Adder FA_3619(s3619, c3619, in3619_1, in3619_2, c1178);
    wire[0:0] s3620, in3620_1, in3620_2;
    wire c3620;
    assign in3620_1 = {c1182};
    assign in3620_2 = {c1183};
    Full_Adder FA_3620(s3620, c3620, in3620_1, in3620_2, c1181);
    wire[0:0] s3621, in3621_1, in3621_2;
    wire c3621;
    assign in3621_1 = {c1185};
    assign in3621_2 = {c1186};
    Full_Adder FA_3621(s3621, c3621, in3621_1, in3621_2, c1184);
    wire[0:0] s3622, in3622_1, in3622_2;
    wire c3622;
    assign in3622_1 = {c1188};
    assign in3622_2 = {c1189};
    Full_Adder FA_3622(s3622, c3622, in3622_1, in3622_2, c1187);
    wire[0:0] s3623, in3623_1, in3623_2;
    wire c3623;
    assign in3623_1 = {c1191};
    assign in3623_2 = {c1192};
    Full_Adder FA_3623(s3623, c3623, in3623_1, in3623_2, c1190);
    wire[0:0] s3624, in3624_1, in3624_2;
    wire c3624;
    assign in3624_1 = {c1194};
    assign in3624_2 = {c1195};
    Full_Adder FA_3624(s3624, c3624, in3624_1, in3624_2, c1193);
    wire[0:0] s3625, in3625_1, in3625_2;
    wire c3625;
    assign in3625_1 = {c1197};
    assign in3625_2 = {c1198};
    Full_Adder FA_3625(s3625, c3625, in3625_1, in3625_2, c1196);
    wire[0:0] s3626, in3626_1, in3626_2;
    wire c3626;
    assign in3626_1 = {c1200};
    assign in3626_2 = {c1201};
    Full_Adder FA_3626(s3626, c3626, in3626_1, in3626_2, c1199);
    wire[0:0] s3627, in3627_1, in3627_2;
    wire c3627;
    assign in3627_1 = {c1203};
    assign in3627_2 = {c1204};
    Full_Adder FA_3627(s3627, c3627, in3627_1, in3627_2, c1202);
    wire[0:0] s3628, in3628_1, in3628_2;
    wire c3628;
    assign in3628_1 = {c1206};
    assign in3628_2 = {c1207};
    Full_Adder FA_3628(s3628, c3628, in3628_1, in3628_2, c1205);
    wire[0:0] s3629, in3629_1, in3629_2;
    wire c3629;
    assign in3629_1 = {c1209};
    assign in3629_2 = {c1210};
    Full_Adder FA_3629(s3629, c3629, in3629_1, in3629_2, c1208);
    wire[0:0] s3630, in3630_1, in3630_2;
    wire c3630;
    assign in3630_1 = {s1212[0]};
    assign in3630_2 = {s1213[0]};
    Full_Adder FA_3630(s3630, c3630, in3630_1, in3630_2, c1211);
    wire[0:0] s3631, in3631_1, in3631_2;
    wire c3631;
    assign in3631_1 = {s1215[0]};
    assign in3631_2 = {s1216[0]};
    Full_Adder FA_3631(s3631, c3631, in3631_1, in3631_2, s1214[0]);
    wire[0:0] s3632, in3632_1, in3632_2;
    wire c3632;
    assign in3632_1 = {s1218[0]};
    assign in3632_2 = {s1219[0]};
    Full_Adder FA_3632(s3632, c3632, in3632_1, in3632_2, s1217[0]);
    wire[0:0] s3633, in3633_1, in3633_2;
    wire c3633;
    assign in3633_1 = {s1221[0]};
    assign in3633_2 = {s1222[0]};
    Full_Adder FA_3633(s3633, c3633, in3633_1, in3633_2, s1220[0]);
    wire[0:0] s3634, in3634_1, in3634_2;
    wire c3634;
    assign in3634_1 = {s1224[0]};
    assign in3634_2 = {s1225[0]};
    Full_Adder FA_3634(s3634, c3634, in3634_1, in3634_2, s1223[0]);
    wire[0:0] s3635, in3635_1, in3635_2;
    wire c3635;
    assign in3635_1 = {s1227[0]};
    assign in3635_2 = {s1228[0]};
    Full_Adder FA_3635(s3635, c3635, in3635_1, in3635_2, s1226[0]);
    wire[0:0] s3636, in3636_1, in3636_2;
    wire c3636;
    assign in3636_1 = {s1230[0]};
    assign in3636_2 = {s1231[0]};
    Full_Adder FA_3636(s3636, c3636, in3636_1, in3636_2, s1229[0]);
    wire[0:0] s3637, in3637_1, in3637_2;
    wire c3637;
    assign in3637_1 = {s1233[0]};
    assign in3637_2 = {s1234[0]};
    Full_Adder FA_3637(s3637, c3637, in3637_1, in3637_2, s1232[0]);
    wire[0:0] s3638, in3638_1, in3638_2;
    wire c3638;
    assign in3638_1 = {s1236[0]};
    assign in3638_2 = {s1237[0]};
    Full_Adder FA_3638(s3638, c3638, in3638_1, in3638_2, s1235[0]);
    wire[0:0] s3639, in3639_1, in3639_2;
    wire c3639;
    assign in3639_1 = {s1239[0]};
    assign in3639_2 = {s1240[0]};
    Full_Adder FA_3639(s3639, c3639, in3639_1, in3639_2, s1238[0]);
    wire[0:0] s3640, in3640_1, in3640_2;
    wire c3640;
    assign in3640_1 = {s1242[0]};
    assign in3640_2 = {s1243[0]};
    Full_Adder FA_3640(s3640, c3640, in3640_1, in3640_2, s1241[0]);
    wire[0:0] s3641, in3641_1, in3641_2;
    wire c3641;
    assign in3641_1 = {pp110[27]};
    assign in3641_2 = {pp111[26]};
    Full_Adder FA_3641(s3641, c3641, in3641_1, in3641_2, pp109[28]);
    wire[0:0] s3642, in3642_1, in3642_2;
    wire c3642;
    assign in3642_1 = {pp113[24]};
    assign in3642_2 = {pp114[23]};
    Full_Adder FA_3642(s3642, c3642, in3642_1, in3642_2, pp112[25]);
    wire[0:0] s3643, in3643_1, in3643_2;
    wire c3643;
    assign in3643_1 = {pp116[21]};
    assign in3643_2 = {pp117[20]};
    Full_Adder FA_3643(s3643, c3643, in3643_1, in3643_2, pp115[22]);
    wire[0:0] s3644, in3644_1, in3644_2;
    wire c3644;
    assign in3644_1 = {pp119[18]};
    assign in3644_2 = {pp120[17]};
    Full_Adder FA_3644(s3644, c3644, in3644_1, in3644_2, pp118[19]);
    wire[0:0] s3645, in3645_1, in3645_2;
    wire c3645;
    assign in3645_1 = {pp122[15]};
    assign in3645_2 = {pp123[14]};
    Full_Adder FA_3645(s3645, c3645, in3645_1, in3645_2, pp121[16]);
    wire[0:0] s3646, in3646_1, in3646_2;
    wire c3646;
    assign in3646_1 = {pp125[12]};
    assign in3646_2 = {pp126[11]};
    Full_Adder FA_3646(s3646, c3646, in3646_1, in3646_2, pp124[13]);
    wire[0:0] s3647, in3647_1, in3647_2;
    wire c3647;
    assign in3647_1 = {c1212};
    assign in3647_2 = {c1213};
    Full_Adder FA_3647(s3647, c3647, in3647_1, in3647_2, pp127[10]);
    wire[0:0] s3648, in3648_1, in3648_2;
    wire c3648;
    assign in3648_1 = {c1215};
    assign in3648_2 = {c1216};
    Full_Adder FA_3648(s3648, c3648, in3648_1, in3648_2, c1214);
    wire[0:0] s3649, in3649_1, in3649_2;
    wire c3649;
    assign in3649_1 = {c1218};
    assign in3649_2 = {c1219};
    Full_Adder FA_3649(s3649, c3649, in3649_1, in3649_2, c1217);
    wire[0:0] s3650, in3650_1, in3650_2;
    wire c3650;
    assign in3650_1 = {c1221};
    assign in3650_2 = {c1222};
    Full_Adder FA_3650(s3650, c3650, in3650_1, in3650_2, c1220);
    wire[0:0] s3651, in3651_1, in3651_2;
    wire c3651;
    assign in3651_1 = {c1224};
    assign in3651_2 = {c1225};
    Full_Adder FA_3651(s3651, c3651, in3651_1, in3651_2, c1223);
    wire[0:0] s3652, in3652_1, in3652_2;
    wire c3652;
    assign in3652_1 = {c1227};
    assign in3652_2 = {c1228};
    Full_Adder FA_3652(s3652, c3652, in3652_1, in3652_2, c1226);
    wire[0:0] s3653, in3653_1, in3653_2;
    wire c3653;
    assign in3653_1 = {c1230};
    assign in3653_2 = {c1231};
    Full_Adder FA_3653(s3653, c3653, in3653_1, in3653_2, c1229);
    wire[0:0] s3654, in3654_1, in3654_2;
    wire c3654;
    assign in3654_1 = {c1233};
    assign in3654_2 = {c1234};
    Full_Adder FA_3654(s3654, c3654, in3654_1, in3654_2, c1232);
    wire[0:0] s3655, in3655_1, in3655_2;
    wire c3655;
    assign in3655_1 = {c1236};
    assign in3655_2 = {c1237};
    Full_Adder FA_3655(s3655, c3655, in3655_1, in3655_2, c1235);
    wire[0:0] s3656, in3656_1, in3656_2;
    wire c3656;
    assign in3656_1 = {c1239};
    assign in3656_2 = {c1240};
    Full_Adder FA_3656(s3656, c3656, in3656_1, in3656_2, c1238);
    wire[0:0] s3657, in3657_1, in3657_2;
    wire c3657;
    assign in3657_1 = {c1242};
    assign in3657_2 = {c1243};
    Full_Adder FA_3657(s3657, c3657, in3657_1, in3657_2, c1241);
    wire[0:0] s3658, in3658_1, in3658_2;
    wire c3658;
    assign in3658_1 = {c1245};
    assign in3658_2 = {s1246[0]};
    Full_Adder FA_3658(s3658, c3658, in3658_1, in3658_2, c1244);
    wire[0:0] s3659, in3659_1, in3659_2;
    wire c3659;
    assign in3659_1 = {s1248[0]};
    assign in3659_2 = {s1249[0]};
    Full_Adder FA_3659(s3659, c3659, in3659_1, in3659_2, s1247[0]);
    wire[0:0] s3660, in3660_1, in3660_2;
    wire c3660;
    assign in3660_1 = {s1251[0]};
    assign in3660_2 = {s1252[0]};
    Full_Adder FA_3660(s3660, c3660, in3660_1, in3660_2, s1250[0]);
    wire[0:0] s3661, in3661_1, in3661_2;
    wire c3661;
    assign in3661_1 = {s1254[0]};
    assign in3661_2 = {s1255[0]};
    Full_Adder FA_3661(s3661, c3661, in3661_1, in3661_2, s1253[0]);
    wire[0:0] s3662, in3662_1, in3662_2;
    wire c3662;
    assign in3662_1 = {s1257[0]};
    assign in3662_2 = {s1258[0]};
    Full_Adder FA_3662(s3662, c3662, in3662_1, in3662_2, s1256[0]);
    wire[0:0] s3663, in3663_1, in3663_2;
    wire c3663;
    assign in3663_1 = {s1260[0]};
    assign in3663_2 = {s1261[0]};
    Full_Adder FA_3663(s3663, c3663, in3663_1, in3663_2, s1259[0]);
    wire[0:0] s3664, in3664_1, in3664_2;
    wire c3664;
    assign in3664_1 = {s1263[0]};
    assign in3664_2 = {s1264[0]};
    Full_Adder FA_3664(s3664, c3664, in3664_1, in3664_2, s1262[0]);
    wire[0:0] s3665, in3665_1, in3665_2;
    wire c3665;
    assign in3665_1 = {s1266[0]};
    assign in3665_2 = {s1267[0]};
    Full_Adder FA_3665(s3665, c3665, in3665_1, in3665_2, s1265[0]);
    wire[0:0] s3666, in3666_1, in3666_2;
    wire c3666;
    assign in3666_1 = {s1269[0]};
    assign in3666_2 = {s1270[0]};
    Full_Adder FA_3666(s3666, c3666, in3666_1, in3666_2, s1268[0]);
    wire[0:0] s3667, in3667_1, in3667_2;
    wire c3667;
    assign in3667_1 = {s1272[0]};
    assign in3667_2 = {s1273[0]};
    Full_Adder FA_3667(s3667, c3667, in3667_1, in3667_2, s1271[0]);
    wire[0:0] s3668, in3668_1, in3668_2;
    wire c3668;
    assign in3668_1 = {s1275[0]};
    assign in3668_2 = {s1276[0]};
    Full_Adder FA_3668(s3668, c3668, in3668_1, in3668_2, s1274[0]);
    wire[0:0] s3669, in3669_1, in3669_2;
    wire c3669;
    assign in3669_1 = {pp108[30]};
    assign in3669_2 = {pp109[29]};
    Full_Adder FA_3669(s3669, c3669, in3669_1, in3669_2, pp107[31]);
    wire[0:0] s3670, in3670_1, in3670_2;
    wire c3670;
    assign in3670_1 = {pp111[27]};
    assign in3670_2 = {pp112[26]};
    Full_Adder FA_3670(s3670, c3670, in3670_1, in3670_2, pp110[28]);
    wire[0:0] s3671, in3671_1, in3671_2;
    wire c3671;
    assign in3671_1 = {pp114[24]};
    assign in3671_2 = {pp115[23]};
    Full_Adder FA_3671(s3671, c3671, in3671_1, in3671_2, pp113[25]);
    wire[0:0] s3672, in3672_1, in3672_2;
    wire c3672;
    assign in3672_1 = {pp117[21]};
    assign in3672_2 = {pp118[20]};
    Full_Adder FA_3672(s3672, c3672, in3672_1, in3672_2, pp116[22]);
    wire[0:0] s3673, in3673_1, in3673_2;
    wire c3673;
    assign in3673_1 = {pp120[18]};
    assign in3673_2 = {pp121[17]};
    Full_Adder FA_3673(s3673, c3673, in3673_1, in3673_2, pp119[19]);
    wire[0:0] s3674, in3674_1, in3674_2;
    wire c3674;
    assign in3674_1 = {pp123[15]};
    assign in3674_2 = {pp124[14]};
    Full_Adder FA_3674(s3674, c3674, in3674_1, in3674_2, pp122[16]);
    wire[0:0] s3675, in3675_1, in3675_2;
    wire c3675;
    assign in3675_1 = {pp126[12]};
    assign in3675_2 = {pp127[11]};
    Full_Adder FA_3675(s3675, c3675, in3675_1, in3675_2, pp125[13]);
    wire[0:0] s3676, in3676_1, in3676_2;
    wire c3676;
    assign in3676_1 = {c1247};
    assign in3676_2 = {c1248};
    Full_Adder FA_3676(s3676, c3676, in3676_1, in3676_2, c1246);
    wire[0:0] s3677, in3677_1, in3677_2;
    wire c3677;
    assign in3677_1 = {c1250};
    assign in3677_2 = {c1251};
    Full_Adder FA_3677(s3677, c3677, in3677_1, in3677_2, c1249);
    wire[0:0] s3678, in3678_1, in3678_2;
    wire c3678;
    assign in3678_1 = {c1253};
    assign in3678_2 = {c1254};
    Full_Adder FA_3678(s3678, c3678, in3678_1, in3678_2, c1252);
    wire[0:0] s3679, in3679_1, in3679_2;
    wire c3679;
    assign in3679_1 = {c1256};
    assign in3679_2 = {c1257};
    Full_Adder FA_3679(s3679, c3679, in3679_1, in3679_2, c1255);
    wire[0:0] s3680, in3680_1, in3680_2;
    wire c3680;
    assign in3680_1 = {c1259};
    assign in3680_2 = {c1260};
    Full_Adder FA_3680(s3680, c3680, in3680_1, in3680_2, c1258);
    wire[0:0] s3681, in3681_1, in3681_2;
    wire c3681;
    assign in3681_1 = {c1262};
    assign in3681_2 = {c1263};
    Full_Adder FA_3681(s3681, c3681, in3681_1, in3681_2, c1261);
    wire[0:0] s3682, in3682_1, in3682_2;
    wire c3682;
    assign in3682_1 = {c1265};
    assign in3682_2 = {c1266};
    Full_Adder FA_3682(s3682, c3682, in3682_1, in3682_2, c1264);
    wire[0:0] s3683, in3683_1, in3683_2;
    wire c3683;
    assign in3683_1 = {c1268};
    assign in3683_2 = {c1269};
    Full_Adder FA_3683(s3683, c3683, in3683_1, in3683_2, c1267);
    wire[0:0] s3684, in3684_1, in3684_2;
    wire c3684;
    assign in3684_1 = {c1271};
    assign in3684_2 = {c1272};
    Full_Adder FA_3684(s3684, c3684, in3684_1, in3684_2, c1270);
    wire[0:0] s3685, in3685_1, in3685_2;
    wire c3685;
    assign in3685_1 = {c1274};
    assign in3685_2 = {c1275};
    Full_Adder FA_3685(s3685, c3685, in3685_1, in3685_2, c1273);
    wire[0:0] s3686, in3686_1, in3686_2;
    wire c3686;
    assign in3686_1 = {c1277};
    assign in3686_2 = {c1278};
    Full_Adder FA_3686(s3686, c3686, in3686_1, in3686_2, c1276);
    wire[0:0] s3687, in3687_1, in3687_2;
    wire c3687;
    assign in3687_1 = {s1280[0]};
    assign in3687_2 = {s1281[0]};
    Full_Adder FA_3687(s3687, c3687, in3687_1, in3687_2, s1279[0]);
    wire[0:0] s3688, in3688_1, in3688_2;
    wire c3688;
    assign in3688_1 = {s1283[0]};
    assign in3688_2 = {s1284[0]};
    Full_Adder FA_3688(s3688, c3688, in3688_1, in3688_2, s1282[0]);
    wire[0:0] s3689, in3689_1, in3689_2;
    wire c3689;
    assign in3689_1 = {s1286[0]};
    assign in3689_2 = {s1287[0]};
    Full_Adder FA_3689(s3689, c3689, in3689_1, in3689_2, s1285[0]);
    wire[0:0] s3690, in3690_1, in3690_2;
    wire c3690;
    assign in3690_1 = {s1289[0]};
    assign in3690_2 = {s1290[0]};
    Full_Adder FA_3690(s3690, c3690, in3690_1, in3690_2, s1288[0]);
    wire[0:0] s3691, in3691_1, in3691_2;
    wire c3691;
    assign in3691_1 = {s1292[0]};
    assign in3691_2 = {s1293[0]};
    Full_Adder FA_3691(s3691, c3691, in3691_1, in3691_2, s1291[0]);
    wire[0:0] s3692, in3692_1, in3692_2;
    wire c3692;
    assign in3692_1 = {s1295[0]};
    assign in3692_2 = {s1296[0]};
    Full_Adder FA_3692(s3692, c3692, in3692_1, in3692_2, s1294[0]);
    wire[0:0] s3693, in3693_1, in3693_2;
    wire c3693;
    assign in3693_1 = {s1298[0]};
    assign in3693_2 = {s1299[0]};
    Full_Adder FA_3693(s3693, c3693, in3693_1, in3693_2, s1297[0]);
    wire[0:0] s3694, in3694_1, in3694_2;
    wire c3694;
    assign in3694_1 = {s1301[0]};
    assign in3694_2 = {s1302[0]};
    Full_Adder FA_3694(s3694, c3694, in3694_1, in3694_2, s1300[0]);
    wire[0:0] s3695, in3695_1, in3695_2;
    wire c3695;
    assign in3695_1 = {s1304[0]};
    assign in3695_2 = {s1305[0]};
    Full_Adder FA_3695(s3695, c3695, in3695_1, in3695_2, s1303[0]);
    wire[0:0] s3696, in3696_1, in3696_2;
    wire c3696;
    assign in3696_1 = {s1307[0]};
    assign in3696_2 = {s1308[0]};
    Full_Adder FA_3696(s3696, c3696, in3696_1, in3696_2, s1306[0]);
    wire[0:0] s3697, in3697_1, in3697_2;
    wire c3697;
    assign in3697_1 = {pp106[33]};
    assign in3697_2 = {pp107[32]};
    Full_Adder FA_3697(s3697, c3697, in3697_1, in3697_2, pp105[34]);
    wire[0:0] s3698, in3698_1, in3698_2;
    wire c3698;
    assign in3698_1 = {pp109[30]};
    assign in3698_2 = {pp110[29]};
    Full_Adder FA_3698(s3698, c3698, in3698_1, in3698_2, pp108[31]);
    wire[0:0] s3699, in3699_1, in3699_2;
    wire c3699;
    assign in3699_1 = {pp112[27]};
    assign in3699_2 = {pp113[26]};
    Full_Adder FA_3699(s3699, c3699, in3699_1, in3699_2, pp111[28]);
    wire[0:0] s3700, in3700_1, in3700_2;
    wire c3700;
    assign in3700_1 = {pp115[24]};
    assign in3700_2 = {pp116[23]};
    Full_Adder FA_3700(s3700, c3700, in3700_1, in3700_2, pp114[25]);
    wire[0:0] s3701, in3701_1, in3701_2;
    wire c3701;
    assign in3701_1 = {pp118[21]};
    assign in3701_2 = {pp119[20]};
    Full_Adder FA_3701(s3701, c3701, in3701_1, in3701_2, pp117[22]);
    wire[0:0] s3702, in3702_1, in3702_2;
    wire c3702;
    assign in3702_1 = {pp121[18]};
    assign in3702_2 = {pp122[17]};
    Full_Adder FA_3702(s3702, c3702, in3702_1, in3702_2, pp120[19]);
    wire[0:0] s3703, in3703_1, in3703_2;
    wire c3703;
    assign in3703_1 = {pp124[15]};
    assign in3703_2 = {pp125[14]};
    Full_Adder FA_3703(s3703, c3703, in3703_1, in3703_2, pp123[16]);
    wire[0:0] s3704, in3704_1, in3704_2;
    wire c3704;
    assign in3704_1 = {pp127[12]};
    assign in3704_2 = {c1279};
    Full_Adder FA_3704(s3704, c3704, in3704_1, in3704_2, pp126[13]);
    wire[0:0] s3705, in3705_1, in3705_2;
    wire c3705;
    assign in3705_1 = {c1281};
    assign in3705_2 = {c1282};
    Full_Adder FA_3705(s3705, c3705, in3705_1, in3705_2, c1280);
    wire[0:0] s3706, in3706_1, in3706_2;
    wire c3706;
    assign in3706_1 = {c1284};
    assign in3706_2 = {c1285};
    Full_Adder FA_3706(s3706, c3706, in3706_1, in3706_2, c1283);
    wire[0:0] s3707, in3707_1, in3707_2;
    wire c3707;
    assign in3707_1 = {c1287};
    assign in3707_2 = {c1288};
    Full_Adder FA_3707(s3707, c3707, in3707_1, in3707_2, c1286);
    wire[0:0] s3708, in3708_1, in3708_2;
    wire c3708;
    assign in3708_1 = {c1290};
    assign in3708_2 = {c1291};
    Full_Adder FA_3708(s3708, c3708, in3708_1, in3708_2, c1289);
    wire[0:0] s3709, in3709_1, in3709_2;
    wire c3709;
    assign in3709_1 = {c1293};
    assign in3709_2 = {c1294};
    Full_Adder FA_3709(s3709, c3709, in3709_1, in3709_2, c1292);
    wire[0:0] s3710, in3710_1, in3710_2;
    wire c3710;
    assign in3710_1 = {c1296};
    assign in3710_2 = {c1297};
    Full_Adder FA_3710(s3710, c3710, in3710_1, in3710_2, c1295);
    wire[0:0] s3711, in3711_1, in3711_2;
    wire c3711;
    assign in3711_1 = {c1299};
    assign in3711_2 = {c1300};
    Full_Adder FA_3711(s3711, c3711, in3711_1, in3711_2, c1298);
    wire[0:0] s3712, in3712_1, in3712_2;
    wire c3712;
    assign in3712_1 = {c1302};
    assign in3712_2 = {c1303};
    Full_Adder FA_3712(s3712, c3712, in3712_1, in3712_2, c1301);
    wire[0:0] s3713, in3713_1, in3713_2;
    wire c3713;
    assign in3713_1 = {c1305};
    assign in3713_2 = {c1306};
    Full_Adder FA_3713(s3713, c3713, in3713_1, in3713_2, c1304);
    wire[0:0] s3714, in3714_1, in3714_2;
    wire c3714;
    assign in3714_1 = {c1308};
    assign in3714_2 = {c1309};
    Full_Adder FA_3714(s3714, c3714, in3714_1, in3714_2, c1307);
    wire[0:0] s3715, in3715_1, in3715_2;
    wire c3715;
    assign in3715_1 = {s1311[0]};
    assign in3715_2 = {s1312[0]};
    Full_Adder FA_3715(s3715, c3715, in3715_1, in3715_2, c1310);
    wire[0:0] s3716, in3716_1, in3716_2;
    wire c3716;
    assign in3716_1 = {s1314[0]};
    assign in3716_2 = {s1315[0]};
    Full_Adder FA_3716(s3716, c3716, in3716_1, in3716_2, s1313[0]);
    wire[0:0] s3717, in3717_1, in3717_2;
    wire c3717;
    assign in3717_1 = {s1317[0]};
    assign in3717_2 = {s1318[0]};
    Full_Adder FA_3717(s3717, c3717, in3717_1, in3717_2, s1316[0]);
    wire[0:0] s3718, in3718_1, in3718_2;
    wire c3718;
    assign in3718_1 = {s1320[0]};
    assign in3718_2 = {s1321[0]};
    Full_Adder FA_3718(s3718, c3718, in3718_1, in3718_2, s1319[0]);
    wire[0:0] s3719, in3719_1, in3719_2;
    wire c3719;
    assign in3719_1 = {s1323[0]};
    assign in3719_2 = {s1324[0]};
    Full_Adder FA_3719(s3719, c3719, in3719_1, in3719_2, s1322[0]);
    wire[0:0] s3720, in3720_1, in3720_2;
    wire c3720;
    assign in3720_1 = {s1326[0]};
    assign in3720_2 = {s1327[0]};
    Full_Adder FA_3720(s3720, c3720, in3720_1, in3720_2, s1325[0]);
    wire[0:0] s3721, in3721_1, in3721_2;
    wire c3721;
    assign in3721_1 = {s1329[0]};
    assign in3721_2 = {s1330[0]};
    Full_Adder FA_3721(s3721, c3721, in3721_1, in3721_2, s1328[0]);
    wire[0:0] s3722, in3722_1, in3722_2;
    wire c3722;
    assign in3722_1 = {s1332[0]};
    assign in3722_2 = {s1333[0]};
    Full_Adder FA_3722(s3722, c3722, in3722_1, in3722_2, s1331[0]);
    wire[0:0] s3723, in3723_1, in3723_2;
    wire c3723;
    assign in3723_1 = {s1335[0]};
    assign in3723_2 = {s1336[0]};
    Full_Adder FA_3723(s3723, c3723, in3723_1, in3723_2, s1334[0]);
    wire[0:0] s3724, in3724_1, in3724_2;
    wire c3724;
    assign in3724_1 = {s1338[0]};
    assign in3724_2 = {s1339[0]};
    Full_Adder FA_3724(s3724, c3724, in3724_1, in3724_2, s1337[0]);
    wire[0:0] s3725, in3725_1, in3725_2;
    wire c3725;
    assign in3725_1 = {pp104[36]};
    assign in3725_2 = {pp105[35]};
    Full_Adder FA_3725(s3725, c3725, in3725_1, in3725_2, pp103[37]);
    wire[0:0] s3726, in3726_1, in3726_2;
    wire c3726;
    assign in3726_1 = {pp107[33]};
    assign in3726_2 = {pp108[32]};
    Full_Adder FA_3726(s3726, c3726, in3726_1, in3726_2, pp106[34]);
    wire[0:0] s3727, in3727_1, in3727_2;
    wire c3727;
    assign in3727_1 = {pp110[30]};
    assign in3727_2 = {pp111[29]};
    Full_Adder FA_3727(s3727, c3727, in3727_1, in3727_2, pp109[31]);
    wire[0:0] s3728, in3728_1, in3728_2;
    wire c3728;
    assign in3728_1 = {pp113[27]};
    assign in3728_2 = {pp114[26]};
    Full_Adder FA_3728(s3728, c3728, in3728_1, in3728_2, pp112[28]);
    wire[0:0] s3729, in3729_1, in3729_2;
    wire c3729;
    assign in3729_1 = {pp116[24]};
    assign in3729_2 = {pp117[23]};
    Full_Adder FA_3729(s3729, c3729, in3729_1, in3729_2, pp115[25]);
    wire[0:0] s3730, in3730_1, in3730_2;
    wire c3730;
    assign in3730_1 = {pp119[21]};
    assign in3730_2 = {pp120[20]};
    Full_Adder FA_3730(s3730, c3730, in3730_1, in3730_2, pp118[22]);
    wire[0:0] s3731, in3731_1, in3731_2;
    wire c3731;
    assign in3731_1 = {pp122[18]};
    assign in3731_2 = {pp123[17]};
    Full_Adder FA_3731(s3731, c3731, in3731_1, in3731_2, pp121[19]);
    wire[0:0] s3732, in3732_1, in3732_2;
    wire c3732;
    assign in3732_1 = {pp125[15]};
    assign in3732_2 = {pp126[14]};
    Full_Adder FA_3732(s3732, c3732, in3732_1, in3732_2, pp124[16]);
    wire[0:0] s3733, in3733_1, in3733_2;
    wire c3733;
    assign in3733_1 = {c1311};
    assign in3733_2 = {c1312};
    Full_Adder FA_3733(s3733, c3733, in3733_1, in3733_2, pp127[13]);
    wire[0:0] s3734, in3734_1, in3734_2;
    wire c3734;
    assign in3734_1 = {c1314};
    assign in3734_2 = {c1315};
    Full_Adder FA_3734(s3734, c3734, in3734_1, in3734_2, c1313);
    wire[0:0] s3735, in3735_1, in3735_2;
    wire c3735;
    assign in3735_1 = {c1317};
    assign in3735_2 = {c1318};
    Full_Adder FA_3735(s3735, c3735, in3735_1, in3735_2, c1316);
    wire[0:0] s3736, in3736_1, in3736_2;
    wire c3736;
    assign in3736_1 = {c1320};
    assign in3736_2 = {c1321};
    Full_Adder FA_3736(s3736, c3736, in3736_1, in3736_2, c1319);
    wire[0:0] s3737, in3737_1, in3737_2;
    wire c3737;
    assign in3737_1 = {c1323};
    assign in3737_2 = {c1324};
    Full_Adder FA_3737(s3737, c3737, in3737_1, in3737_2, c1322);
    wire[0:0] s3738, in3738_1, in3738_2;
    wire c3738;
    assign in3738_1 = {c1326};
    assign in3738_2 = {c1327};
    Full_Adder FA_3738(s3738, c3738, in3738_1, in3738_2, c1325);
    wire[0:0] s3739, in3739_1, in3739_2;
    wire c3739;
    assign in3739_1 = {c1329};
    assign in3739_2 = {c1330};
    Full_Adder FA_3739(s3739, c3739, in3739_1, in3739_2, c1328);
    wire[0:0] s3740, in3740_1, in3740_2;
    wire c3740;
    assign in3740_1 = {c1332};
    assign in3740_2 = {c1333};
    Full_Adder FA_3740(s3740, c3740, in3740_1, in3740_2, c1331);
    wire[0:0] s3741, in3741_1, in3741_2;
    wire c3741;
    assign in3741_1 = {c1335};
    assign in3741_2 = {c1336};
    Full_Adder FA_3741(s3741, c3741, in3741_1, in3741_2, c1334);
    wire[0:0] s3742, in3742_1, in3742_2;
    wire c3742;
    assign in3742_1 = {c1338};
    assign in3742_2 = {c1339};
    Full_Adder FA_3742(s3742, c3742, in3742_1, in3742_2, c1337);
    wire[0:0] s3743, in3743_1, in3743_2;
    wire c3743;
    assign in3743_1 = {c1341};
    assign in3743_2 = {s1342[0]};
    Full_Adder FA_3743(s3743, c3743, in3743_1, in3743_2, c1340);
    wire[0:0] s3744, in3744_1, in3744_2;
    wire c3744;
    assign in3744_1 = {s1344[0]};
    assign in3744_2 = {s1345[0]};
    Full_Adder FA_3744(s3744, c3744, in3744_1, in3744_2, s1343[0]);
    wire[0:0] s3745, in3745_1, in3745_2;
    wire c3745;
    assign in3745_1 = {s1347[0]};
    assign in3745_2 = {s1348[0]};
    Full_Adder FA_3745(s3745, c3745, in3745_1, in3745_2, s1346[0]);
    wire[0:0] s3746, in3746_1, in3746_2;
    wire c3746;
    assign in3746_1 = {s1350[0]};
    assign in3746_2 = {s1351[0]};
    Full_Adder FA_3746(s3746, c3746, in3746_1, in3746_2, s1349[0]);
    wire[0:0] s3747, in3747_1, in3747_2;
    wire c3747;
    assign in3747_1 = {s1353[0]};
    assign in3747_2 = {s1354[0]};
    Full_Adder FA_3747(s3747, c3747, in3747_1, in3747_2, s1352[0]);
    wire[0:0] s3748, in3748_1, in3748_2;
    wire c3748;
    assign in3748_1 = {s1356[0]};
    assign in3748_2 = {s1357[0]};
    Full_Adder FA_3748(s3748, c3748, in3748_1, in3748_2, s1355[0]);
    wire[0:0] s3749, in3749_1, in3749_2;
    wire c3749;
    assign in3749_1 = {s1359[0]};
    assign in3749_2 = {s1360[0]};
    Full_Adder FA_3749(s3749, c3749, in3749_1, in3749_2, s1358[0]);
    wire[0:0] s3750, in3750_1, in3750_2;
    wire c3750;
    assign in3750_1 = {s1362[0]};
    assign in3750_2 = {s1363[0]};
    Full_Adder FA_3750(s3750, c3750, in3750_1, in3750_2, s1361[0]);
    wire[0:0] s3751, in3751_1, in3751_2;
    wire c3751;
    assign in3751_1 = {s1365[0]};
    assign in3751_2 = {s1366[0]};
    Full_Adder FA_3751(s3751, c3751, in3751_1, in3751_2, s1364[0]);
    wire[0:0] s3752, in3752_1, in3752_2;
    wire c3752;
    assign in3752_1 = {s1368[0]};
    assign in3752_2 = {s1369[0]};
    Full_Adder FA_3752(s3752, c3752, in3752_1, in3752_2, s1367[0]);
    wire[0:0] s3753, in3753_1, in3753_2;
    wire c3753;
    assign in3753_1 = {pp102[39]};
    assign in3753_2 = {pp103[38]};
    Full_Adder FA_3753(s3753, c3753, in3753_1, in3753_2, pp101[40]);
    wire[0:0] s3754, in3754_1, in3754_2;
    wire c3754;
    assign in3754_1 = {pp105[36]};
    assign in3754_2 = {pp106[35]};
    Full_Adder FA_3754(s3754, c3754, in3754_1, in3754_2, pp104[37]);
    wire[0:0] s3755, in3755_1, in3755_2;
    wire c3755;
    assign in3755_1 = {pp108[33]};
    assign in3755_2 = {pp109[32]};
    Full_Adder FA_3755(s3755, c3755, in3755_1, in3755_2, pp107[34]);
    wire[0:0] s3756, in3756_1, in3756_2;
    wire c3756;
    assign in3756_1 = {pp111[30]};
    assign in3756_2 = {pp112[29]};
    Full_Adder FA_3756(s3756, c3756, in3756_1, in3756_2, pp110[31]);
    wire[0:0] s3757, in3757_1, in3757_2;
    wire c3757;
    assign in3757_1 = {pp114[27]};
    assign in3757_2 = {pp115[26]};
    Full_Adder FA_3757(s3757, c3757, in3757_1, in3757_2, pp113[28]);
    wire[0:0] s3758, in3758_1, in3758_2;
    wire c3758;
    assign in3758_1 = {pp117[24]};
    assign in3758_2 = {pp118[23]};
    Full_Adder FA_3758(s3758, c3758, in3758_1, in3758_2, pp116[25]);
    wire[0:0] s3759, in3759_1, in3759_2;
    wire c3759;
    assign in3759_1 = {pp120[21]};
    assign in3759_2 = {pp121[20]};
    Full_Adder FA_3759(s3759, c3759, in3759_1, in3759_2, pp119[22]);
    wire[0:0] s3760, in3760_1, in3760_2;
    wire c3760;
    assign in3760_1 = {pp123[18]};
    assign in3760_2 = {pp124[17]};
    Full_Adder FA_3760(s3760, c3760, in3760_1, in3760_2, pp122[19]);
    wire[0:0] s3761, in3761_1, in3761_2;
    wire c3761;
    assign in3761_1 = {pp126[15]};
    assign in3761_2 = {pp127[14]};
    Full_Adder FA_3761(s3761, c3761, in3761_1, in3761_2, pp125[16]);
    wire[0:0] s3762, in3762_1, in3762_2;
    wire c3762;
    assign in3762_1 = {c1343};
    assign in3762_2 = {c1344};
    Full_Adder FA_3762(s3762, c3762, in3762_1, in3762_2, c1342);
    wire[0:0] s3763, in3763_1, in3763_2;
    wire c3763;
    assign in3763_1 = {c1346};
    assign in3763_2 = {c1347};
    Full_Adder FA_3763(s3763, c3763, in3763_1, in3763_2, c1345);
    wire[0:0] s3764, in3764_1, in3764_2;
    wire c3764;
    assign in3764_1 = {c1349};
    assign in3764_2 = {c1350};
    Full_Adder FA_3764(s3764, c3764, in3764_1, in3764_2, c1348);
    wire[0:0] s3765, in3765_1, in3765_2;
    wire c3765;
    assign in3765_1 = {c1352};
    assign in3765_2 = {c1353};
    Full_Adder FA_3765(s3765, c3765, in3765_1, in3765_2, c1351);
    wire[0:0] s3766, in3766_1, in3766_2;
    wire c3766;
    assign in3766_1 = {c1355};
    assign in3766_2 = {c1356};
    Full_Adder FA_3766(s3766, c3766, in3766_1, in3766_2, c1354);
    wire[0:0] s3767, in3767_1, in3767_2;
    wire c3767;
    assign in3767_1 = {c1358};
    assign in3767_2 = {c1359};
    Full_Adder FA_3767(s3767, c3767, in3767_1, in3767_2, c1357);
    wire[0:0] s3768, in3768_1, in3768_2;
    wire c3768;
    assign in3768_1 = {c1361};
    assign in3768_2 = {c1362};
    Full_Adder FA_3768(s3768, c3768, in3768_1, in3768_2, c1360);
    wire[0:0] s3769, in3769_1, in3769_2;
    wire c3769;
    assign in3769_1 = {c1364};
    assign in3769_2 = {c1365};
    Full_Adder FA_3769(s3769, c3769, in3769_1, in3769_2, c1363);
    wire[0:0] s3770, in3770_1, in3770_2;
    wire c3770;
    assign in3770_1 = {c1367};
    assign in3770_2 = {c1368};
    Full_Adder FA_3770(s3770, c3770, in3770_1, in3770_2, c1366);
    wire[0:0] s3771, in3771_1, in3771_2;
    wire c3771;
    assign in3771_1 = {c1370};
    assign in3771_2 = {c1371};
    Full_Adder FA_3771(s3771, c3771, in3771_1, in3771_2, c1369);
    wire[0:0] s3772, in3772_1, in3772_2;
    wire c3772;
    assign in3772_1 = {s1373[0]};
    assign in3772_2 = {s1374[0]};
    Full_Adder FA_3772(s3772, c3772, in3772_1, in3772_2, s1372[0]);
    wire[0:0] s3773, in3773_1, in3773_2;
    wire c3773;
    assign in3773_1 = {s1376[0]};
    assign in3773_2 = {s1377[0]};
    Full_Adder FA_3773(s3773, c3773, in3773_1, in3773_2, s1375[0]);
    wire[0:0] s3774, in3774_1, in3774_2;
    wire c3774;
    assign in3774_1 = {s1379[0]};
    assign in3774_2 = {s1380[0]};
    Full_Adder FA_3774(s3774, c3774, in3774_1, in3774_2, s1378[0]);
    wire[0:0] s3775, in3775_1, in3775_2;
    wire c3775;
    assign in3775_1 = {s1382[0]};
    assign in3775_2 = {s1383[0]};
    Full_Adder FA_3775(s3775, c3775, in3775_1, in3775_2, s1381[0]);
    wire[0:0] s3776, in3776_1, in3776_2;
    wire c3776;
    assign in3776_1 = {s1385[0]};
    assign in3776_2 = {s1386[0]};
    Full_Adder FA_3776(s3776, c3776, in3776_1, in3776_2, s1384[0]);
    wire[0:0] s3777, in3777_1, in3777_2;
    wire c3777;
    assign in3777_1 = {s1388[0]};
    assign in3777_2 = {s1389[0]};
    Full_Adder FA_3777(s3777, c3777, in3777_1, in3777_2, s1387[0]);
    wire[0:0] s3778, in3778_1, in3778_2;
    wire c3778;
    assign in3778_1 = {s1391[0]};
    assign in3778_2 = {s1392[0]};
    Full_Adder FA_3778(s3778, c3778, in3778_1, in3778_2, s1390[0]);
    wire[0:0] s3779, in3779_1, in3779_2;
    wire c3779;
    assign in3779_1 = {s1394[0]};
    assign in3779_2 = {s1395[0]};
    Full_Adder FA_3779(s3779, c3779, in3779_1, in3779_2, s1393[0]);
    wire[0:0] s3780, in3780_1, in3780_2;
    wire c3780;
    assign in3780_1 = {s1397[0]};
    assign in3780_2 = {s1398[0]};
    Full_Adder FA_3780(s3780, c3780, in3780_1, in3780_2, s1396[0]);
    wire[0:0] s3781, in3781_1, in3781_2;
    wire c3781;
    assign in3781_1 = {pp100[42]};
    assign in3781_2 = {pp101[41]};
    Full_Adder FA_3781(s3781, c3781, in3781_1, in3781_2, pp99[43]);
    wire[0:0] s3782, in3782_1, in3782_2;
    wire c3782;
    assign in3782_1 = {pp103[39]};
    assign in3782_2 = {pp104[38]};
    Full_Adder FA_3782(s3782, c3782, in3782_1, in3782_2, pp102[40]);
    wire[0:0] s3783, in3783_1, in3783_2;
    wire c3783;
    assign in3783_1 = {pp106[36]};
    assign in3783_2 = {pp107[35]};
    Full_Adder FA_3783(s3783, c3783, in3783_1, in3783_2, pp105[37]);
    wire[0:0] s3784, in3784_1, in3784_2;
    wire c3784;
    assign in3784_1 = {pp109[33]};
    assign in3784_2 = {pp110[32]};
    Full_Adder FA_3784(s3784, c3784, in3784_1, in3784_2, pp108[34]);
    wire[0:0] s3785, in3785_1, in3785_2;
    wire c3785;
    assign in3785_1 = {pp112[30]};
    assign in3785_2 = {pp113[29]};
    Full_Adder FA_3785(s3785, c3785, in3785_1, in3785_2, pp111[31]);
    wire[0:0] s3786, in3786_1, in3786_2;
    wire c3786;
    assign in3786_1 = {pp115[27]};
    assign in3786_2 = {pp116[26]};
    Full_Adder FA_3786(s3786, c3786, in3786_1, in3786_2, pp114[28]);
    wire[0:0] s3787, in3787_1, in3787_2;
    wire c3787;
    assign in3787_1 = {pp118[24]};
    assign in3787_2 = {pp119[23]};
    Full_Adder FA_3787(s3787, c3787, in3787_1, in3787_2, pp117[25]);
    wire[0:0] s3788, in3788_1, in3788_2;
    wire c3788;
    assign in3788_1 = {pp121[21]};
    assign in3788_2 = {pp122[20]};
    Full_Adder FA_3788(s3788, c3788, in3788_1, in3788_2, pp120[22]);
    wire[0:0] s3789, in3789_1, in3789_2;
    wire c3789;
    assign in3789_1 = {pp124[18]};
    assign in3789_2 = {pp125[17]};
    Full_Adder FA_3789(s3789, c3789, in3789_1, in3789_2, pp123[19]);
    wire[0:0] s3790, in3790_1, in3790_2;
    wire c3790;
    assign in3790_1 = {pp127[15]};
    assign in3790_2 = {c1372};
    Full_Adder FA_3790(s3790, c3790, in3790_1, in3790_2, pp126[16]);
    wire[0:0] s3791, in3791_1, in3791_2;
    wire c3791;
    assign in3791_1 = {c1374};
    assign in3791_2 = {c1375};
    Full_Adder FA_3791(s3791, c3791, in3791_1, in3791_2, c1373);
    wire[0:0] s3792, in3792_1, in3792_2;
    wire c3792;
    assign in3792_1 = {c1377};
    assign in3792_2 = {c1378};
    Full_Adder FA_3792(s3792, c3792, in3792_1, in3792_2, c1376);
    wire[0:0] s3793, in3793_1, in3793_2;
    wire c3793;
    assign in3793_1 = {c1380};
    assign in3793_2 = {c1381};
    Full_Adder FA_3793(s3793, c3793, in3793_1, in3793_2, c1379);
    wire[0:0] s3794, in3794_1, in3794_2;
    wire c3794;
    assign in3794_1 = {c1383};
    assign in3794_2 = {c1384};
    Full_Adder FA_3794(s3794, c3794, in3794_1, in3794_2, c1382);
    wire[0:0] s3795, in3795_1, in3795_2;
    wire c3795;
    assign in3795_1 = {c1386};
    assign in3795_2 = {c1387};
    Full_Adder FA_3795(s3795, c3795, in3795_1, in3795_2, c1385);
    wire[0:0] s3796, in3796_1, in3796_2;
    wire c3796;
    assign in3796_1 = {c1389};
    assign in3796_2 = {c1390};
    Full_Adder FA_3796(s3796, c3796, in3796_1, in3796_2, c1388);
    wire[0:0] s3797, in3797_1, in3797_2;
    wire c3797;
    assign in3797_1 = {c1392};
    assign in3797_2 = {c1393};
    Full_Adder FA_3797(s3797, c3797, in3797_1, in3797_2, c1391);
    wire[0:0] s3798, in3798_1, in3798_2;
    wire c3798;
    assign in3798_1 = {c1395};
    assign in3798_2 = {c1396};
    Full_Adder FA_3798(s3798, c3798, in3798_1, in3798_2, c1394);
    wire[0:0] s3799, in3799_1, in3799_2;
    wire c3799;
    assign in3799_1 = {c1398};
    assign in3799_2 = {c1399};
    Full_Adder FA_3799(s3799, c3799, in3799_1, in3799_2, c1397);
    wire[0:0] s3800, in3800_1, in3800_2;
    wire c3800;
    assign in3800_1 = {s1401[0]};
    assign in3800_2 = {s1402[0]};
    Full_Adder FA_3800(s3800, c3800, in3800_1, in3800_2, c1400);
    wire[0:0] s3801, in3801_1, in3801_2;
    wire c3801;
    assign in3801_1 = {s1404[0]};
    assign in3801_2 = {s1405[0]};
    Full_Adder FA_3801(s3801, c3801, in3801_1, in3801_2, s1403[0]);
    wire[0:0] s3802, in3802_1, in3802_2;
    wire c3802;
    assign in3802_1 = {s1407[0]};
    assign in3802_2 = {s1408[0]};
    Full_Adder FA_3802(s3802, c3802, in3802_1, in3802_2, s1406[0]);
    wire[0:0] s3803, in3803_1, in3803_2;
    wire c3803;
    assign in3803_1 = {s1410[0]};
    assign in3803_2 = {s1411[0]};
    Full_Adder FA_3803(s3803, c3803, in3803_1, in3803_2, s1409[0]);
    wire[0:0] s3804, in3804_1, in3804_2;
    wire c3804;
    assign in3804_1 = {s1413[0]};
    assign in3804_2 = {s1414[0]};
    Full_Adder FA_3804(s3804, c3804, in3804_1, in3804_2, s1412[0]);
    wire[0:0] s3805, in3805_1, in3805_2;
    wire c3805;
    assign in3805_1 = {s1416[0]};
    assign in3805_2 = {s1417[0]};
    Full_Adder FA_3805(s3805, c3805, in3805_1, in3805_2, s1415[0]);
    wire[0:0] s3806, in3806_1, in3806_2;
    wire c3806;
    assign in3806_1 = {s1419[0]};
    assign in3806_2 = {s1420[0]};
    Full_Adder FA_3806(s3806, c3806, in3806_1, in3806_2, s1418[0]);
    wire[0:0] s3807, in3807_1, in3807_2;
    wire c3807;
    assign in3807_1 = {s1422[0]};
    assign in3807_2 = {s1423[0]};
    Full_Adder FA_3807(s3807, c3807, in3807_1, in3807_2, s1421[0]);
    wire[0:0] s3808, in3808_1, in3808_2;
    wire c3808;
    assign in3808_1 = {s1425[0]};
    assign in3808_2 = {s1426[0]};
    Full_Adder FA_3808(s3808, c3808, in3808_1, in3808_2, s1424[0]);
    wire[0:0] s3809, in3809_1, in3809_2;
    wire c3809;
    assign in3809_1 = {pp98[45]};
    assign in3809_2 = {pp99[44]};
    Full_Adder FA_3809(s3809, c3809, in3809_1, in3809_2, pp97[46]);
    wire[0:0] s3810, in3810_1, in3810_2;
    wire c3810;
    assign in3810_1 = {pp101[42]};
    assign in3810_2 = {pp102[41]};
    Full_Adder FA_3810(s3810, c3810, in3810_1, in3810_2, pp100[43]);
    wire[0:0] s3811, in3811_1, in3811_2;
    wire c3811;
    assign in3811_1 = {pp104[39]};
    assign in3811_2 = {pp105[38]};
    Full_Adder FA_3811(s3811, c3811, in3811_1, in3811_2, pp103[40]);
    wire[0:0] s3812, in3812_1, in3812_2;
    wire c3812;
    assign in3812_1 = {pp107[36]};
    assign in3812_2 = {pp108[35]};
    Full_Adder FA_3812(s3812, c3812, in3812_1, in3812_2, pp106[37]);
    wire[0:0] s3813, in3813_1, in3813_2;
    wire c3813;
    assign in3813_1 = {pp110[33]};
    assign in3813_2 = {pp111[32]};
    Full_Adder FA_3813(s3813, c3813, in3813_1, in3813_2, pp109[34]);
    wire[0:0] s3814, in3814_1, in3814_2;
    wire c3814;
    assign in3814_1 = {pp113[30]};
    assign in3814_2 = {pp114[29]};
    Full_Adder FA_3814(s3814, c3814, in3814_1, in3814_2, pp112[31]);
    wire[0:0] s3815, in3815_1, in3815_2;
    wire c3815;
    assign in3815_1 = {pp116[27]};
    assign in3815_2 = {pp117[26]};
    Full_Adder FA_3815(s3815, c3815, in3815_1, in3815_2, pp115[28]);
    wire[0:0] s3816, in3816_1, in3816_2;
    wire c3816;
    assign in3816_1 = {pp119[24]};
    assign in3816_2 = {pp120[23]};
    Full_Adder FA_3816(s3816, c3816, in3816_1, in3816_2, pp118[25]);
    wire[0:0] s3817, in3817_1, in3817_2;
    wire c3817;
    assign in3817_1 = {pp122[21]};
    assign in3817_2 = {pp123[20]};
    Full_Adder FA_3817(s3817, c3817, in3817_1, in3817_2, pp121[22]);
    wire[0:0] s3818, in3818_1, in3818_2;
    wire c3818;
    assign in3818_1 = {pp125[18]};
    assign in3818_2 = {pp126[17]};
    Full_Adder FA_3818(s3818, c3818, in3818_1, in3818_2, pp124[19]);
    wire[0:0] s3819, in3819_1, in3819_2;
    wire c3819;
    assign in3819_1 = {c1401};
    assign in3819_2 = {c1402};
    Full_Adder FA_3819(s3819, c3819, in3819_1, in3819_2, pp127[16]);
    wire[0:0] s3820, in3820_1, in3820_2;
    wire c3820;
    assign in3820_1 = {c1404};
    assign in3820_2 = {c1405};
    Full_Adder FA_3820(s3820, c3820, in3820_1, in3820_2, c1403);
    wire[0:0] s3821, in3821_1, in3821_2;
    wire c3821;
    assign in3821_1 = {c1407};
    assign in3821_2 = {c1408};
    Full_Adder FA_3821(s3821, c3821, in3821_1, in3821_2, c1406);
    wire[0:0] s3822, in3822_1, in3822_2;
    wire c3822;
    assign in3822_1 = {c1410};
    assign in3822_2 = {c1411};
    Full_Adder FA_3822(s3822, c3822, in3822_1, in3822_2, c1409);
    wire[0:0] s3823, in3823_1, in3823_2;
    wire c3823;
    assign in3823_1 = {c1413};
    assign in3823_2 = {c1414};
    Full_Adder FA_3823(s3823, c3823, in3823_1, in3823_2, c1412);
    wire[0:0] s3824, in3824_1, in3824_2;
    wire c3824;
    assign in3824_1 = {c1416};
    assign in3824_2 = {c1417};
    Full_Adder FA_3824(s3824, c3824, in3824_1, in3824_2, c1415);
    wire[0:0] s3825, in3825_1, in3825_2;
    wire c3825;
    assign in3825_1 = {c1419};
    assign in3825_2 = {c1420};
    Full_Adder FA_3825(s3825, c3825, in3825_1, in3825_2, c1418);
    wire[0:0] s3826, in3826_1, in3826_2;
    wire c3826;
    assign in3826_1 = {c1422};
    assign in3826_2 = {c1423};
    Full_Adder FA_3826(s3826, c3826, in3826_1, in3826_2, c1421);
    wire[0:0] s3827, in3827_1, in3827_2;
    wire c3827;
    assign in3827_1 = {c1425};
    assign in3827_2 = {c1426};
    Full_Adder FA_3827(s3827, c3827, in3827_1, in3827_2, c1424);
    wire[0:0] s3828, in3828_1, in3828_2;
    wire c3828;
    assign in3828_1 = {c1428};
    assign in3828_2 = {s1429[0]};
    Full_Adder FA_3828(s3828, c3828, in3828_1, in3828_2, c1427);
    wire[0:0] s3829, in3829_1, in3829_2;
    wire c3829;
    assign in3829_1 = {s1431[0]};
    assign in3829_2 = {s1432[0]};
    Full_Adder FA_3829(s3829, c3829, in3829_1, in3829_2, s1430[0]);
    wire[0:0] s3830, in3830_1, in3830_2;
    wire c3830;
    assign in3830_1 = {s1434[0]};
    assign in3830_2 = {s1435[0]};
    Full_Adder FA_3830(s3830, c3830, in3830_1, in3830_2, s1433[0]);
    wire[0:0] s3831, in3831_1, in3831_2;
    wire c3831;
    assign in3831_1 = {s1437[0]};
    assign in3831_2 = {s1438[0]};
    Full_Adder FA_3831(s3831, c3831, in3831_1, in3831_2, s1436[0]);
    wire[0:0] s3832, in3832_1, in3832_2;
    wire c3832;
    assign in3832_1 = {s1440[0]};
    assign in3832_2 = {s1441[0]};
    Full_Adder FA_3832(s3832, c3832, in3832_1, in3832_2, s1439[0]);
    wire[0:0] s3833, in3833_1, in3833_2;
    wire c3833;
    assign in3833_1 = {s1443[0]};
    assign in3833_2 = {s1444[0]};
    Full_Adder FA_3833(s3833, c3833, in3833_1, in3833_2, s1442[0]);
    wire[0:0] s3834, in3834_1, in3834_2;
    wire c3834;
    assign in3834_1 = {s1446[0]};
    assign in3834_2 = {s1447[0]};
    Full_Adder FA_3834(s3834, c3834, in3834_1, in3834_2, s1445[0]);
    wire[0:0] s3835, in3835_1, in3835_2;
    wire c3835;
    assign in3835_1 = {s1449[0]};
    assign in3835_2 = {s1450[0]};
    Full_Adder FA_3835(s3835, c3835, in3835_1, in3835_2, s1448[0]);
    wire[0:0] s3836, in3836_1, in3836_2;
    wire c3836;
    assign in3836_1 = {s1452[0]};
    assign in3836_2 = {s1453[0]};
    Full_Adder FA_3836(s3836, c3836, in3836_1, in3836_2, s1451[0]);
    wire[0:0] s3837, in3837_1, in3837_2;
    wire c3837;
    assign in3837_1 = {pp96[48]};
    assign in3837_2 = {pp97[47]};
    Full_Adder FA_3837(s3837, c3837, in3837_1, in3837_2, pp95[49]);
    wire[0:0] s3838, in3838_1, in3838_2;
    wire c3838;
    assign in3838_1 = {pp99[45]};
    assign in3838_2 = {pp100[44]};
    Full_Adder FA_3838(s3838, c3838, in3838_1, in3838_2, pp98[46]);
    wire[0:0] s3839, in3839_1, in3839_2;
    wire c3839;
    assign in3839_1 = {pp102[42]};
    assign in3839_2 = {pp103[41]};
    Full_Adder FA_3839(s3839, c3839, in3839_1, in3839_2, pp101[43]);
    wire[0:0] s3840, in3840_1, in3840_2;
    wire c3840;
    assign in3840_1 = {pp105[39]};
    assign in3840_2 = {pp106[38]};
    Full_Adder FA_3840(s3840, c3840, in3840_1, in3840_2, pp104[40]);
    wire[0:0] s3841, in3841_1, in3841_2;
    wire c3841;
    assign in3841_1 = {pp108[36]};
    assign in3841_2 = {pp109[35]};
    Full_Adder FA_3841(s3841, c3841, in3841_1, in3841_2, pp107[37]);
    wire[0:0] s3842, in3842_1, in3842_2;
    wire c3842;
    assign in3842_1 = {pp111[33]};
    assign in3842_2 = {pp112[32]};
    Full_Adder FA_3842(s3842, c3842, in3842_1, in3842_2, pp110[34]);
    wire[0:0] s3843, in3843_1, in3843_2;
    wire c3843;
    assign in3843_1 = {pp114[30]};
    assign in3843_2 = {pp115[29]};
    Full_Adder FA_3843(s3843, c3843, in3843_1, in3843_2, pp113[31]);
    wire[0:0] s3844, in3844_1, in3844_2;
    wire c3844;
    assign in3844_1 = {pp117[27]};
    assign in3844_2 = {pp118[26]};
    Full_Adder FA_3844(s3844, c3844, in3844_1, in3844_2, pp116[28]);
    wire[0:0] s3845, in3845_1, in3845_2;
    wire c3845;
    assign in3845_1 = {pp120[24]};
    assign in3845_2 = {pp121[23]};
    Full_Adder FA_3845(s3845, c3845, in3845_1, in3845_2, pp119[25]);
    wire[0:0] s3846, in3846_1, in3846_2;
    wire c3846;
    assign in3846_1 = {pp123[21]};
    assign in3846_2 = {pp124[20]};
    Full_Adder FA_3846(s3846, c3846, in3846_1, in3846_2, pp122[22]);
    wire[0:0] s3847, in3847_1, in3847_2;
    wire c3847;
    assign in3847_1 = {pp126[18]};
    assign in3847_2 = {pp127[17]};
    Full_Adder FA_3847(s3847, c3847, in3847_1, in3847_2, pp125[19]);
    wire[0:0] s3848, in3848_1, in3848_2;
    wire c3848;
    assign in3848_1 = {c1430};
    assign in3848_2 = {c1431};
    Full_Adder FA_3848(s3848, c3848, in3848_1, in3848_2, c1429);
    wire[0:0] s3849, in3849_1, in3849_2;
    wire c3849;
    assign in3849_1 = {c1433};
    assign in3849_2 = {c1434};
    Full_Adder FA_3849(s3849, c3849, in3849_1, in3849_2, c1432);
    wire[0:0] s3850, in3850_1, in3850_2;
    wire c3850;
    assign in3850_1 = {c1436};
    assign in3850_2 = {c1437};
    Full_Adder FA_3850(s3850, c3850, in3850_1, in3850_2, c1435);
    wire[0:0] s3851, in3851_1, in3851_2;
    wire c3851;
    assign in3851_1 = {c1439};
    assign in3851_2 = {c1440};
    Full_Adder FA_3851(s3851, c3851, in3851_1, in3851_2, c1438);
    wire[0:0] s3852, in3852_1, in3852_2;
    wire c3852;
    assign in3852_1 = {c1442};
    assign in3852_2 = {c1443};
    Full_Adder FA_3852(s3852, c3852, in3852_1, in3852_2, c1441);
    wire[0:0] s3853, in3853_1, in3853_2;
    wire c3853;
    assign in3853_1 = {c1445};
    assign in3853_2 = {c1446};
    Full_Adder FA_3853(s3853, c3853, in3853_1, in3853_2, c1444);
    wire[0:0] s3854, in3854_1, in3854_2;
    wire c3854;
    assign in3854_1 = {c1448};
    assign in3854_2 = {c1449};
    Full_Adder FA_3854(s3854, c3854, in3854_1, in3854_2, c1447);
    wire[0:0] s3855, in3855_1, in3855_2;
    wire c3855;
    assign in3855_1 = {c1451};
    assign in3855_2 = {c1452};
    Full_Adder FA_3855(s3855, c3855, in3855_1, in3855_2, c1450);
    wire[0:0] s3856, in3856_1, in3856_2;
    wire c3856;
    assign in3856_1 = {c1454};
    assign in3856_2 = {c1455};
    Full_Adder FA_3856(s3856, c3856, in3856_1, in3856_2, c1453);
    wire[0:0] s3857, in3857_1, in3857_2;
    wire c3857;
    assign in3857_1 = {s1457[0]};
    assign in3857_2 = {s1458[0]};
    Full_Adder FA_3857(s3857, c3857, in3857_1, in3857_2, s1456[0]);
    wire[0:0] s3858, in3858_1, in3858_2;
    wire c3858;
    assign in3858_1 = {s1460[0]};
    assign in3858_2 = {s1461[0]};
    Full_Adder FA_3858(s3858, c3858, in3858_1, in3858_2, s1459[0]);
    wire[0:0] s3859, in3859_1, in3859_2;
    wire c3859;
    assign in3859_1 = {s1463[0]};
    assign in3859_2 = {s1464[0]};
    Full_Adder FA_3859(s3859, c3859, in3859_1, in3859_2, s1462[0]);
    wire[0:0] s3860, in3860_1, in3860_2;
    wire c3860;
    assign in3860_1 = {s1466[0]};
    assign in3860_2 = {s1467[0]};
    Full_Adder FA_3860(s3860, c3860, in3860_1, in3860_2, s1465[0]);
    wire[0:0] s3861, in3861_1, in3861_2;
    wire c3861;
    assign in3861_1 = {s1469[0]};
    assign in3861_2 = {s1470[0]};
    Full_Adder FA_3861(s3861, c3861, in3861_1, in3861_2, s1468[0]);
    wire[0:0] s3862, in3862_1, in3862_2;
    wire c3862;
    assign in3862_1 = {s1472[0]};
    assign in3862_2 = {s1473[0]};
    Full_Adder FA_3862(s3862, c3862, in3862_1, in3862_2, s1471[0]);
    wire[0:0] s3863, in3863_1, in3863_2;
    wire c3863;
    assign in3863_1 = {s1475[0]};
    assign in3863_2 = {s1476[0]};
    Full_Adder FA_3863(s3863, c3863, in3863_1, in3863_2, s1474[0]);
    wire[0:0] s3864, in3864_1, in3864_2;
    wire c3864;
    assign in3864_1 = {s1478[0]};
    assign in3864_2 = {s1479[0]};
    Full_Adder FA_3864(s3864, c3864, in3864_1, in3864_2, s1477[0]);
    wire[0:0] s3865, in3865_1, in3865_2;
    wire c3865;
    assign in3865_1 = {pp94[51]};
    assign in3865_2 = {pp95[50]};
    Full_Adder FA_3865(s3865, c3865, in3865_1, in3865_2, pp93[52]);
    wire[0:0] s3866, in3866_1, in3866_2;
    wire c3866;
    assign in3866_1 = {pp97[48]};
    assign in3866_2 = {pp98[47]};
    Full_Adder FA_3866(s3866, c3866, in3866_1, in3866_2, pp96[49]);
    wire[0:0] s3867, in3867_1, in3867_2;
    wire c3867;
    assign in3867_1 = {pp100[45]};
    assign in3867_2 = {pp101[44]};
    Full_Adder FA_3867(s3867, c3867, in3867_1, in3867_2, pp99[46]);
    wire[0:0] s3868, in3868_1, in3868_2;
    wire c3868;
    assign in3868_1 = {pp103[42]};
    assign in3868_2 = {pp104[41]};
    Full_Adder FA_3868(s3868, c3868, in3868_1, in3868_2, pp102[43]);
    wire[0:0] s3869, in3869_1, in3869_2;
    wire c3869;
    assign in3869_1 = {pp106[39]};
    assign in3869_2 = {pp107[38]};
    Full_Adder FA_3869(s3869, c3869, in3869_1, in3869_2, pp105[40]);
    wire[0:0] s3870, in3870_1, in3870_2;
    wire c3870;
    assign in3870_1 = {pp109[36]};
    assign in3870_2 = {pp110[35]};
    Full_Adder FA_3870(s3870, c3870, in3870_1, in3870_2, pp108[37]);
    wire[0:0] s3871, in3871_1, in3871_2;
    wire c3871;
    assign in3871_1 = {pp112[33]};
    assign in3871_2 = {pp113[32]};
    Full_Adder FA_3871(s3871, c3871, in3871_1, in3871_2, pp111[34]);
    wire[0:0] s3872, in3872_1, in3872_2;
    wire c3872;
    assign in3872_1 = {pp115[30]};
    assign in3872_2 = {pp116[29]};
    Full_Adder FA_3872(s3872, c3872, in3872_1, in3872_2, pp114[31]);
    wire[0:0] s3873, in3873_1, in3873_2;
    wire c3873;
    assign in3873_1 = {pp118[27]};
    assign in3873_2 = {pp119[26]};
    Full_Adder FA_3873(s3873, c3873, in3873_1, in3873_2, pp117[28]);
    wire[0:0] s3874, in3874_1, in3874_2;
    wire c3874;
    assign in3874_1 = {pp121[24]};
    assign in3874_2 = {pp122[23]};
    Full_Adder FA_3874(s3874, c3874, in3874_1, in3874_2, pp120[25]);
    wire[0:0] s3875, in3875_1, in3875_2;
    wire c3875;
    assign in3875_1 = {pp124[21]};
    assign in3875_2 = {pp125[20]};
    Full_Adder FA_3875(s3875, c3875, in3875_1, in3875_2, pp123[22]);
    wire[0:0] s3876, in3876_1, in3876_2;
    wire c3876;
    assign in3876_1 = {pp127[18]};
    assign in3876_2 = {c1456};
    Full_Adder FA_3876(s3876, c3876, in3876_1, in3876_2, pp126[19]);
    wire[0:0] s3877, in3877_1, in3877_2;
    wire c3877;
    assign in3877_1 = {c1458};
    assign in3877_2 = {c1459};
    Full_Adder FA_3877(s3877, c3877, in3877_1, in3877_2, c1457);
    wire[0:0] s3878, in3878_1, in3878_2;
    wire c3878;
    assign in3878_1 = {c1461};
    assign in3878_2 = {c1462};
    Full_Adder FA_3878(s3878, c3878, in3878_1, in3878_2, c1460);
    wire[0:0] s3879, in3879_1, in3879_2;
    wire c3879;
    assign in3879_1 = {c1464};
    assign in3879_2 = {c1465};
    Full_Adder FA_3879(s3879, c3879, in3879_1, in3879_2, c1463);
    wire[0:0] s3880, in3880_1, in3880_2;
    wire c3880;
    assign in3880_1 = {c1467};
    assign in3880_2 = {c1468};
    Full_Adder FA_3880(s3880, c3880, in3880_1, in3880_2, c1466);
    wire[0:0] s3881, in3881_1, in3881_2;
    wire c3881;
    assign in3881_1 = {c1470};
    assign in3881_2 = {c1471};
    Full_Adder FA_3881(s3881, c3881, in3881_1, in3881_2, c1469);
    wire[0:0] s3882, in3882_1, in3882_2;
    wire c3882;
    assign in3882_1 = {c1473};
    assign in3882_2 = {c1474};
    Full_Adder FA_3882(s3882, c3882, in3882_1, in3882_2, c1472);
    wire[0:0] s3883, in3883_1, in3883_2;
    wire c3883;
    assign in3883_1 = {c1476};
    assign in3883_2 = {c1477};
    Full_Adder FA_3883(s3883, c3883, in3883_1, in3883_2, c1475);
    wire[0:0] s3884, in3884_1, in3884_2;
    wire c3884;
    assign in3884_1 = {c1479};
    assign in3884_2 = {c1480};
    Full_Adder FA_3884(s3884, c3884, in3884_1, in3884_2, c1478);
    wire[0:0] s3885, in3885_1, in3885_2;
    wire c3885;
    assign in3885_1 = {s1482[0]};
    assign in3885_2 = {s1483[0]};
    Full_Adder FA_3885(s3885, c3885, in3885_1, in3885_2, c1481);
    wire[0:0] s3886, in3886_1, in3886_2;
    wire c3886;
    assign in3886_1 = {s1485[0]};
    assign in3886_2 = {s1486[0]};
    Full_Adder FA_3886(s3886, c3886, in3886_1, in3886_2, s1484[0]);
    wire[0:0] s3887, in3887_1, in3887_2;
    wire c3887;
    assign in3887_1 = {s1488[0]};
    assign in3887_2 = {s1489[0]};
    Full_Adder FA_3887(s3887, c3887, in3887_1, in3887_2, s1487[0]);
    wire[0:0] s3888, in3888_1, in3888_2;
    wire c3888;
    assign in3888_1 = {s1491[0]};
    assign in3888_2 = {s1492[0]};
    Full_Adder FA_3888(s3888, c3888, in3888_1, in3888_2, s1490[0]);
    wire[0:0] s3889, in3889_1, in3889_2;
    wire c3889;
    assign in3889_1 = {s1494[0]};
    assign in3889_2 = {s1495[0]};
    Full_Adder FA_3889(s3889, c3889, in3889_1, in3889_2, s1493[0]);
    wire[0:0] s3890, in3890_1, in3890_2;
    wire c3890;
    assign in3890_1 = {s1497[0]};
    assign in3890_2 = {s1498[0]};
    Full_Adder FA_3890(s3890, c3890, in3890_1, in3890_2, s1496[0]);
    wire[0:0] s3891, in3891_1, in3891_2;
    wire c3891;
    assign in3891_1 = {s1500[0]};
    assign in3891_2 = {s1501[0]};
    Full_Adder FA_3891(s3891, c3891, in3891_1, in3891_2, s1499[0]);
    wire[0:0] s3892, in3892_1, in3892_2;
    wire c3892;
    assign in3892_1 = {s1503[0]};
    assign in3892_2 = {s1504[0]};
    Full_Adder FA_3892(s3892, c3892, in3892_1, in3892_2, s1502[0]);
    wire[0:0] s3893, in3893_1, in3893_2;
    wire c3893;
    assign in3893_1 = {pp92[54]};
    assign in3893_2 = {pp93[53]};
    Full_Adder FA_3893(s3893, c3893, in3893_1, in3893_2, pp91[55]);
    wire[0:0] s3894, in3894_1, in3894_2;
    wire c3894;
    assign in3894_1 = {pp95[51]};
    assign in3894_2 = {pp96[50]};
    Full_Adder FA_3894(s3894, c3894, in3894_1, in3894_2, pp94[52]);
    wire[0:0] s3895, in3895_1, in3895_2;
    wire c3895;
    assign in3895_1 = {pp98[48]};
    assign in3895_2 = {pp99[47]};
    Full_Adder FA_3895(s3895, c3895, in3895_1, in3895_2, pp97[49]);
    wire[0:0] s3896, in3896_1, in3896_2;
    wire c3896;
    assign in3896_1 = {pp101[45]};
    assign in3896_2 = {pp102[44]};
    Full_Adder FA_3896(s3896, c3896, in3896_1, in3896_2, pp100[46]);
    wire[0:0] s3897, in3897_1, in3897_2;
    wire c3897;
    assign in3897_1 = {pp104[42]};
    assign in3897_2 = {pp105[41]};
    Full_Adder FA_3897(s3897, c3897, in3897_1, in3897_2, pp103[43]);
    wire[0:0] s3898, in3898_1, in3898_2;
    wire c3898;
    assign in3898_1 = {pp107[39]};
    assign in3898_2 = {pp108[38]};
    Full_Adder FA_3898(s3898, c3898, in3898_1, in3898_2, pp106[40]);
    wire[0:0] s3899, in3899_1, in3899_2;
    wire c3899;
    assign in3899_1 = {pp110[36]};
    assign in3899_2 = {pp111[35]};
    Full_Adder FA_3899(s3899, c3899, in3899_1, in3899_2, pp109[37]);
    wire[0:0] s3900, in3900_1, in3900_2;
    wire c3900;
    assign in3900_1 = {pp113[33]};
    assign in3900_2 = {pp114[32]};
    Full_Adder FA_3900(s3900, c3900, in3900_1, in3900_2, pp112[34]);
    wire[0:0] s3901, in3901_1, in3901_2;
    wire c3901;
    assign in3901_1 = {pp116[30]};
    assign in3901_2 = {pp117[29]};
    Full_Adder FA_3901(s3901, c3901, in3901_1, in3901_2, pp115[31]);
    wire[0:0] s3902, in3902_1, in3902_2;
    wire c3902;
    assign in3902_1 = {pp119[27]};
    assign in3902_2 = {pp120[26]};
    Full_Adder FA_3902(s3902, c3902, in3902_1, in3902_2, pp118[28]);
    wire[0:0] s3903, in3903_1, in3903_2;
    wire c3903;
    assign in3903_1 = {pp122[24]};
    assign in3903_2 = {pp123[23]};
    Full_Adder FA_3903(s3903, c3903, in3903_1, in3903_2, pp121[25]);
    wire[0:0] s3904, in3904_1, in3904_2;
    wire c3904;
    assign in3904_1 = {pp125[21]};
    assign in3904_2 = {pp126[20]};
    Full_Adder FA_3904(s3904, c3904, in3904_1, in3904_2, pp124[22]);
    wire[0:0] s3905, in3905_1, in3905_2;
    wire c3905;
    assign in3905_1 = {c1482};
    assign in3905_2 = {c1483};
    Full_Adder FA_3905(s3905, c3905, in3905_1, in3905_2, pp127[19]);
    wire[0:0] s3906, in3906_1, in3906_2;
    wire c3906;
    assign in3906_1 = {c1485};
    assign in3906_2 = {c1486};
    Full_Adder FA_3906(s3906, c3906, in3906_1, in3906_2, c1484);
    wire[0:0] s3907, in3907_1, in3907_2;
    wire c3907;
    assign in3907_1 = {c1488};
    assign in3907_2 = {c1489};
    Full_Adder FA_3907(s3907, c3907, in3907_1, in3907_2, c1487);
    wire[0:0] s3908, in3908_1, in3908_2;
    wire c3908;
    assign in3908_1 = {c1491};
    assign in3908_2 = {c1492};
    Full_Adder FA_3908(s3908, c3908, in3908_1, in3908_2, c1490);
    wire[0:0] s3909, in3909_1, in3909_2;
    wire c3909;
    assign in3909_1 = {c1494};
    assign in3909_2 = {c1495};
    Full_Adder FA_3909(s3909, c3909, in3909_1, in3909_2, c1493);
    wire[0:0] s3910, in3910_1, in3910_2;
    wire c3910;
    assign in3910_1 = {c1497};
    assign in3910_2 = {c1498};
    Full_Adder FA_3910(s3910, c3910, in3910_1, in3910_2, c1496);
    wire[0:0] s3911, in3911_1, in3911_2;
    wire c3911;
    assign in3911_1 = {c1500};
    assign in3911_2 = {c1501};
    Full_Adder FA_3911(s3911, c3911, in3911_1, in3911_2, c1499);
    wire[0:0] s3912, in3912_1, in3912_2;
    wire c3912;
    assign in3912_1 = {c1503};
    assign in3912_2 = {c1504};
    Full_Adder FA_3912(s3912, c3912, in3912_1, in3912_2, c1502);
    wire[0:0] s3913, in3913_1, in3913_2;
    wire c3913;
    assign in3913_1 = {c1506};
    assign in3913_2 = {s1507[0]};
    Full_Adder FA_3913(s3913, c3913, in3913_1, in3913_2, c1505);
    wire[0:0] s3914, in3914_1, in3914_2;
    wire c3914;
    assign in3914_1 = {s1509[0]};
    assign in3914_2 = {s1510[0]};
    Full_Adder FA_3914(s3914, c3914, in3914_1, in3914_2, s1508[0]);
    wire[0:0] s3915, in3915_1, in3915_2;
    wire c3915;
    assign in3915_1 = {s1512[0]};
    assign in3915_2 = {s1513[0]};
    Full_Adder FA_3915(s3915, c3915, in3915_1, in3915_2, s1511[0]);
    wire[0:0] s3916, in3916_1, in3916_2;
    wire c3916;
    assign in3916_1 = {s1515[0]};
    assign in3916_2 = {s1516[0]};
    Full_Adder FA_3916(s3916, c3916, in3916_1, in3916_2, s1514[0]);
    wire[0:0] s3917, in3917_1, in3917_2;
    wire c3917;
    assign in3917_1 = {s1518[0]};
    assign in3917_2 = {s1519[0]};
    Full_Adder FA_3917(s3917, c3917, in3917_1, in3917_2, s1517[0]);
    wire[0:0] s3918, in3918_1, in3918_2;
    wire c3918;
    assign in3918_1 = {s1521[0]};
    assign in3918_2 = {s1522[0]};
    Full_Adder FA_3918(s3918, c3918, in3918_1, in3918_2, s1520[0]);
    wire[0:0] s3919, in3919_1, in3919_2;
    wire c3919;
    assign in3919_1 = {s1524[0]};
    assign in3919_2 = {s1525[0]};
    Full_Adder FA_3919(s3919, c3919, in3919_1, in3919_2, s1523[0]);
    wire[0:0] s3920, in3920_1, in3920_2;
    wire c3920;
    assign in3920_1 = {s1527[0]};
    assign in3920_2 = {s1528[0]};
    Full_Adder FA_3920(s3920, c3920, in3920_1, in3920_2, s1526[0]);
    wire[0:0] s3921, in3921_1, in3921_2;
    wire c3921;
    assign in3921_1 = {pp90[57]};
    assign in3921_2 = {pp91[56]};
    Full_Adder FA_3921(s3921, c3921, in3921_1, in3921_2, pp89[58]);
    wire[0:0] s3922, in3922_1, in3922_2;
    wire c3922;
    assign in3922_1 = {pp93[54]};
    assign in3922_2 = {pp94[53]};
    Full_Adder FA_3922(s3922, c3922, in3922_1, in3922_2, pp92[55]);
    wire[0:0] s3923, in3923_1, in3923_2;
    wire c3923;
    assign in3923_1 = {pp96[51]};
    assign in3923_2 = {pp97[50]};
    Full_Adder FA_3923(s3923, c3923, in3923_1, in3923_2, pp95[52]);
    wire[0:0] s3924, in3924_1, in3924_2;
    wire c3924;
    assign in3924_1 = {pp99[48]};
    assign in3924_2 = {pp100[47]};
    Full_Adder FA_3924(s3924, c3924, in3924_1, in3924_2, pp98[49]);
    wire[0:0] s3925, in3925_1, in3925_2;
    wire c3925;
    assign in3925_1 = {pp102[45]};
    assign in3925_2 = {pp103[44]};
    Full_Adder FA_3925(s3925, c3925, in3925_1, in3925_2, pp101[46]);
    wire[0:0] s3926, in3926_1, in3926_2;
    wire c3926;
    assign in3926_1 = {pp105[42]};
    assign in3926_2 = {pp106[41]};
    Full_Adder FA_3926(s3926, c3926, in3926_1, in3926_2, pp104[43]);
    wire[0:0] s3927, in3927_1, in3927_2;
    wire c3927;
    assign in3927_1 = {pp108[39]};
    assign in3927_2 = {pp109[38]};
    Full_Adder FA_3927(s3927, c3927, in3927_1, in3927_2, pp107[40]);
    wire[0:0] s3928, in3928_1, in3928_2;
    wire c3928;
    assign in3928_1 = {pp111[36]};
    assign in3928_2 = {pp112[35]};
    Full_Adder FA_3928(s3928, c3928, in3928_1, in3928_2, pp110[37]);
    wire[0:0] s3929, in3929_1, in3929_2;
    wire c3929;
    assign in3929_1 = {pp114[33]};
    assign in3929_2 = {pp115[32]};
    Full_Adder FA_3929(s3929, c3929, in3929_1, in3929_2, pp113[34]);
    wire[0:0] s3930, in3930_1, in3930_2;
    wire c3930;
    assign in3930_1 = {pp117[30]};
    assign in3930_2 = {pp118[29]};
    Full_Adder FA_3930(s3930, c3930, in3930_1, in3930_2, pp116[31]);
    wire[0:0] s3931, in3931_1, in3931_2;
    wire c3931;
    assign in3931_1 = {pp120[27]};
    assign in3931_2 = {pp121[26]};
    Full_Adder FA_3931(s3931, c3931, in3931_1, in3931_2, pp119[28]);
    wire[0:0] s3932, in3932_1, in3932_2;
    wire c3932;
    assign in3932_1 = {pp123[24]};
    assign in3932_2 = {pp124[23]};
    Full_Adder FA_3932(s3932, c3932, in3932_1, in3932_2, pp122[25]);
    wire[0:0] s3933, in3933_1, in3933_2;
    wire c3933;
    assign in3933_1 = {pp126[21]};
    assign in3933_2 = {pp127[20]};
    Full_Adder FA_3933(s3933, c3933, in3933_1, in3933_2, pp125[22]);
    wire[0:0] s3934, in3934_1, in3934_2;
    wire c3934;
    assign in3934_1 = {c1508};
    assign in3934_2 = {c1509};
    Full_Adder FA_3934(s3934, c3934, in3934_1, in3934_2, c1507);
    wire[0:0] s3935, in3935_1, in3935_2;
    wire c3935;
    assign in3935_1 = {c1511};
    assign in3935_2 = {c1512};
    Full_Adder FA_3935(s3935, c3935, in3935_1, in3935_2, c1510);
    wire[0:0] s3936, in3936_1, in3936_2;
    wire c3936;
    assign in3936_1 = {c1514};
    assign in3936_2 = {c1515};
    Full_Adder FA_3936(s3936, c3936, in3936_1, in3936_2, c1513);
    wire[0:0] s3937, in3937_1, in3937_2;
    wire c3937;
    assign in3937_1 = {c1517};
    assign in3937_2 = {c1518};
    Full_Adder FA_3937(s3937, c3937, in3937_1, in3937_2, c1516);
    wire[0:0] s3938, in3938_1, in3938_2;
    wire c3938;
    assign in3938_1 = {c1520};
    assign in3938_2 = {c1521};
    Full_Adder FA_3938(s3938, c3938, in3938_1, in3938_2, c1519);
    wire[0:0] s3939, in3939_1, in3939_2;
    wire c3939;
    assign in3939_1 = {c1523};
    assign in3939_2 = {c1524};
    Full_Adder FA_3939(s3939, c3939, in3939_1, in3939_2, c1522);
    wire[0:0] s3940, in3940_1, in3940_2;
    wire c3940;
    assign in3940_1 = {c1526};
    assign in3940_2 = {c1527};
    Full_Adder FA_3940(s3940, c3940, in3940_1, in3940_2, c1525);
    wire[0:0] s3941, in3941_1, in3941_2;
    wire c3941;
    assign in3941_1 = {c1529};
    assign in3941_2 = {c1530};
    Full_Adder FA_3941(s3941, c3941, in3941_1, in3941_2, c1528);
    wire[0:0] s3942, in3942_1, in3942_2;
    wire c3942;
    assign in3942_1 = {s1532[0]};
    assign in3942_2 = {s1533[0]};
    Full_Adder FA_3942(s3942, c3942, in3942_1, in3942_2, s1531[0]);
    wire[0:0] s3943, in3943_1, in3943_2;
    wire c3943;
    assign in3943_1 = {s1535[0]};
    assign in3943_2 = {s1536[0]};
    Full_Adder FA_3943(s3943, c3943, in3943_1, in3943_2, s1534[0]);
    wire[0:0] s3944, in3944_1, in3944_2;
    wire c3944;
    assign in3944_1 = {s1538[0]};
    assign in3944_2 = {s1539[0]};
    Full_Adder FA_3944(s3944, c3944, in3944_1, in3944_2, s1537[0]);
    wire[0:0] s3945, in3945_1, in3945_2;
    wire c3945;
    assign in3945_1 = {s1541[0]};
    assign in3945_2 = {s1542[0]};
    Full_Adder FA_3945(s3945, c3945, in3945_1, in3945_2, s1540[0]);
    wire[0:0] s3946, in3946_1, in3946_2;
    wire c3946;
    assign in3946_1 = {s1544[0]};
    assign in3946_2 = {s1545[0]};
    Full_Adder FA_3946(s3946, c3946, in3946_1, in3946_2, s1543[0]);
    wire[0:0] s3947, in3947_1, in3947_2;
    wire c3947;
    assign in3947_1 = {s1547[0]};
    assign in3947_2 = {s1548[0]};
    Full_Adder FA_3947(s3947, c3947, in3947_1, in3947_2, s1546[0]);
    wire[0:0] s3948, in3948_1, in3948_2;
    wire c3948;
    assign in3948_1 = {s1550[0]};
    assign in3948_2 = {s1551[0]};
    Full_Adder FA_3948(s3948, c3948, in3948_1, in3948_2, s1549[0]);
    wire[0:0] s3949, in3949_1, in3949_2;
    wire c3949;
    assign in3949_1 = {pp88[60]};
    assign in3949_2 = {pp89[59]};
    Full_Adder FA_3949(s3949, c3949, in3949_1, in3949_2, pp87[61]);
    wire[0:0] s3950, in3950_1, in3950_2;
    wire c3950;
    assign in3950_1 = {pp91[57]};
    assign in3950_2 = {pp92[56]};
    Full_Adder FA_3950(s3950, c3950, in3950_1, in3950_2, pp90[58]);
    wire[0:0] s3951, in3951_1, in3951_2;
    wire c3951;
    assign in3951_1 = {pp94[54]};
    assign in3951_2 = {pp95[53]};
    Full_Adder FA_3951(s3951, c3951, in3951_1, in3951_2, pp93[55]);
    wire[0:0] s3952, in3952_1, in3952_2;
    wire c3952;
    assign in3952_1 = {pp97[51]};
    assign in3952_2 = {pp98[50]};
    Full_Adder FA_3952(s3952, c3952, in3952_1, in3952_2, pp96[52]);
    wire[0:0] s3953, in3953_1, in3953_2;
    wire c3953;
    assign in3953_1 = {pp100[48]};
    assign in3953_2 = {pp101[47]};
    Full_Adder FA_3953(s3953, c3953, in3953_1, in3953_2, pp99[49]);
    wire[0:0] s3954, in3954_1, in3954_2;
    wire c3954;
    assign in3954_1 = {pp103[45]};
    assign in3954_2 = {pp104[44]};
    Full_Adder FA_3954(s3954, c3954, in3954_1, in3954_2, pp102[46]);
    wire[0:0] s3955, in3955_1, in3955_2;
    wire c3955;
    assign in3955_1 = {pp106[42]};
    assign in3955_2 = {pp107[41]};
    Full_Adder FA_3955(s3955, c3955, in3955_1, in3955_2, pp105[43]);
    wire[0:0] s3956, in3956_1, in3956_2;
    wire c3956;
    assign in3956_1 = {pp109[39]};
    assign in3956_2 = {pp110[38]};
    Full_Adder FA_3956(s3956, c3956, in3956_1, in3956_2, pp108[40]);
    wire[0:0] s3957, in3957_1, in3957_2;
    wire c3957;
    assign in3957_1 = {pp112[36]};
    assign in3957_2 = {pp113[35]};
    Full_Adder FA_3957(s3957, c3957, in3957_1, in3957_2, pp111[37]);
    wire[0:0] s3958, in3958_1, in3958_2;
    wire c3958;
    assign in3958_1 = {pp115[33]};
    assign in3958_2 = {pp116[32]};
    Full_Adder FA_3958(s3958, c3958, in3958_1, in3958_2, pp114[34]);
    wire[0:0] s3959, in3959_1, in3959_2;
    wire c3959;
    assign in3959_1 = {pp118[30]};
    assign in3959_2 = {pp119[29]};
    Full_Adder FA_3959(s3959, c3959, in3959_1, in3959_2, pp117[31]);
    wire[0:0] s3960, in3960_1, in3960_2;
    wire c3960;
    assign in3960_1 = {pp121[27]};
    assign in3960_2 = {pp122[26]};
    Full_Adder FA_3960(s3960, c3960, in3960_1, in3960_2, pp120[28]);
    wire[0:0] s3961, in3961_1, in3961_2;
    wire c3961;
    assign in3961_1 = {pp124[24]};
    assign in3961_2 = {pp125[23]};
    Full_Adder FA_3961(s3961, c3961, in3961_1, in3961_2, pp123[25]);
    wire[0:0] s3962, in3962_1, in3962_2;
    wire c3962;
    assign in3962_1 = {pp127[21]};
    assign in3962_2 = {c1531};
    Full_Adder FA_3962(s3962, c3962, in3962_1, in3962_2, pp126[22]);
    wire[0:0] s3963, in3963_1, in3963_2;
    wire c3963;
    assign in3963_1 = {c1533};
    assign in3963_2 = {c1534};
    Full_Adder FA_3963(s3963, c3963, in3963_1, in3963_2, c1532);
    wire[0:0] s3964, in3964_1, in3964_2;
    wire c3964;
    assign in3964_1 = {c1536};
    assign in3964_2 = {c1537};
    Full_Adder FA_3964(s3964, c3964, in3964_1, in3964_2, c1535);
    wire[0:0] s3965, in3965_1, in3965_2;
    wire c3965;
    assign in3965_1 = {c1539};
    assign in3965_2 = {c1540};
    Full_Adder FA_3965(s3965, c3965, in3965_1, in3965_2, c1538);
    wire[0:0] s3966, in3966_1, in3966_2;
    wire c3966;
    assign in3966_1 = {c1542};
    assign in3966_2 = {c1543};
    Full_Adder FA_3966(s3966, c3966, in3966_1, in3966_2, c1541);
    wire[0:0] s3967, in3967_1, in3967_2;
    wire c3967;
    assign in3967_1 = {c1545};
    assign in3967_2 = {c1546};
    Full_Adder FA_3967(s3967, c3967, in3967_1, in3967_2, c1544);
    wire[0:0] s3968, in3968_1, in3968_2;
    wire c3968;
    assign in3968_1 = {c1548};
    assign in3968_2 = {c1549};
    Full_Adder FA_3968(s3968, c3968, in3968_1, in3968_2, c1547);
    wire[0:0] s3969, in3969_1, in3969_2;
    wire c3969;
    assign in3969_1 = {c1551};
    assign in3969_2 = {c1552};
    Full_Adder FA_3969(s3969, c3969, in3969_1, in3969_2, c1550);
    wire[0:0] s3970, in3970_1, in3970_2;
    wire c3970;
    assign in3970_1 = {s1554[0]};
    assign in3970_2 = {s1555[0]};
    Full_Adder FA_3970(s3970, c3970, in3970_1, in3970_2, c1553);
    wire[0:0] s3971, in3971_1, in3971_2;
    wire c3971;
    assign in3971_1 = {s1557[0]};
    assign in3971_2 = {s1558[0]};
    Full_Adder FA_3971(s3971, c3971, in3971_1, in3971_2, s1556[0]);
    wire[0:0] s3972, in3972_1, in3972_2;
    wire c3972;
    assign in3972_1 = {s1560[0]};
    assign in3972_2 = {s1561[0]};
    Full_Adder FA_3972(s3972, c3972, in3972_1, in3972_2, s1559[0]);
    wire[0:0] s3973, in3973_1, in3973_2;
    wire c3973;
    assign in3973_1 = {s1563[0]};
    assign in3973_2 = {s1564[0]};
    Full_Adder FA_3973(s3973, c3973, in3973_1, in3973_2, s1562[0]);
    wire[0:0] s3974, in3974_1, in3974_2;
    wire c3974;
    assign in3974_1 = {s1566[0]};
    assign in3974_2 = {s1567[0]};
    Full_Adder FA_3974(s3974, c3974, in3974_1, in3974_2, s1565[0]);
    wire[0:0] s3975, in3975_1, in3975_2;
    wire c3975;
    assign in3975_1 = {s1569[0]};
    assign in3975_2 = {s1570[0]};
    Full_Adder FA_3975(s3975, c3975, in3975_1, in3975_2, s1568[0]);
    wire[0:0] s3976, in3976_1, in3976_2;
    wire c3976;
    assign in3976_1 = {s1572[0]};
    assign in3976_2 = {s1573[0]};
    Full_Adder FA_3976(s3976, c3976, in3976_1, in3976_2, s1571[0]);
    wire[0:0] s3977, in3977_1, in3977_2;
    wire c3977;
    assign in3977_1 = {pp86[63]};
    assign in3977_2 = {pp87[62]};
    Full_Adder FA_3977(s3977, c3977, in3977_1, in3977_2, pp85[64]);
    wire[0:0] s3978, in3978_1, in3978_2;
    wire c3978;
    assign in3978_1 = {pp89[60]};
    assign in3978_2 = {pp90[59]};
    Full_Adder FA_3978(s3978, c3978, in3978_1, in3978_2, pp88[61]);
    wire[0:0] s3979, in3979_1, in3979_2;
    wire c3979;
    assign in3979_1 = {pp92[57]};
    assign in3979_2 = {pp93[56]};
    Full_Adder FA_3979(s3979, c3979, in3979_1, in3979_2, pp91[58]);
    wire[0:0] s3980, in3980_1, in3980_2;
    wire c3980;
    assign in3980_1 = {pp95[54]};
    assign in3980_2 = {pp96[53]};
    Full_Adder FA_3980(s3980, c3980, in3980_1, in3980_2, pp94[55]);
    wire[0:0] s3981, in3981_1, in3981_2;
    wire c3981;
    assign in3981_1 = {pp98[51]};
    assign in3981_2 = {pp99[50]};
    Full_Adder FA_3981(s3981, c3981, in3981_1, in3981_2, pp97[52]);
    wire[0:0] s3982, in3982_1, in3982_2;
    wire c3982;
    assign in3982_1 = {pp101[48]};
    assign in3982_2 = {pp102[47]};
    Full_Adder FA_3982(s3982, c3982, in3982_1, in3982_2, pp100[49]);
    wire[0:0] s3983, in3983_1, in3983_2;
    wire c3983;
    assign in3983_1 = {pp104[45]};
    assign in3983_2 = {pp105[44]};
    Full_Adder FA_3983(s3983, c3983, in3983_1, in3983_2, pp103[46]);
    wire[0:0] s3984, in3984_1, in3984_2;
    wire c3984;
    assign in3984_1 = {pp107[42]};
    assign in3984_2 = {pp108[41]};
    Full_Adder FA_3984(s3984, c3984, in3984_1, in3984_2, pp106[43]);
    wire[0:0] s3985, in3985_1, in3985_2;
    wire c3985;
    assign in3985_1 = {pp110[39]};
    assign in3985_2 = {pp111[38]};
    Full_Adder FA_3985(s3985, c3985, in3985_1, in3985_2, pp109[40]);
    wire[0:0] s3986, in3986_1, in3986_2;
    wire c3986;
    assign in3986_1 = {pp113[36]};
    assign in3986_2 = {pp114[35]};
    Full_Adder FA_3986(s3986, c3986, in3986_1, in3986_2, pp112[37]);
    wire[0:0] s3987, in3987_1, in3987_2;
    wire c3987;
    assign in3987_1 = {pp116[33]};
    assign in3987_2 = {pp117[32]};
    Full_Adder FA_3987(s3987, c3987, in3987_1, in3987_2, pp115[34]);
    wire[0:0] s3988, in3988_1, in3988_2;
    wire c3988;
    assign in3988_1 = {pp119[30]};
    assign in3988_2 = {pp120[29]};
    Full_Adder FA_3988(s3988, c3988, in3988_1, in3988_2, pp118[31]);
    wire[0:0] s3989, in3989_1, in3989_2;
    wire c3989;
    assign in3989_1 = {pp122[27]};
    assign in3989_2 = {pp123[26]};
    Full_Adder FA_3989(s3989, c3989, in3989_1, in3989_2, pp121[28]);
    wire[0:0] s3990, in3990_1, in3990_2;
    wire c3990;
    assign in3990_1 = {pp125[24]};
    assign in3990_2 = {pp126[23]};
    Full_Adder FA_3990(s3990, c3990, in3990_1, in3990_2, pp124[25]);
    wire[0:0] s3991, in3991_1, in3991_2;
    wire c3991;
    assign in3991_1 = {c1554};
    assign in3991_2 = {c1555};
    Full_Adder FA_3991(s3991, c3991, in3991_1, in3991_2, pp127[22]);
    wire[0:0] s3992, in3992_1, in3992_2;
    wire c3992;
    assign in3992_1 = {c1557};
    assign in3992_2 = {c1558};
    Full_Adder FA_3992(s3992, c3992, in3992_1, in3992_2, c1556);
    wire[0:0] s3993, in3993_1, in3993_2;
    wire c3993;
    assign in3993_1 = {c1560};
    assign in3993_2 = {c1561};
    Full_Adder FA_3993(s3993, c3993, in3993_1, in3993_2, c1559);
    wire[0:0] s3994, in3994_1, in3994_2;
    wire c3994;
    assign in3994_1 = {c1563};
    assign in3994_2 = {c1564};
    Full_Adder FA_3994(s3994, c3994, in3994_1, in3994_2, c1562);
    wire[0:0] s3995, in3995_1, in3995_2;
    wire c3995;
    assign in3995_1 = {c1566};
    assign in3995_2 = {c1567};
    Full_Adder FA_3995(s3995, c3995, in3995_1, in3995_2, c1565);
    wire[0:0] s3996, in3996_1, in3996_2;
    wire c3996;
    assign in3996_1 = {c1569};
    assign in3996_2 = {c1570};
    Full_Adder FA_3996(s3996, c3996, in3996_1, in3996_2, c1568);
    wire[0:0] s3997, in3997_1, in3997_2;
    wire c3997;
    assign in3997_1 = {c1572};
    assign in3997_2 = {c1573};
    Full_Adder FA_3997(s3997, c3997, in3997_1, in3997_2, c1571);
    wire[0:0] s3998, in3998_1, in3998_2;
    wire c3998;
    assign in3998_1 = {c1575};
    assign in3998_2 = {s1576[0]};
    Full_Adder FA_3998(s3998, c3998, in3998_1, in3998_2, c1574);
    wire[0:0] s3999, in3999_1, in3999_2;
    wire c3999;
    assign in3999_1 = {s1578[0]};
    assign in3999_2 = {s1579[0]};
    Full_Adder FA_3999(s3999, c3999, in3999_1, in3999_2, s1577[0]);
    wire[0:0] s4000, in4000_1, in4000_2;
    wire c4000;
    assign in4000_1 = {s1581[0]};
    assign in4000_2 = {s1582[0]};
    Full_Adder FA_4000(s4000, c4000, in4000_1, in4000_2, s1580[0]);
    wire[0:0] s4001, in4001_1, in4001_2;
    wire c4001;
    assign in4001_1 = {s1584[0]};
    assign in4001_2 = {s1585[0]};
    Full_Adder FA_4001(s4001, c4001, in4001_1, in4001_2, s1583[0]);
    wire[0:0] s4002, in4002_1, in4002_2;
    wire c4002;
    assign in4002_1 = {s1587[0]};
    assign in4002_2 = {s1588[0]};
    Full_Adder FA_4002(s4002, c4002, in4002_1, in4002_2, s1586[0]);
    wire[0:0] s4003, in4003_1, in4003_2;
    wire c4003;
    assign in4003_1 = {s1590[0]};
    assign in4003_2 = {s1591[0]};
    Full_Adder FA_4003(s4003, c4003, in4003_1, in4003_2, s1589[0]);
    wire[0:0] s4004, in4004_1, in4004_2;
    wire c4004;
    assign in4004_1 = {s1593[0]};
    assign in4004_2 = {s1594[0]};
    Full_Adder FA_4004(s4004, c4004, in4004_1, in4004_2, s1592[0]);
    wire[0:0] s4005, in4005_1, in4005_2;
    wire c4005;
    assign in4005_1 = {pp84[66]};
    assign in4005_2 = {pp85[65]};
    Full_Adder FA_4005(s4005, c4005, in4005_1, in4005_2, pp83[67]);
    wire[0:0] s4006, in4006_1, in4006_2;
    wire c4006;
    assign in4006_1 = {pp87[63]};
    assign in4006_2 = {pp88[62]};
    Full_Adder FA_4006(s4006, c4006, in4006_1, in4006_2, pp86[64]);
    wire[0:0] s4007, in4007_1, in4007_2;
    wire c4007;
    assign in4007_1 = {pp90[60]};
    assign in4007_2 = {pp91[59]};
    Full_Adder FA_4007(s4007, c4007, in4007_1, in4007_2, pp89[61]);
    wire[0:0] s4008, in4008_1, in4008_2;
    wire c4008;
    assign in4008_1 = {pp93[57]};
    assign in4008_2 = {pp94[56]};
    Full_Adder FA_4008(s4008, c4008, in4008_1, in4008_2, pp92[58]);
    wire[0:0] s4009, in4009_1, in4009_2;
    wire c4009;
    assign in4009_1 = {pp96[54]};
    assign in4009_2 = {pp97[53]};
    Full_Adder FA_4009(s4009, c4009, in4009_1, in4009_2, pp95[55]);
    wire[0:0] s4010, in4010_1, in4010_2;
    wire c4010;
    assign in4010_1 = {pp99[51]};
    assign in4010_2 = {pp100[50]};
    Full_Adder FA_4010(s4010, c4010, in4010_1, in4010_2, pp98[52]);
    wire[0:0] s4011, in4011_1, in4011_2;
    wire c4011;
    assign in4011_1 = {pp102[48]};
    assign in4011_2 = {pp103[47]};
    Full_Adder FA_4011(s4011, c4011, in4011_1, in4011_2, pp101[49]);
    wire[0:0] s4012, in4012_1, in4012_2;
    wire c4012;
    assign in4012_1 = {pp105[45]};
    assign in4012_2 = {pp106[44]};
    Full_Adder FA_4012(s4012, c4012, in4012_1, in4012_2, pp104[46]);
    wire[0:0] s4013, in4013_1, in4013_2;
    wire c4013;
    assign in4013_1 = {pp108[42]};
    assign in4013_2 = {pp109[41]};
    Full_Adder FA_4013(s4013, c4013, in4013_1, in4013_2, pp107[43]);
    wire[0:0] s4014, in4014_1, in4014_2;
    wire c4014;
    assign in4014_1 = {pp111[39]};
    assign in4014_2 = {pp112[38]};
    Full_Adder FA_4014(s4014, c4014, in4014_1, in4014_2, pp110[40]);
    wire[0:0] s4015, in4015_1, in4015_2;
    wire c4015;
    assign in4015_1 = {pp114[36]};
    assign in4015_2 = {pp115[35]};
    Full_Adder FA_4015(s4015, c4015, in4015_1, in4015_2, pp113[37]);
    wire[0:0] s4016, in4016_1, in4016_2;
    wire c4016;
    assign in4016_1 = {pp117[33]};
    assign in4016_2 = {pp118[32]};
    Full_Adder FA_4016(s4016, c4016, in4016_1, in4016_2, pp116[34]);
    wire[0:0] s4017, in4017_1, in4017_2;
    wire c4017;
    assign in4017_1 = {pp120[30]};
    assign in4017_2 = {pp121[29]};
    Full_Adder FA_4017(s4017, c4017, in4017_1, in4017_2, pp119[31]);
    wire[0:0] s4018, in4018_1, in4018_2;
    wire c4018;
    assign in4018_1 = {pp123[27]};
    assign in4018_2 = {pp124[26]};
    Full_Adder FA_4018(s4018, c4018, in4018_1, in4018_2, pp122[28]);
    wire[0:0] s4019, in4019_1, in4019_2;
    wire c4019;
    assign in4019_1 = {pp126[24]};
    assign in4019_2 = {pp127[23]};
    Full_Adder FA_4019(s4019, c4019, in4019_1, in4019_2, pp125[25]);
    wire[0:0] s4020, in4020_1, in4020_2;
    wire c4020;
    assign in4020_1 = {c1577};
    assign in4020_2 = {c1578};
    Full_Adder FA_4020(s4020, c4020, in4020_1, in4020_2, c1576);
    wire[0:0] s4021, in4021_1, in4021_2;
    wire c4021;
    assign in4021_1 = {c1580};
    assign in4021_2 = {c1581};
    Full_Adder FA_4021(s4021, c4021, in4021_1, in4021_2, c1579);
    wire[0:0] s4022, in4022_1, in4022_2;
    wire c4022;
    assign in4022_1 = {c1583};
    assign in4022_2 = {c1584};
    Full_Adder FA_4022(s4022, c4022, in4022_1, in4022_2, c1582);
    wire[0:0] s4023, in4023_1, in4023_2;
    wire c4023;
    assign in4023_1 = {c1586};
    assign in4023_2 = {c1587};
    Full_Adder FA_4023(s4023, c4023, in4023_1, in4023_2, c1585);
    wire[0:0] s4024, in4024_1, in4024_2;
    wire c4024;
    assign in4024_1 = {c1589};
    assign in4024_2 = {c1590};
    Full_Adder FA_4024(s4024, c4024, in4024_1, in4024_2, c1588);
    wire[0:0] s4025, in4025_1, in4025_2;
    wire c4025;
    assign in4025_1 = {c1592};
    assign in4025_2 = {c1593};
    Full_Adder FA_4025(s4025, c4025, in4025_1, in4025_2, c1591);
    wire[0:0] s4026, in4026_1, in4026_2;
    wire c4026;
    assign in4026_1 = {c1595};
    assign in4026_2 = {c1596};
    Full_Adder FA_4026(s4026, c4026, in4026_1, in4026_2, c1594);
    wire[0:0] s4027, in4027_1, in4027_2;
    wire c4027;
    assign in4027_1 = {s1598[0]};
    assign in4027_2 = {s1599[0]};
    Full_Adder FA_4027(s4027, c4027, in4027_1, in4027_2, s1597[0]);
    wire[0:0] s4028, in4028_1, in4028_2;
    wire c4028;
    assign in4028_1 = {s1601[0]};
    assign in4028_2 = {s1602[0]};
    Full_Adder FA_4028(s4028, c4028, in4028_1, in4028_2, s1600[0]);
    wire[0:0] s4029, in4029_1, in4029_2;
    wire c4029;
    assign in4029_1 = {s1604[0]};
    assign in4029_2 = {s1605[0]};
    Full_Adder FA_4029(s4029, c4029, in4029_1, in4029_2, s1603[0]);
    wire[0:0] s4030, in4030_1, in4030_2;
    wire c4030;
    assign in4030_1 = {s1607[0]};
    assign in4030_2 = {s1608[0]};
    Full_Adder FA_4030(s4030, c4030, in4030_1, in4030_2, s1606[0]);
    wire[0:0] s4031, in4031_1, in4031_2;
    wire c4031;
    assign in4031_1 = {s1610[0]};
    assign in4031_2 = {s1611[0]};
    Full_Adder FA_4031(s4031, c4031, in4031_1, in4031_2, s1609[0]);
    wire[0:0] s4032, in4032_1, in4032_2;
    wire c4032;
    assign in4032_1 = {s1613[0]};
    assign in4032_2 = {s1614[0]};
    Full_Adder FA_4032(s4032, c4032, in4032_1, in4032_2, s1612[0]);
    wire[0:0] s4033, in4033_1, in4033_2;
    wire c4033;
    assign in4033_1 = {pp82[69]};
    assign in4033_2 = {pp83[68]};
    Full_Adder FA_4033(s4033, c4033, in4033_1, in4033_2, pp81[70]);
    wire[0:0] s4034, in4034_1, in4034_2;
    wire c4034;
    assign in4034_1 = {pp85[66]};
    assign in4034_2 = {pp86[65]};
    Full_Adder FA_4034(s4034, c4034, in4034_1, in4034_2, pp84[67]);
    wire[0:0] s4035, in4035_1, in4035_2;
    wire c4035;
    assign in4035_1 = {pp88[63]};
    assign in4035_2 = {pp89[62]};
    Full_Adder FA_4035(s4035, c4035, in4035_1, in4035_2, pp87[64]);
    wire[0:0] s4036, in4036_1, in4036_2;
    wire c4036;
    assign in4036_1 = {pp91[60]};
    assign in4036_2 = {pp92[59]};
    Full_Adder FA_4036(s4036, c4036, in4036_1, in4036_2, pp90[61]);
    wire[0:0] s4037, in4037_1, in4037_2;
    wire c4037;
    assign in4037_1 = {pp94[57]};
    assign in4037_2 = {pp95[56]};
    Full_Adder FA_4037(s4037, c4037, in4037_1, in4037_2, pp93[58]);
    wire[0:0] s4038, in4038_1, in4038_2;
    wire c4038;
    assign in4038_1 = {pp97[54]};
    assign in4038_2 = {pp98[53]};
    Full_Adder FA_4038(s4038, c4038, in4038_1, in4038_2, pp96[55]);
    wire[0:0] s4039, in4039_1, in4039_2;
    wire c4039;
    assign in4039_1 = {pp100[51]};
    assign in4039_2 = {pp101[50]};
    Full_Adder FA_4039(s4039, c4039, in4039_1, in4039_2, pp99[52]);
    wire[0:0] s4040, in4040_1, in4040_2;
    wire c4040;
    assign in4040_1 = {pp103[48]};
    assign in4040_2 = {pp104[47]};
    Full_Adder FA_4040(s4040, c4040, in4040_1, in4040_2, pp102[49]);
    wire[0:0] s4041, in4041_1, in4041_2;
    wire c4041;
    assign in4041_1 = {pp106[45]};
    assign in4041_2 = {pp107[44]};
    Full_Adder FA_4041(s4041, c4041, in4041_1, in4041_2, pp105[46]);
    wire[0:0] s4042, in4042_1, in4042_2;
    wire c4042;
    assign in4042_1 = {pp109[42]};
    assign in4042_2 = {pp110[41]};
    Full_Adder FA_4042(s4042, c4042, in4042_1, in4042_2, pp108[43]);
    wire[0:0] s4043, in4043_1, in4043_2;
    wire c4043;
    assign in4043_1 = {pp112[39]};
    assign in4043_2 = {pp113[38]};
    Full_Adder FA_4043(s4043, c4043, in4043_1, in4043_2, pp111[40]);
    wire[0:0] s4044, in4044_1, in4044_2;
    wire c4044;
    assign in4044_1 = {pp115[36]};
    assign in4044_2 = {pp116[35]};
    Full_Adder FA_4044(s4044, c4044, in4044_1, in4044_2, pp114[37]);
    wire[0:0] s4045, in4045_1, in4045_2;
    wire c4045;
    assign in4045_1 = {pp118[33]};
    assign in4045_2 = {pp119[32]};
    Full_Adder FA_4045(s4045, c4045, in4045_1, in4045_2, pp117[34]);
    wire[0:0] s4046, in4046_1, in4046_2;
    wire c4046;
    assign in4046_1 = {pp121[30]};
    assign in4046_2 = {pp122[29]};
    Full_Adder FA_4046(s4046, c4046, in4046_1, in4046_2, pp120[31]);
    wire[0:0] s4047, in4047_1, in4047_2;
    wire c4047;
    assign in4047_1 = {pp124[27]};
    assign in4047_2 = {pp125[26]};
    Full_Adder FA_4047(s4047, c4047, in4047_1, in4047_2, pp123[28]);
    wire[0:0] s4048, in4048_1, in4048_2;
    wire c4048;
    assign in4048_1 = {pp127[24]};
    assign in4048_2 = {c1597};
    Full_Adder FA_4048(s4048, c4048, in4048_1, in4048_2, pp126[25]);
    wire[0:0] s4049, in4049_1, in4049_2;
    wire c4049;
    assign in4049_1 = {c1599};
    assign in4049_2 = {c1600};
    Full_Adder FA_4049(s4049, c4049, in4049_1, in4049_2, c1598);
    wire[0:0] s4050, in4050_1, in4050_2;
    wire c4050;
    assign in4050_1 = {c1602};
    assign in4050_2 = {c1603};
    Full_Adder FA_4050(s4050, c4050, in4050_1, in4050_2, c1601);
    wire[0:0] s4051, in4051_1, in4051_2;
    wire c4051;
    assign in4051_1 = {c1605};
    assign in4051_2 = {c1606};
    Full_Adder FA_4051(s4051, c4051, in4051_1, in4051_2, c1604);
    wire[0:0] s4052, in4052_1, in4052_2;
    wire c4052;
    assign in4052_1 = {c1608};
    assign in4052_2 = {c1609};
    Full_Adder FA_4052(s4052, c4052, in4052_1, in4052_2, c1607);
    wire[0:0] s4053, in4053_1, in4053_2;
    wire c4053;
    assign in4053_1 = {c1611};
    assign in4053_2 = {c1612};
    Full_Adder FA_4053(s4053, c4053, in4053_1, in4053_2, c1610);
    wire[0:0] s4054, in4054_1, in4054_2;
    wire c4054;
    assign in4054_1 = {c1614};
    assign in4054_2 = {c1615};
    Full_Adder FA_4054(s4054, c4054, in4054_1, in4054_2, c1613);
    wire[0:0] s4055, in4055_1, in4055_2;
    wire c4055;
    assign in4055_1 = {s1617[0]};
    assign in4055_2 = {s1618[0]};
    Full_Adder FA_4055(s4055, c4055, in4055_1, in4055_2, c1616);
    wire[0:0] s4056, in4056_1, in4056_2;
    wire c4056;
    assign in4056_1 = {s1620[0]};
    assign in4056_2 = {s1621[0]};
    Full_Adder FA_4056(s4056, c4056, in4056_1, in4056_2, s1619[0]);
    wire[0:0] s4057, in4057_1, in4057_2;
    wire c4057;
    assign in4057_1 = {s1623[0]};
    assign in4057_2 = {s1624[0]};
    Full_Adder FA_4057(s4057, c4057, in4057_1, in4057_2, s1622[0]);
    wire[0:0] s4058, in4058_1, in4058_2;
    wire c4058;
    assign in4058_1 = {s1626[0]};
    assign in4058_2 = {s1627[0]};
    Full_Adder FA_4058(s4058, c4058, in4058_1, in4058_2, s1625[0]);
    wire[0:0] s4059, in4059_1, in4059_2;
    wire c4059;
    assign in4059_1 = {s1629[0]};
    assign in4059_2 = {s1630[0]};
    Full_Adder FA_4059(s4059, c4059, in4059_1, in4059_2, s1628[0]);
    wire[0:0] s4060, in4060_1, in4060_2;
    wire c4060;
    assign in4060_1 = {s1632[0]};
    assign in4060_2 = {s1633[0]};
    Full_Adder FA_4060(s4060, c4060, in4060_1, in4060_2, s1631[0]);
    wire[0:0] s4061, in4061_1, in4061_2;
    wire c4061;
    assign in4061_1 = {pp80[72]};
    assign in4061_2 = {pp81[71]};
    Full_Adder FA_4061(s4061, c4061, in4061_1, in4061_2, pp79[73]);
    wire[0:0] s4062, in4062_1, in4062_2;
    wire c4062;
    assign in4062_1 = {pp83[69]};
    assign in4062_2 = {pp84[68]};
    Full_Adder FA_4062(s4062, c4062, in4062_1, in4062_2, pp82[70]);
    wire[0:0] s4063, in4063_1, in4063_2;
    wire c4063;
    assign in4063_1 = {pp86[66]};
    assign in4063_2 = {pp87[65]};
    Full_Adder FA_4063(s4063, c4063, in4063_1, in4063_2, pp85[67]);
    wire[0:0] s4064, in4064_1, in4064_2;
    wire c4064;
    assign in4064_1 = {pp89[63]};
    assign in4064_2 = {pp90[62]};
    Full_Adder FA_4064(s4064, c4064, in4064_1, in4064_2, pp88[64]);
    wire[0:0] s4065, in4065_1, in4065_2;
    wire c4065;
    assign in4065_1 = {pp92[60]};
    assign in4065_2 = {pp93[59]};
    Full_Adder FA_4065(s4065, c4065, in4065_1, in4065_2, pp91[61]);
    wire[0:0] s4066, in4066_1, in4066_2;
    wire c4066;
    assign in4066_1 = {pp95[57]};
    assign in4066_2 = {pp96[56]};
    Full_Adder FA_4066(s4066, c4066, in4066_1, in4066_2, pp94[58]);
    wire[0:0] s4067, in4067_1, in4067_2;
    wire c4067;
    assign in4067_1 = {pp98[54]};
    assign in4067_2 = {pp99[53]};
    Full_Adder FA_4067(s4067, c4067, in4067_1, in4067_2, pp97[55]);
    wire[0:0] s4068, in4068_1, in4068_2;
    wire c4068;
    assign in4068_1 = {pp101[51]};
    assign in4068_2 = {pp102[50]};
    Full_Adder FA_4068(s4068, c4068, in4068_1, in4068_2, pp100[52]);
    wire[0:0] s4069, in4069_1, in4069_2;
    wire c4069;
    assign in4069_1 = {pp104[48]};
    assign in4069_2 = {pp105[47]};
    Full_Adder FA_4069(s4069, c4069, in4069_1, in4069_2, pp103[49]);
    wire[0:0] s4070, in4070_1, in4070_2;
    wire c4070;
    assign in4070_1 = {pp107[45]};
    assign in4070_2 = {pp108[44]};
    Full_Adder FA_4070(s4070, c4070, in4070_1, in4070_2, pp106[46]);
    wire[0:0] s4071, in4071_1, in4071_2;
    wire c4071;
    assign in4071_1 = {pp110[42]};
    assign in4071_2 = {pp111[41]};
    Full_Adder FA_4071(s4071, c4071, in4071_1, in4071_2, pp109[43]);
    wire[0:0] s4072, in4072_1, in4072_2;
    wire c4072;
    assign in4072_1 = {pp113[39]};
    assign in4072_2 = {pp114[38]};
    Full_Adder FA_4072(s4072, c4072, in4072_1, in4072_2, pp112[40]);
    wire[0:0] s4073, in4073_1, in4073_2;
    wire c4073;
    assign in4073_1 = {pp116[36]};
    assign in4073_2 = {pp117[35]};
    Full_Adder FA_4073(s4073, c4073, in4073_1, in4073_2, pp115[37]);
    wire[0:0] s4074, in4074_1, in4074_2;
    wire c4074;
    assign in4074_1 = {pp119[33]};
    assign in4074_2 = {pp120[32]};
    Full_Adder FA_4074(s4074, c4074, in4074_1, in4074_2, pp118[34]);
    wire[0:0] s4075, in4075_1, in4075_2;
    wire c4075;
    assign in4075_1 = {pp122[30]};
    assign in4075_2 = {pp123[29]};
    Full_Adder FA_4075(s4075, c4075, in4075_1, in4075_2, pp121[31]);
    wire[0:0] s4076, in4076_1, in4076_2;
    wire c4076;
    assign in4076_1 = {pp125[27]};
    assign in4076_2 = {pp126[26]};
    Full_Adder FA_4076(s4076, c4076, in4076_1, in4076_2, pp124[28]);
    wire[0:0] s4077, in4077_1, in4077_2;
    wire c4077;
    assign in4077_1 = {c1617};
    assign in4077_2 = {c1618};
    Full_Adder FA_4077(s4077, c4077, in4077_1, in4077_2, pp127[25]);
    wire[0:0] s4078, in4078_1, in4078_2;
    wire c4078;
    assign in4078_1 = {c1620};
    assign in4078_2 = {c1621};
    Full_Adder FA_4078(s4078, c4078, in4078_1, in4078_2, c1619);
    wire[0:0] s4079, in4079_1, in4079_2;
    wire c4079;
    assign in4079_1 = {c1623};
    assign in4079_2 = {c1624};
    Full_Adder FA_4079(s4079, c4079, in4079_1, in4079_2, c1622);
    wire[0:0] s4080, in4080_1, in4080_2;
    wire c4080;
    assign in4080_1 = {c1626};
    assign in4080_2 = {c1627};
    Full_Adder FA_4080(s4080, c4080, in4080_1, in4080_2, c1625);
    wire[0:0] s4081, in4081_1, in4081_2;
    wire c4081;
    assign in4081_1 = {c1629};
    assign in4081_2 = {c1630};
    Full_Adder FA_4081(s4081, c4081, in4081_1, in4081_2, c1628);
    wire[0:0] s4082, in4082_1, in4082_2;
    wire c4082;
    assign in4082_1 = {c1632};
    assign in4082_2 = {c1633};
    Full_Adder FA_4082(s4082, c4082, in4082_1, in4082_2, c1631);
    wire[0:0] s4083, in4083_1, in4083_2;
    wire c4083;
    assign in4083_1 = {c1635};
    assign in4083_2 = {s1636[0]};
    Full_Adder FA_4083(s4083, c4083, in4083_1, in4083_2, c1634);
    wire[0:0] s4084, in4084_1, in4084_2;
    wire c4084;
    assign in4084_1 = {s1638[0]};
    assign in4084_2 = {s1639[0]};
    Full_Adder FA_4084(s4084, c4084, in4084_1, in4084_2, s1637[0]);
    wire[0:0] s4085, in4085_1, in4085_2;
    wire c4085;
    assign in4085_1 = {s1641[0]};
    assign in4085_2 = {s1642[0]};
    Full_Adder FA_4085(s4085, c4085, in4085_1, in4085_2, s1640[0]);
    wire[0:0] s4086, in4086_1, in4086_2;
    wire c4086;
    assign in4086_1 = {s1644[0]};
    assign in4086_2 = {s1645[0]};
    Full_Adder FA_4086(s4086, c4086, in4086_1, in4086_2, s1643[0]);
    wire[0:0] s4087, in4087_1, in4087_2;
    wire c4087;
    assign in4087_1 = {s1647[0]};
    assign in4087_2 = {s1648[0]};
    Full_Adder FA_4087(s4087, c4087, in4087_1, in4087_2, s1646[0]);
    wire[0:0] s4088, in4088_1, in4088_2;
    wire c4088;
    assign in4088_1 = {s1650[0]};
    assign in4088_2 = {s1651[0]};
    Full_Adder FA_4088(s4088, c4088, in4088_1, in4088_2, s1649[0]);
    wire[0:0] s4089, in4089_1, in4089_2;
    wire c4089;
    assign in4089_1 = {pp78[75]};
    assign in4089_2 = {pp79[74]};
    Full_Adder FA_4089(s4089, c4089, in4089_1, in4089_2, pp77[76]);
    wire[0:0] s4090, in4090_1, in4090_2;
    wire c4090;
    assign in4090_1 = {pp81[72]};
    assign in4090_2 = {pp82[71]};
    Full_Adder FA_4090(s4090, c4090, in4090_1, in4090_2, pp80[73]);
    wire[0:0] s4091, in4091_1, in4091_2;
    wire c4091;
    assign in4091_1 = {pp84[69]};
    assign in4091_2 = {pp85[68]};
    Full_Adder FA_4091(s4091, c4091, in4091_1, in4091_2, pp83[70]);
    wire[0:0] s4092, in4092_1, in4092_2;
    wire c4092;
    assign in4092_1 = {pp87[66]};
    assign in4092_2 = {pp88[65]};
    Full_Adder FA_4092(s4092, c4092, in4092_1, in4092_2, pp86[67]);
    wire[0:0] s4093, in4093_1, in4093_2;
    wire c4093;
    assign in4093_1 = {pp90[63]};
    assign in4093_2 = {pp91[62]};
    Full_Adder FA_4093(s4093, c4093, in4093_1, in4093_2, pp89[64]);
    wire[0:0] s4094, in4094_1, in4094_2;
    wire c4094;
    assign in4094_1 = {pp93[60]};
    assign in4094_2 = {pp94[59]};
    Full_Adder FA_4094(s4094, c4094, in4094_1, in4094_2, pp92[61]);
    wire[0:0] s4095, in4095_1, in4095_2;
    wire c4095;
    assign in4095_1 = {pp96[57]};
    assign in4095_2 = {pp97[56]};
    Full_Adder FA_4095(s4095, c4095, in4095_1, in4095_2, pp95[58]);
    wire[0:0] s4096, in4096_1, in4096_2;
    wire c4096;
    assign in4096_1 = {pp99[54]};
    assign in4096_2 = {pp100[53]};
    Full_Adder FA_4096(s4096, c4096, in4096_1, in4096_2, pp98[55]);
    wire[0:0] s4097, in4097_1, in4097_2;
    wire c4097;
    assign in4097_1 = {pp102[51]};
    assign in4097_2 = {pp103[50]};
    Full_Adder FA_4097(s4097, c4097, in4097_1, in4097_2, pp101[52]);
    wire[0:0] s4098, in4098_1, in4098_2;
    wire c4098;
    assign in4098_1 = {pp105[48]};
    assign in4098_2 = {pp106[47]};
    Full_Adder FA_4098(s4098, c4098, in4098_1, in4098_2, pp104[49]);
    wire[0:0] s4099, in4099_1, in4099_2;
    wire c4099;
    assign in4099_1 = {pp108[45]};
    assign in4099_2 = {pp109[44]};
    Full_Adder FA_4099(s4099, c4099, in4099_1, in4099_2, pp107[46]);
    wire[0:0] s4100, in4100_1, in4100_2;
    wire c4100;
    assign in4100_1 = {pp111[42]};
    assign in4100_2 = {pp112[41]};
    Full_Adder FA_4100(s4100, c4100, in4100_1, in4100_2, pp110[43]);
    wire[0:0] s4101, in4101_1, in4101_2;
    wire c4101;
    assign in4101_1 = {pp114[39]};
    assign in4101_2 = {pp115[38]};
    Full_Adder FA_4101(s4101, c4101, in4101_1, in4101_2, pp113[40]);
    wire[0:0] s4102, in4102_1, in4102_2;
    wire c4102;
    assign in4102_1 = {pp117[36]};
    assign in4102_2 = {pp118[35]};
    Full_Adder FA_4102(s4102, c4102, in4102_1, in4102_2, pp116[37]);
    wire[0:0] s4103, in4103_1, in4103_2;
    wire c4103;
    assign in4103_1 = {pp120[33]};
    assign in4103_2 = {pp121[32]};
    Full_Adder FA_4103(s4103, c4103, in4103_1, in4103_2, pp119[34]);
    wire[0:0] s4104, in4104_1, in4104_2;
    wire c4104;
    assign in4104_1 = {pp123[30]};
    assign in4104_2 = {pp124[29]};
    Full_Adder FA_4104(s4104, c4104, in4104_1, in4104_2, pp122[31]);
    wire[0:0] s4105, in4105_1, in4105_2;
    wire c4105;
    assign in4105_1 = {pp126[27]};
    assign in4105_2 = {pp127[26]};
    Full_Adder FA_4105(s4105, c4105, in4105_1, in4105_2, pp125[28]);
    wire[0:0] s4106, in4106_1, in4106_2;
    wire c4106;
    assign in4106_1 = {c1637};
    assign in4106_2 = {c1638};
    Full_Adder FA_4106(s4106, c4106, in4106_1, in4106_2, c1636);
    wire[0:0] s4107, in4107_1, in4107_2;
    wire c4107;
    assign in4107_1 = {c1640};
    assign in4107_2 = {c1641};
    Full_Adder FA_4107(s4107, c4107, in4107_1, in4107_2, c1639);
    wire[0:0] s4108, in4108_1, in4108_2;
    wire c4108;
    assign in4108_1 = {c1643};
    assign in4108_2 = {c1644};
    Full_Adder FA_4108(s4108, c4108, in4108_1, in4108_2, c1642);
    wire[0:0] s4109, in4109_1, in4109_2;
    wire c4109;
    assign in4109_1 = {c1646};
    assign in4109_2 = {c1647};
    Full_Adder FA_4109(s4109, c4109, in4109_1, in4109_2, c1645);
    wire[0:0] s4110, in4110_1, in4110_2;
    wire c4110;
    assign in4110_1 = {c1649};
    assign in4110_2 = {c1650};
    Full_Adder FA_4110(s4110, c4110, in4110_1, in4110_2, c1648);
    wire[0:0] s4111, in4111_1, in4111_2;
    wire c4111;
    assign in4111_1 = {c1652};
    assign in4111_2 = {c1653};
    Full_Adder FA_4111(s4111, c4111, in4111_1, in4111_2, c1651);
    wire[0:0] s4112, in4112_1, in4112_2;
    wire c4112;
    assign in4112_1 = {s1655[0]};
    assign in4112_2 = {s1656[0]};
    Full_Adder FA_4112(s4112, c4112, in4112_1, in4112_2, s1654[0]);
    wire[0:0] s4113, in4113_1, in4113_2;
    wire c4113;
    assign in4113_1 = {s1658[0]};
    assign in4113_2 = {s1659[0]};
    Full_Adder FA_4113(s4113, c4113, in4113_1, in4113_2, s1657[0]);
    wire[0:0] s4114, in4114_1, in4114_2;
    wire c4114;
    assign in4114_1 = {s1661[0]};
    assign in4114_2 = {s1662[0]};
    Full_Adder FA_4114(s4114, c4114, in4114_1, in4114_2, s1660[0]);
    wire[0:0] s4115, in4115_1, in4115_2;
    wire c4115;
    assign in4115_1 = {s1664[0]};
    assign in4115_2 = {s1665[0]};
    Full_Adder FA_4115(s4115, c4115, in4115_1, in4115_2, s1663[0]);
    wire[0:0] s4116, in4116_1, in4116_2;
    wire c4116;
    assign in4116_1 = {s1667[0]};
    assign in4116_2 = {s1668[0]};
    Full_Adder FA_4116(s4116, c4116, in4116_1, in4116_2, s1666[0]);
    wire[0:0] s4117, in4117_1, in4117_2;
    wire c4117;
    assign in4117_1 = {pp76[78]};
    assign in4117_2 = {pp77[77]};
    Full_Adder FA_4117(s4117, c4117, in4117_1, in4117_2, pp75[79]);
    wire[0:0] s4118, in4118_1, in4118_2;
    wire c4118;
    assign in4118_1 = {pp79[75]};
    assign in4118_2 = {pp80[74]};
    Full_Adder FA_4118(s4118, c4118, in4118_1, in4118_2, pp78[76]);
    wire[0:0] s4119, in4119_1, in4119_2;
    wire c4119;
    assign in4119_1 = {pp82[72]};
    assign in4119_2 = {pp83[71]};
    Full_Adder FA_4119(s4119, c4119, in4119_1, in4119_2, pp81[73]);
    wire[0:0] s4120, in4120_1, in4120_2;
    wire c4120;
    assign in4120_1 = {pp85[69]};
    assign in4120_2 = {pp86[68]};
    Full_Adder FA_4120(s4120, c4120, in4120_1, in4120_2, pp84[70]);
    wire[0:0] s4121, in4121_1, in4121_2;
    wire c4121;
    assign in4121_1 = {pp88[66]};
    assign in4121_2 = {pp89[65]};
    Full_Adder FA_4121(s4121, c4121, in4121_1, in4121_2, pp87[67]);
    wire[0:0] s4122, in4122_1, in4122_2;
    wire c4122;
    assign in4122_1 = {pp91[63]};
    assign in4122_2 = {pp92[62]};
    Full_Adder FA_4122(s4122, c4122, in4122_1, in4122_2, pp90[64]);
    wire[0:0] s4123, in4123_1, in4123_2;
    wire c4123;
    assign in4123_1 = {pp94[60]};
    assign in4123_2 = {pp95[59]};
    Full_Adder FA_4123(s4123, c4123, in4123_1, in4123_2, pp93[61]);
    wire[0:0] s4124, in4124_1, in4124_2;
    wire c4124;
    assign in4124_1 = {pp97[57]};
    assign in4124_2 = {pp98[56]};
    Full_Adder FA_4124(s4124, c4124, in4124_1, in4124_2, pp96[58]);
    wire[0:0] s4125, in4125_1, in4125_2;
    wire c4125;
    assign in4125_1 = {pp100[54]};
    assign in4125_2 = {pp101[53]};
    Full_Adder FA_4125(s4125, c4125, in4125_1, in4125_2, pp99[55]);
    wire[0:0] s4126, in4126_1, in4126_2;
    wire c4126;
    assign in4126_1 = {pp103[51]};
    assign in4126_2 = {pp104[50]};
    Full_Adder FA_4126(s4126, c4126, in4126_1, in4126_2, pp102[52]);
    wire[0:0] s4127, in4127_1, in4127_2;
    wire c4127;
    assign in4127_1 = {pp106[48]};
    assign in4127_2 = {pp107[47]};
    Full_Adder FA_4127(s4127, c4127, in4127_1, in4127_2, pp105[49]);
    wire[0:0] s4128, in4128_1, in4128_2;
    wire c4128;
    assign in4128_1 = {pp109[45]};
    assign in4128_2 = {pp110[44]};
    Full_Adder FA_4128(s4128, c4128, in4128_1, in4128_2, pp108[46]);
    wire[0:0] s4129, in4129_1, in4129_2;
    wire c4129;
    assign in4129_1 = {pp112[42]};
    assign in4129_2 = {pp113[41]};
    Full_Adder FA_4129(s4129, c4129, in4129_1, in4129_2, pp111[43]);
    wire[0:0] s4130, in4130_1, in4130_2;
    wire c4130;
    assign in4130_1 = {pp115[39]};
    assign in4130_2 = {pp116[38]};
    Full_Adder FA_4130(s4130, c4130, in4130_1, in4130_2, pp114[40]);
    wire[0:0] s4131, in4131_1, in4131_2;
    wire c4131;
    assign in4131_1 = {pp118[36]};
    assign in4131_2 = {pp119[35]};
    Full_Adder FA_4131(s4131, c4131, in4131_1, in4131_2, pp117[37]);
    wire[0:0] s4132, in4132_1, in4132_2;
    wire c4132;
    assign in4132_1 = {pp121[33]};
    assign in4132_2 = {pp122[32]};
    Full_Adder FA_4132(s4132, c4132, in4132_1, in4132_2, pp120[34]);
    wire[0:0] s4133, in4133_1, in4133_2;
    wire c4133;
    assign in4133_1 = {pp124[30]};
    assign in4133_2 = {pp125[29]};
    Full_Adder FA_4133(s4133, c4133, in4133_1, in4133_2, pp123[31]);
    wire[0:0] s4134, in4134_1, in4134_2;
    wire c4134;
    assign in4134_1 = {pp127[27]};
    assign in4134_2 = {c1654};
    Full_Adder FA_4134(s4134, c4134, in4134_1, in4134_2, pp126[28]);
    wire[0:0] s4135, in4135_1, in4135_2;
    wire c4135;
    assign in4135_1 = {c1656};
    assign in4135_2 = {c1657};
    Full_Adder FA_4135(s4135, c4135, in4135_1, in4135_2, c1655);
    wire[0:0] s4136, in4136_1, in4136_2;
    wire c4136;
    assign in4136_1 = {c1659};
    assign in4136_2 = {c1660};
    Full_Adder FA_4136(s4136, c4136, in4136_1, in4136_2, c1658);
    wire[0:0] s4137, in4137_1, in4137_2;
    wire c4137;
    assign in4137_1 = {c1662};
    assign in4137_2 = {c1663};
    Full_Adder FA_4137(s4137, c4137, in4137_1, in4137_2, c1661);
    wire[0:0] s4138, in4138_1, in4138_2;
    wire c4138;
    assign in4138_1 = {c1665};
    assign in4138_2 = {c1666};
    Full_Adder FA_4138(s4138, c4138, in4138_1, in4138_2, c1664);
    wire[0:0] s4139, in4139_1, in4139_2;
    wire c4139;
    assign in4139_1 = {c1668};
    assign in4139_2 = {c1669};
    Full_Adder FA_4139(s4139, c4139, in4139_1, in4139_2, c1667);
    wire[0:0] s4140, in4140_1, in4140_2;
    wire c4140;
    assign in4140_1 = {s1671[0]};
    assign in4140_2 = {s1672[0]};
    Full_Adder FA_4140(s4140, c4140, in4140_1, in4140_2, c1670);
    wire[0:0] s4141, in4141_1, in4141_2;
    wire c4141;
    assign in4141_1 = {s1674[0]};
    assign in4141_2 = {s1675[0]};
    Full_Adder FA_4141(s4141, c4141, in4141_1, in4141_2, s1673[0]);
    wire[0:0] s4142, in4142_1, in4142_2;
    wire c4142;
    assign in4142_1 = {s1677[0]};
    assign in4142_2 = {s1678[0]};
    Full_Adder FA_4142(s4142, c4142, in4142_1, in4142_2, s1676[0]);
    wire[0:0] s4143, in4143_1, in4143_2;
    wire c4143;
    assign in4143_1 = {s1680[0]};
    assign in4143_2 = {s1681[0]};
    Full_Adder FA_4143(s4143, c4143, in4143_1, in4143_2, s1679[0]);
    wire[0:0] s4144, in4144_1, in4144_2;
    wire c4144;
    assign in4144_1 = {s1683[0]};
    assign in4144_2 = {s1684[0]};
    Full_Adder FA_4144(s4144, c4144, in4144_1, in4144_2, s1682[0]);
    wire[0:0] s4145, in4145_1, in4145_2;
    wire c4145;
    assign in4145_1 = {pp74[81]};
    assign in4145_2 = {pp75[80]};
    Full_Adder FA_4145(s4145, c4145, in4145_1, in4145_2, pp73[82]);
    wire[0:0] s4146, in4146_1, in4146_2;
    wire c4146;
    assign in4146_1 = {pp77[78]};
    assign in4146_2 = {pp78[77]};
    Full_Adder FA_4146(s4146, c4146, in4146_1, in4146_2, pp76[79]);
    wire[0:0] s4147, in4147_1, in4147_2;
    wire c4147;
    assign in4147_1 = {pp80[75]};
    assign in4147_2 = {pp81[74]};
    Full_Adder FA_4147(s4147, c4147, in4147_1, in4147_2, pp79[76]);
    wire[0:0] s4148, in4148_1, in4148_2;
    wire c4148;
    assign in4148_1 = {pp83[72]};
    assign in4148_2 = {pp84[71]};
    Full_Adder FA_4148(s4148, c4148, in4148_1, in4148_2, pp82[73]);
    wire[0:0] s4149, in4149_1, in4149_2;
    wire c4149;
    assign in4149_1 = {pp86[69]};
    assign in4149_2 = {pp87[68]};
    Full_Adder FA_4149(s4149, c4149, in4149_1, in4149_2, pp85[70]);
    wire[0:0] s4150, in4150_1, in4150_2;
    wire c4150;
    assign in4150_1 = {pp89[66]};
    assign in4150_2 = {pp90[65]};
    Full_Adder FA_4150(s4150, c4150, in4150_1, in4150_2, pp88[67]);
    wire[0:0] s4151, in4151_1, in4151_2;
    wire c4151;
    assign in4151_1 = {pp92[63]};
    assign in4151_2 = {pp93[62]};
    Full_Adder FA_4151(s4151, c4151, in4151_1, in4151_2, pp91[64]);
    wire[0:0] s4152, in4152_1, in4152_2;
    wire c4152;
    assign in4152_1 = {pp95[60]};
    assign in4152_2 = {pp96[59]};
    Full_Adder FA_4152(s4152, c4152, in4152_1, in4152_2, pp94[61]);
    wire[0:0] s4153, in4153_1, in4153_2;
    wire c4153;
    assign in4153_1 = {pp98[57]};
    assign in4153_2 = {pp99[56]};
    Full_Adder FA_4153(s4153, c4153, in4153_1, in4153_2, pp97[58]);
    wire[0:0] s4154, in4154_1, in4154_2;
    wire c4154;
    assign in4154_1 = {pp101[54]};
    assign in4154_2 = {pp102[53]};
    Full_Adder FA_4154(s4154, c4154, in4154_1, in4154_2, pp100[55]);
    wire[0:0] s4155, in4155_1, in4155_2;
    wire c4155;
    assign in4155_1 = {pp104[51]};
    assign in4155_2 = {pp105[50]};
    Full_Adder FA_4155(s4155, c4155, in4155_1, in4155_2, pp103[52]);
    wire[0:0] s4156, in4156_1, in4156_2;
    wire c4156;
    assign in4156_1 = {pp107[48]};
    assign in4156_2 = {pp108[47]};
    Full_Adder FA_4156(s4156, c4156, in4156_1, in4156_2, pp106[49]);
    wire[0:0] s4157, in4157_1, in4157_2;
    wire c4157;
    assign in4157_1 = {pp110[45]};
    assign in4157_2 = {pp111[44]};
    Full_Adder FA_4157(s4157, c4157, in4157_1, in4157_2, pp109[46]);
    wire[0:0] s4158, in4158_1, in4158_2;
    wire c4158;
    assign in4158_1 = {pp113[42]};
    assign in4158_2 = {pp114[41]};
    Full_Adder FA_4158(s4158, c4158, in4158_1, in4158_2, pp112[43]);
    wire[0:0] s4159, in4159_1, in4159_2;
    wire c4159;
    assign in4159_1 = {pp116[39]};
    assign in4159_2 = {pp117[38]};
    Full_Adder FA_4159(s4159, c4159, in4159_1, in4159_2, pp115[40]);
    wire[0:0] s4160, in4160_1, in4160_2;
    wire c4160;
    assign in4160_1 = {pp119[36]};
    assign in4160_2 = {pp120[35]};
    Full_Adder FA_4160(s4160, c4160, in4160_1, in4160_2, pp118[37]);
    wire[0:0] s4161, in4161_1, in4161_2;
    wire c4161;
    assign in4161_1 = {pp122[33]};
    assign in4161_2 = {pp123[32]};
    Full_Adder FA_4161(s4161, c4161, in4161_1, in4161_2, pp121[34]);
    wire[0:0] s4162, in4162_1, in4162_2;
    wire c4162;
    assign in4162_1 = {pp125[30]};
    assign in4162_2 = {pp126[29]};
    Full_Adder FA_4162(s4162, c4162, in4162_1, in4162_2, pp124[31]);
    wire[0:0] s4163, in4163_1, in4163_2;
    wire c4163;
    assign in4163_1 = {c1671};
    assign in4163_2 = {c1672};
    Full_Adder FA_4163(s4163, c4163, in4163_1, in4163_2, pp127[28]);
    wire[0:0] s4164, in4164_1, in4164_2;
    wire c4164;
    assign in4164_1 = {c1674};
    assign in4164_2 = {c1675};
    Full_Adder FA_4164(s4164, c4164, in4164_1, in4164_2, c1673);
    wire[0:0] s4165, in4165_1, in4165_2;
    wire c4165;
    assign in4165_1 = {c1677};
    assign in4165_2 = {c1678};
    Full_Adder FA_4165(s4165, c4165, in4165_1, in4165_2, c1676);
    wire[0:0] s4166, in4166_1, in4166_2;
    wire c4166;
    assign in4166_1 = {c1680};
    assign in4166_2 = {c1681};
    Full_Adder FA_4166(s4166, c4166, in4166_1, in4166_2, c1679);
    wire[0:0] s4167, in4167_1, in4167_2;
    wire c4167;
    assign in4167_1 = {c1683};
    assign in4167_2 = {c1684};
    Full_Adder FA_4167(s4167, c4167, in4167_1, in4167_2, c1682);
    wire[0:0] s4168, in4168_1, in4168_2;
    wire c4168;
    assign in4168_1 = {c1686};
    assign in4168_2 = {s1687[0]};
    Full_Adder FA_4168(s4168, c4168, in4168_1, in4168_2, c1685);
    wire[0:0] s4169, in4169_1, in4169_2;
    wire c4169;
    assign in4169_1 = {s1689[0]};
    assign in4169_2 = {s1690[0]};
    Full_Adder FA_4169(s4169, c4169, in4169_1, in4169_2, s1688[0]);
    wire[0:0] s4170, in4170_1, in4170_2;
    wire c4170;
    assign in4170_1 = {s1692[0]};
    assign in4170_2 = {s1693[0]};
    Full_Adder FA_4170(s4170, c4170, in4170_1, in4170_2, s1691[0]);
    wire[0:0] s4171, in4171_1, in4171_2;
    wire c4171;
    assign in4171_1 = {s1695[0]};
    assign in4171_2 = {s1696[0]};
    Full_Adder FA_4171(s4171, c4171, in4171_1, in4171_2, s1694[0]);
    wire[0:0] s4172, in4172_1, in4172_2;
    wire c4172;
    assign in4172_1 = {s1698[0]};
    assign in4172_2 = {s1699[0]};
    Full_Adder FA_4172(s4172, c4172, in4172_1, in4172_2, s1697[0]);
    wire[0:0] s4173, in4173_1, in4173_2;
    wire c4173;
    assign in4173_1 = {pp72[84]};
    assign in4173_2 = {pp73[83]};
    Full_Adder FA_4173(s4173, c4173, in4173_1, in4173_2, pp71[85]);
    wire[0:0] s4174, in4174_1, in4174_2;
    wire c4174;
    assign in4174_1 = {pp75[81]};
    assign in4174_2 = {pp76[80]};
    Full_Adder FA_4174(s4174, c4174, in4174_1, in4174_2, pp74[82]);
    wire[0:0] s4175, in4175_1, in4175_2;
    wire c4175;
    assign in4175_1 = {pp78[78]};
    assign in4175_2 = {pp79[77]};
    Full_Adder FA_4175(s4175, c4175, in4175_1, in4175_2, pp77[79]);
    wire[0:0] s4176, in4176_1, in4176_2;
    wire c4176;
    assign in4176_1 = {pp81[75]};
    assign in4176_2 = {pp82[74]};
    Full_Adder FA_4176(s4176, c4176, in4176_1, in4176_2, pp80[76]);
    wire[0:0] s4177, in4177_1, in4177_2;
    wire c4177;
    assign in4177_1 = {pp84[72]};
    assign in4177_2 = {pp85[71]};
    Full_Adder FA_4177(s4177, c4177, in4177_1, in4177_2, pp83[73]);
    wire[0:0] s4178, in4178_1, in4178_2;
    wire c4178;
    assign in4178_1 = {pp87[69]};
    assign in4178_2 = {pp88[68]};
    Full_Adder FA_4178(s4178, c4178, in4178_1, in4178_2, pp86[70]);
    wire[0:0] s4179, in4179_1, in4179_2;
    wire c4179;
    assign in4179_1 = {pp90[66]};
    assign in4179_2 = {pp91[65]};
    Full_Adder FA_4179(s4179, c4179, in4179_1, in4179_2, pp89[67]);
    wire[0:0] s4180, in4180_1, in4180_2;
    wire c4180;
    assign in4180_1 = {pp93[63]};
    assign in4180_2 = {pp94[62]};
    Full_Adder FA_4180(s4180, c4180, in4180_1, in4180_2, pp92[64]);
    wire[0:0] s4181, in4181_1, in4181_2;
    wire c4181;
    assign in4181_1 = {pp96[60]};
    assign in4181_2 = {pp97[59]};
    Full_Adder FA_4181(s4181, c4181, in4181_1, in4181_2, pp95[61]);
    wire[0:0] s4182, in4182_1, in4182_2;
    wire c4182;
    assign in4182_1 = {pp99[57]};
    assign in4182_2 = {pp100[56]};
    Full_Adder FA_4182(s4182, c4182, in4182_1, in4182_2, pp98[58]);
    wire[0:0] s4183, in4183_1, in4183_2;
    wire c4183;
    assign in4183_1 = {pp102[54]};
    assign in4183_2 = {pp103[53]};
    Full_Adder FA_4183(s4183, c4183, in4183_1, in4183_2, pp101[55]);
    wire[0:0] s4184, in4184_1, in4184_2;
    wire c4184;
    assign in4184_1 = {pp105[51]};
    assign in4184_2 = {pp106[50]};
    Full_Adder FA_4184(s4184, c4184, in4184_1, in4184_2, pp104[52]);
    wire[0:0] s4185, in4185_1, in4185_2;
    wire c4185;
    assign in4185_1 = {pp108[48]};
    assign in4185_2 = {pp109[47]};
    Full_Adder FA_4185(s4185, c4185, in4185_1, in4185_2, pp107[49]);
    wire[0:0] s4186, in4186_1, in4186_2;
    wire c4186;
    assign in4186_1 = {pp111[45]};
    assign in4186_2 = {pp112[44]};
    Full_Adder FA_4186(s4186, c4186, in4186_1, in4186_2, pp110[46]);
    wire[0:0] s4187, in4187_1, in4187_2;
    wire c4187;
    assign in4187_1 = {pp114[42]};
    assign in4187_2 = {pp115[41]};
    Full_Adder FA_4187(s4187, c4187, in4187_1, in4187_2, pp113[43]);
    wire[0:0] s4188, in4188_1, in4188_2;
    wire c4188;
    assign in4188_1 = {pp117[39]};
    assign in4188_2 = {pp118[38]};
    Full_Adder FA_4188(s4188, c4188, in4188_1, in4188_2, pp116[40]);
    wire[0:0] s4189, in4189_1, in4189_2;
    wire c4189;
    assign in4189_1 = {pp120[36]};
    assign in4189_2 = {pp121[35]};
    Full_Adder FA_4189(s4189, c4189, in4189_1, in4189_2, pp119[37]);
    wire[0:0] s4190, in4190_1, in4190_2;
    wire c4190;
    assign in4190_1 = {pp123[33]};
    assign in4190_2 = {pp124[32]};
    Full_Adder FA_4190(s4190, c4190, in4190_1, in4190_2, pp122[34]);
    wire[0:0] s4191, in4191_1, in4191_2;
    wire c4191;
    assign in4191_1 = {pp126[30]};
    assign in4191_2 = {pp127[29]};
    Full_Adder FA_4191(s4191, c4191, in4191_1, in4191_2, pp125[31]);
    wire[0:0] s4192, in4192_1, in4192_2;
    wire c4192;
    assign in4192_1 = {c1688};
    assign in4192_2 = {c1689};
    Full_Adder FA_4192(s4192, c4192, in4192_1, in4192_2, c1687);
    wire[0:0] s4193, in4193_1, in4193_2;
    wire c4193;
    assign in4193_1 = {c1691};
    assign in4193_2 = {c1692};
    Full_Adder FA_4193(s4193, c4193, in4193_1, in4193_2, c1690);
    wire[0:0] s4194, in4194_1, in4194_2;
    wire c4194;
    assign in4194_1 = {c1694};
    assign in4194_2 = {c1695};
    Full_Adder FA_4194(s4194, c4194, in4194_1, in4194_2, c1693);
    wire[0:0] s4195, in4195_1, in4195_2;
    wire c4195;
    assign in4195_1 = {c1697};
    assign in4195_2 = {c1698};
    Full_Adder FA_4195(s4195, c4195, in4195_1, in4195_2, c1696);
    wire[0:0] s4196, in4196_1, in4196_2;
    wire c4196;
    assign in4196_1 = {c1700};
    assign in4196_2 = {c1701};
    Full_Adder FA_4196(s4196, c4196, in4196_1, in4196_2, c1699);
    wire[0:0] s4197, in4197_1, in4197_2;
    wire c4197;
    assign in4197_1 = {s1703[0]};
    assign in4197_2 = {s1704[0]};
    Full_Adder FA_4197(s4197, c4197, in4197_1, in4197_2, s1702[0]);
    wire[0:0] s4198, in4198_1, in4198_2;
    wire c4198;
    assign in4198_1 = {s1706[0]};
    assign in4198_2 = {s1707[0]};
    Full_Adder FA_4198(s4198, c4198, in4198_1, in4198_2, s1705[0]);
    wire[0:0] s4199, in4199_1, in4199_2;
    wire c4199;
    assign in4199_1 = {s1709[0]};
    assign in4199_2 = {s1710[0]};
    Full_Adder FA_4199(s4199, c4199, in4199_1, in4199_2, s1708[0]);
    wire[0:0] s4200, in4200_1, in4200_2;
    wire c4200;
    assign in4200_1 = {s1712[0]};
    assign in4200_2 = {s1713[0]};
    Full_Adder FA_4200(s4200, c4200, in4200_1, in4200_2, s1711[0]);
    wire[0:0] s4201, in4201_1, in4201_2;
    wire c4201;
    assign in4201_1 = {pp70[87]};
    assign in4201_2 = {pp71[86]};
    Full_Adder FA_4201(s4201, c4201, in4201_1, in4201_2, pp69[88]);
    wire[0:0] s4202, in4202_1, in4202_2;
    wire c4202;
    assign in4202_1 = {pp73[84]};
    assign in4202_2 = {pp74[83]};
    Full_Adder FA_4202(s4202, c4202, in4202_1, in4202_2, pp72[85]);
    wire[0:0] s4203, in4203_1, in4203_2;
    wire c4203;
    assign in4203_1 = {pp76[81]};
    assign in4203_2 = {pp77[80]};
    Full_Adder FA_4203(s4203, c4203, in4203_1, in4203_2, pp75[82]);
    wire[0:0] s4204, in4204_1, in4204_2;
    wire c4204;
    assign in4204_1 = {pp79[78]};
    assign in4204_2 = {pp80[77]};
    Full_Adder FA_4204(s4204, c4204, in4204_1, in4204_2, pp78[79]);
    wire[0:0] s4205, in4205_1, in4205_2;
    wire c4205;
    assign in4205_1 = {pp82[75]};
    assign in4205_2 = {pp83[74]};
    Full_Adder FA_4205(s4205, c4205, in4205_1, in4205_2, pp81[76]);
    wire[0:0] s4206, in4206_1, in4206_2;
    wire c4206;
    assign in4206_1 = {pp85[72]};
    assign in4206_2 = {pp86[71]};
    Full_Adder FA_4206(s4206, c4206, in4206_1, in4206_2, pp84[73]);
    wire[0:0] s4207, in4207_1, in4207_2;
    wire c4207;
    assign in4207_1 = {pp88[69]};
    assign in4207_2 = {pp89[68]};
    Full_Adder FA_4207(s4207, c4207, in4207_1, in4207_2, pp87[70]);
    wire[0:0] s4208, in4208_1, in4208_2;
    wire c4208;
    assign in4208_1 = {pp91[66]};
    assign in4208_2 = {pp92[65]};
    Full_Adder FA_4208(s4208, c4208, in4208_1, in4208_2, pp90[67]);
    wire[0:0] s4209, in4209_1, in4209_2;
    wire c4209;
    assign in4209_1 = {pp94[63]};
    assign in4209_2 = {pp95[62]};
    Full_Adder FA_4209(s4209, c4209, in4209_1, in4209_2, pp93[64]);
    wire[0:0] s4210, in4210_1, in4210_2;
    wire c4210;
    assign in4210_1 = {pp97[60]};
    assign in4210_2 = {pp98[59]};
    Full_Adder FA_4210(s4210, c4210, in4210_1, in4210_2, pp96[61]);
    wire[0:0] s4211, in4211_1, in4211_2;
    wire c4211;
    assign in4211_1 = {pp100[57]};
    assign in4211_2 = {pp101[56]};
    Full_Adder FA_4211(s4211, c4211, in4211_1, in4211_2, pp99[58]);
    wire[0:0] s4212, in4212_1, in4212_2;
    wire c4212;
    assign in4212_1 = {pp103[54]};
    assign in4212_2 = {pp104[53]};
    Full_Adder FA_4212(s4212, c4212, in4212_1, in4212_2, pp102[55]);
    wire[0:0] s4213, in4213_1, in4213_2;
    wire c4213;
    assign in4213_1 = {pp106[51]};
    assign in4213_2 = {pp107[50]};
    Full_Adder FA_4213(s4213, c4213, in4213_1, in4213_2, pp105[52]);
    wire[0:0] s4214, in4214_1, in4214_2;
    wire c4214;
    assign in4214_1 = {pp109[48]};
    assign in4214_2 = {pp110[47]};
    Full_Adder FA_4214(s4214, c4214, in4214_1, in4214_2, pp108[49]);
    wire[0:0] s4215, in4215_1, in4215_2;
    wire c4215;
    assign in4215_1 = {pp112[45]};
    assign in4215_2 = {pp113[44]};
    Full_Adder FA_4215(s4215, c4215, in4215_1, in4215_2, pp111[46]);
    wire[0:0] s4216, in4216_1, in4216_2;
    wire c4216;
    assign in4216_1 = {pp115[42]};
    assign in4216_2 = {pp116[41]};
    Full_Adder FA_4216(s4216, c4216, in4216_1, in4216_2, pp114[43]);
    wire[0:0] s4217, in4217_1, in4217_2;
    wire c4217;
    assign in4217_1 = {pp118[39]};
    assign in4217_2 = {pp119[38]};
    Full_Adder FA_4217(s4217, c4217, in4217_1, in4217_2, pp117[40]);
    wire[0:0] s4218, in4218_1, in4218_2;
    wire c4218;
    assign in4218_1 = {pp121[36]};
    assign in4218_2 = {pp122[35]};
    Full_Adder FA_4218(s4218, c4218, in4218_1, in4218_2, pp120[37]);
    wire[0:0] s4219, in4219_1, in4219_2;
    wire c4219;
    assign in4219_1 = {pp124[33]};
    assign in4219_2 = {pp125[32]};
    Full_Adder FA_4219(s4219, c4219, in4219_1, in4219_2, pp123[34]);
    wire[0:0] s4220, in4220_1, in4220_2;
    wire c4220;
    assign in4220_1 = {pp127[30]};
    assign in4220_2 = {c1702};
    Full_Adder FA_4220(s4220, c4220, in4220_1, in4220_2, pp126[31]);
    wire[0:0] s4221, in4221_1, in4221_2;
    wire c4221;
    assign in4221_1 = {c1704};
    assign in4221_2 = {c1705};
    Full_Adder FA_4221(s4221, c4221, in4221_1, in4221_2, c1703);
    wire[0:0] s4222, in4222_1, in4222_2;
    wire c4222;
    assign in4222_1 = {c1707};
    assign in4222_2 = {c1708};
    Full_Adder FA_4222(s4222, c4222, in4222_1, in4222_2, c1706);
    wire[0:0] s4223, in4223_1, in4223_2;
    wire c4223;
    assign in4223_1 = {c1710};
    assign in4223_2 = {c1711};
    Full_Adder FA_4223(s4223, c4223, in4223_1, in4223_2, c1709);
    wire[0:0] s4224, in4224_1, in4224_2;
    wire c4224;
    assign in4224_1 = {c1713};
    assign in4224_2 = {c1714};
    Full_Adder FA_4224(s4224, c4224, in4224_1, in4224_2, c1712);
    wire[0:0] s4225, in4225_1, in4225_2;
    wire c4225;
    assign in4225_1 = {s1716[0]};
    assign in4225_2 = {s1717[0]};
    Full_Adder FA_4225(s4225, c4225, in4225_1, in4225_2, c1715);
    wire[0:0] s4226, in4226_1, in4226_2;
    wire c4226;
    assign in4226_1 = {s1719[0]};
    assign in4226_2 = {s1720[0]};
    Full_Adder FA_4226(s4226, c4226, in4226_1, in4226_2, s1718[0]);
    wire[0:0] s4227, in4227_1, in4227_2;
    wire c4227;
    assign in4227_1 = {s1722[0]};
    assign in4227_2 = {s1723[0]};
    Full_Adder FA_4227(s4227, c4227, in4227_1, in4227_2, s1721[0]);
    wire[0:0] s4228, in4228_1, in4228_2;
    wire c4228;
    assign in4228_1 = {s1725[0]};
    assign in4228_2 = {s1726[0]};
    Full_Adder FA_4228(s4228, c4228, in4228_1, in4228_2, s1724[0]);
    wire[0:0] s4229, in4229_1, in4229_2;
    wire c4229;
    assign in4229_1 = {pp68[90]};
    assign in4229_2 = {pp69[89]};
    Full_Adder FA_4229(s4229, c4229, in4229_1, in4229_2, pp67[91]);
    wire[0:0] s4230, in4230_1, in4230_2;
    wire c4230;
    assign in4230_1 = {pp71[87]};
    assign in4230_2 = {pp72[86]};
    Full_Adder FA_4230(s4230, c4230, in4230_1, in4230_2, pp70[88]);
    wire[0:0] s4231, in4231_1, in4231_2;
    wire c4231;
    assign in4231_1 = {pp74[84]};
    assign in4231_2 = {pp75[83]};
    Full_Adder FA_4231(s4231, c4231, in4231_1, in4231_2, pp73[85]);
    wire[0:0] s4232, in4232_1, in4232_2;
    wire c4232;
    assign in4232_1 = {pp77[81]};
    assign in4232_2 = {pp78[80]};
    Full_Adder FA_4232(s4232, c4232, in4232_1, in4232_2, pp76[82]);
    wire[0:0] s4233, in4233_1, in4233_2;
    wire c4233;
    assign in4233_1 = {pp80[78]};
    assign in4233_2 = {pp81[77]};
    Full_Adder FA_4233(s4233, c4233, in4233_1, in4233_2, pp79[79]);
    wire[0:0] s4234, in4234_1, in4234_2;
    wire c4234;
    assign in4234_1 = {pp83[75]};
    assign in4234_2 = {pp84[74]};
    Full_Adder FA_4234(s4234, c4234, in4234_1, in4234_2, pp82[76]);
    wire[0:0] s4235, in4235_1, in4235_2;
    wire c4235;
    assign in4235_1 = {pp86[72]};
    assign in4235_2 = {pp87[71]};
    Full_Adder FA_4235(s4235, c4235, in4235_1, in4235_2, pp85[73]);
    wire[0:0] s4236, in4236_1, in4236_2;
    wire c4236;
    assign in4236_1 = {pp89[69]};
    assign in4236_2 = {pp90[68]};
    Full_Adder FA_4236(s4236, c4236, in4236_1, in4236_2, pp88[70]);
    wire[0:0] s4237, in4237_1, in4237_2;
    wire c4237;
    assign in4237_1 = {pp92[66]};
    assign in4237_2 = {pp93[65]};
    Full_Adder FA_4237(s4237, c4237, in4237_1, in4237_2, pp91[67]);
    wire[0:0] s4238, in4238_1, in4238_2;
    wire c4238;
    assign in4238_1 = {pp95[63]};
    assign in4238_2 = {pp96[62]};
    Full_Adder FA_4238(s4238, c4238, in4238_1, in4238_2, pp94[64]);
    wire[0:0] s4239, in4239_1, in4239_2;
    wire c4239;
    assign in4239_1 = {pp98[60]};
    assign in4239_2 = {pp99[59]};
    Full_Adder FA_4239(s4239, c4239, in4239_1, in4239_2, pp97[61]);
    wire[0:0] s4240, in4240_1, in4240_2;
    wire c4240;
    assign in4240_1 = {pp101[57]};
    assign in4240_2 = {pp102[56]};
    Full_Adder FA_4240(s4240, c4240, in4240_1, in4240_2, pp100[58]);
    wire[0:0] s4241, in4241_1, in4241_2;
    wire c4241;
    assign in4241_1 = {pp104[54]};
    assign in4241_2 = {pp105[53]};
    Full_Adder FA_4241(s4241, c4241, in4241_1, in4241_2, pp103[55]);
    wire[0:0] s4242, in4242_1, in4242_2;
    wire c4242;
    assign in4242_1 = {pp107[51]};
    assign in4242_2 = {pp108[50]};
    Full_Adder FA_4242(s4242, c4242, in4242_1, in4242_2, pp106[52]);
    wire[0:0] s4243, in4243_1, in4243_2;
    wire c4243;
    assign in4243_1 = {pp110[48]};
    assign in4243_2 = {pp111[47]};
    Full_Adder FA_4243(s4243, c4243, in4243_1, in4243_2, pp109[49]);
    wire[0:0] s4244, in4244_1, in4244_2;
    wire c4244;
    assign in4244_1 = {pp113[45]};
    assign in4244_2 = {pp114[44]};
    Full_Adder FA_4244(s4244, c4244, in4244_1, in4244_2, pp112[46]);
    wire[0:0] s4245, in4245_1, in4245_2;
    wire c4245;
    assign in4245_1 = {pp116[42]};
    assign in4245_2 = {pp117[41]};
    Full_Adder FA_4245(s4245, c4245, in4245_1, in4245_2, pp115[43]);
    wire[0:0] s4246, in4246_1, in4246_2;
    wire c4246;
    assign in4246_1 = {pp119[39]};
    assign in4246_2 = {pp120[38]};
    Full_Adder FA_4246(s4246, c4246, in4246_1, in4246_2, pp118[40]);
    wire[0:0] s4247, in4247_1, in4247_2;
    wire c4247;
    assign in4247_1 = {pp122[36]};
    assign in4247_2 = {pp123[35]};
    Full_Adder FA_4247(s4247, c4247, in4247_1, in4247_2, pp121[37]);
    wire[0:0] s4248, in4248_1, in4248_2;
    wire c4248;
    assign in4248_1 = {pp125[33]};
    assign in4248_2 = {pp126[32]};
    Full_Adder FA_4248(s4248, c4248, in4248_1, in4248_2, pp124[34]);
    wire[0:0] s4249, in4249_1, in4249_2;
    wire c4249;
    assign in4249_1 = {c1716};
    assign in4249_2 = {c1717};
    Full_Adder FA_4249(s4249, c4249, in4249_1, in4249_2, pp127[31]);
    wire[0:0] s4250, in4250_1, in4250_2;
    wire c4250;
    assign in4250_1 = {c1719};
    assign in4250_2 = {c1720};
    Full_Adder FA_4250(s4250, c4250, in4250_1, in4250_2, c1718);
    wire[0:0] s4251, in4251_1, in4251_2;
    wire c4251;
    assign in4251_1 = {c1722};
    assign in4251_2 = {c1723};
    Full_Adder FA_4251(s4251, c4251, in4251_1, in4251_2, c1721);
    wire[0:0] s4252, in4252_1, in4252_2;
    wire c4252;
    assign in4252_1 = {c1725};
    assign in4252_2 = {c1726};
    Full_Adder FA_4252(s4252, c4252, in4252_1, in4252_2, c1724);
    wire[0:0] s4253, in4253_1, in4253_2;
    wire c4253;
    assign in4253_1 = {c1728};
    assign in4253_2 = {s1729[0]};
    Full_Adder FA_4253(s4253, c4253, in4253_1, in4253_2, c1727);
    wire[0:0] s4254, in4254_1, in4254_2;
    wire c4254;
    assign in4254_1 = {s1731[0]};
    assign in4254_2 = {s1732[0]};
    Full_Adder FA_4254(s4254, c4254, in4254_1, in4254_2, s1730[0]);
    wire[0:0] s4255, in4255_1, in4255_2;
    wire c4255;
    assign in4255_1 = {s1734[0]};
    assign in4255_2 = {s1735[0]};
    Full_Adder FA_4255(s4255, c4255, in4255_1, in4255_2, s1733[0]);
    wire[0:0] s4256, in4256_1, in4256_2;
    wire c4256;
    assign in4256_1 = {s1737[0]};
    assign in4256_2 = {s1738[0]};
    Full_Adder FA_4256(s4256, c4256, in4256_1, in4256_2, s1736[0]);
    wire[0:0] s4257, in4257_1, in4257_2;
    wire c4257;
    assign in4257_1 = {pp66[93]};
    assign in4257_2 = {pp67[92]};
    Full_Adder FA_4257(s4257, c4257, in4257_1, in4257_2, pp65[94]);
    wire[0:0] s4258, in4258_1, in4258_2;
    wire c4258;
    assign in4258_1 = {pp69[90]};
    assign in4258_2 = {pp70[89]};
    Full_Adder FA_4258(s4258, c4258, in4258_1, in4258_2, pp68[91]);
    wire[0:0] s4259, in4259_1, in4259_2;
    wire c4259;
    assign in4259_1 = {pp72[87]};
    assign in4259_2 = {pp73[86]};
    Full_Adder FA_4259(s4259, c4259, in4259_1, in4259_2, pp71[88]);
    wire[0:0] s4260, in4260_1, in4260_2;
    wire c4260;
    assign in4260_1 = {pp75[84]};
    assign in4260_2 = {pp76[83]};
    Full_Adder FA_4260(s4260, c4260, in4260_1, in4260_2, pp74[85]);
    wire[0:0] s4261, in4261_1, in4261_2;
    wire c4261;
    assign in4261_1 = {pp78[81]};
    assign in4261_2 = {pp79[80]};
    Full_Adder FA_4261(s4261, c4261, in4261_1, in4261_2, pp77[82]);
    wire[0:0] s4262, in4262_1, in4262_2;
    wire c4262;
    assign in4262_1 = {pp81[78]};
    assign in4262_2 = {pp82[77]};
    Full_Adder FA_4262(s4262, c4262, in4262_1, in4262_2, pp80[79]);
    wire[0:0] s4263, in4263_1, in4263_2;
    wire c4263;
    assign in4263_1 = {pp84[75]};
    assign in4263_2 = {pp85[74]};
    Full_Adder FA_4263(s4263, c4263, in4263_1, in4263_2, pp83[76]);
    wire[0:0] s4264, in4264_1, in4264_2;
    wire c4264;
    assign in4264_1 = {pp87[72]};
    assign in4264_2 = {pp88[71]};
    Full_Adder FA_4264(s4264, c4264, in4264_1, in4264_2, pp86[73]);
    wire[0:0] s4265, in4265_1, in4265_2;
    wire c4265;
    assign in4265_1 = {pp90[69]};
    assign in4265_2 = {pp91[68]};
    Full_Adder FA_4265(s4265, c4265, in4265_1, in4265_2, pp89[70]);
    wire[0:0] s4266, in4266_1, in4266_2;
    wire c4266;
    assign in4266_1 = {pp93[66]};
    assign in4266_2 = {pp94[65]};
    Full_Adder FA_4266(s4266, c4266, in4266_1, in4266_2, pp92[67]);
    wire[0:0] s4267, in4267_1, in4267_2;
    wire c4267;
    assign in4267_1 = {pp96[63]};
    assign in4267_2 = {pp97[62]};
    Full_Adder FA_4267(s4267, c4267, in4267_1, in4267_2, pp95[64]);
    wire[0:0] s4268, in4268_1, in4268_2;
    wire c4268;
    assign in4268_1 = {pp99[60]};
    assign in4268_2 = {pp100[59]};
    Full_Adder FA_4268(s4268, c4268, in4268_1, in4268_2, pp98[61]);
    wire[0:0] s4269, in4269_1, in4269_2;
    wire c4269;
    assign in4269_1 = {pp102[57]};
    assign in4269_2 = {pp103[56]};
    Full_Adder FA_4269(s4269, c4269, in4269_1, in4269_2, pp101[58]);
    wire[0:0] s4270, in4270_1, in4270_2;
    wire c4270;
    assign in4270_1 = {pp105[54]};
    assign in4270_2 = {pp106[53]};
    Full_Adder FA_4270(s4270, c4270, in4270_1, in4270_2, pp104[55]);
    wire[0:0] s4271, in4271_1, in4271_2;
    wire c4271;
    assign in4271_1 = {pp108[51]};
    assign in4271_2 = {pp109[50]};
    Full_Adder FA_4271(s4271, c4271, in4271_1, in4271_2, pp107[52]);
    wire[0:0] s4272, in4272_1, in4272_2;
    wire c4272;
    assign in4272_1 = {pp111[48]};
    assign in4272_2 = {pp112[47]};
    Full_Adder FA_4272(s4272, c4272, in4272_1, in4272_2, pp110[49]);
    wire[0:0] s4273, in4273_1, in4273_2;
    wire c4273;
    assign in4273_1 = {pp114[45]};
    assign in4273_2 = {pp115[44]};
    Full_Adder FA_4273(s4273, c4273, in4273_1, in4273_2, pp113[46]);
    wire[0:0] s4274, in4274_1, in4274_2;
    wire c4274;
    assign in4274_1 = {pp117[42]};
    assign in4274_2 = {pp118[41]};
    Full_Adder FA_4274(s4274, c4274, in4274_1, in4274_2, pp116[43]);
    wire[0:0] s4275, in4275_1, in4275_2;
    wire c4275;
    assign in4275_1 = {pp120[39]};
    assign in4275_2 = {pp121[38]};
    Full_Adder FA_4275(s4275, c4275, in4275_1, in4275_2, pp119[40]);
    wire[0:0] s4276, in4276_1, in4276_2;
    wire c4276;
    assign in4276_1 = {pp123[36]};
    assign in4276_2 = {pp124[35]};
    Full_Adder FA_4276(s4276, c4276, in4276_1, in4276_2, pp122[37]);
    wire[0:0] s4277, in4277_1, in4277_2;
    wire c4277;
    assign in4277_1 = {pp126[33]};
    assign in4277_2 = {pp127[32]};
    Full_Adder FA_4277(s4277, c4277, in4277_1, in4277_2, pp125[34]);
    wire[0:0] s4278, in4278_1, in4278_2;
    wire c4278;
    assign in4278_1 = {c1730};
    assign in4278_2 = {c1731};
    Full_Adder FA_4278(s4278, c4278, in4278_1, in4278_2, c1729);
    wire[0:0] s4279, in4279_1, in4279_2;
    wire c4279;
    assign in4279_1 = {c1733};
    assign in4279_2 = {c1734};
    Full_Adder FA_4279(s4279, c4279, in4279_1, in4279_2, c1732);
    wire[0:0] s4280, in4280_1, in4280_2;
    wire c4280;
    assign in4280_1 = {c1736};
    assign in4280_2 = {c1737};
    Full_Adder FA_4280(s4280, c4280, in4280_1, in4280_2, c1735);
    wire[0:0] s4281, in4281_1, in4281_2;
    wire c4281;
    assign in4281_1 = {c1739};
    assign in4281_2 = {c1740};
    Full_Adder FA_4281(s4281, c4281, in4281_1, in4281_2, c1738);
    wire[0:0] s4282, in4282_1, in4282_2;
    wire c4282;
    assign in4282_1 = {s1742[0]};
    assign in4282_2 = {s1743[0]};
    Full_Adder FA_4282(s4282, c4282, in4282_1, in4282_2, s1741[0]);
    wire[0:0] s4283, in4283_1, in4283_2;
    wire c4283;
    assign in4283_1 = {s1745[0]};
    assign in4283_2 = {s1746[0]};
    Full_Adder FA_4283(s4283, c4283, in4283_1, in4283_2, s1744[0]);
    wire[0:0] s4284, in4284_1, in4284_2;
    wire c4284;
    assign in4284_1 = {s1748[0]};
    assign in4284_2 = {s1749[0]};
    Full_Adder FA_4284(s4284, c4284, in4284_1, in4284_2, s1747[0]);
    wire[0:0] s4285, in4285_1, in4285_2;
    wire c4285;
    assign in4285_1 = {pp64[96]};
    assign in4285_2 = {pp65[95]};
    Full_Adder FA_4285(s4285, c4285, in4285_1, in4285_2, pp63[97]);
    wire[0:0] s4286, in4286_1, in4286_2;
    wire c4286;
    assign in4286_1 = {pp67[93]};
    assign in4286_2 = {pp68[92]};
    Full_Adder FA_4286(s4286, c4286, in4286_1, in4286_2, pp66[94]);
    wire[0:0] s4287, in4287_1, in4287_2;
    wire c4287;
    assign in4287_1 = {pp70[90]};
    assign in4287_2 = {pp71[89]};
    Full_Adder FA_4287(s4287, c4287, in4287_1, in4287_2, pp69[91]);
    wire[0:0] s4288, in4288_1, in4288_2;
    wire c4288;
    assign in4288_1 = {pp73[87]};
    assign in4288_2 = {pp74[86]};
    Full_Adder FA_4288(s4288, c4288, in4288_1, in4288_2, pp72[88]);
    wire[0:0] s4289, in4289_1, in4289_2;
    wire c4289;
    assign in4289_1 = {pp76[84]};
    assign in4289_2 = {pp77[83]};
    Full_Adder FA_4289(s4289, c4289, in4289_1, in4289_2, pp75[85]);
    wire[0:0] s4290, in4290_1, in4290_2;
    wire c4290;
    assign in4290_1 = {pp79[81]};
    assign in4290_2 = {pp80[80]};
    Full_Adder FA_4290(s4290, c4290, in4290_1, in4290_2, pp78[82]);
    wire[0:0] s4291, in4291_1, in4291_2;
    wire c4291;
    assign in4291_1 = {pp82[78]};
    assign in4291_2 = {pp83[77]};
    Full_Adder FA_4291(s4291, c4291, in4291_1, in4291_2, pp81[79]);
    wire[0:0] s4292, in4292_1, in4292_2;
    wire c4292;
    assign in4292_1 = {pp85[75]};
    assign in4292_2 = {pp86[74]};
    Full_Adder FA_4292(s4292, c4292, in4292_1, in4292_2, pp84[76]);
    wire[0:0] s4293, in4293_1, in4293_2;
    wire c4293;
    assign in4293_1 = {pp88[72]};
    assign in4293_2 = {pp89[71]};
    Full_Adder FA_4293(s4293, c4293, in4293_1, in4293_2, pp87[73]);
    wire[0:0] s4294, in4294_1, in4294_2;
    wire c4294;
    assign in4294_1 = {pp91[69]};
    assign in4294_2 = {pp92[68]};
    Full_Adder FA_4294(s4294, c4294, in4294_1, in4294_2, pp90[70]);
    wire[0:0] s4295, in4295_1, in4295_2;
    wire c4295;
    assign in4295_1 = {pp94[66]};
    assign in4295_2 = {pp95[65]};
    Full_Adder FA_4295(s4295, c4295, in4295_1, in4295_2, pp93[67]);
    wire[0:0] s4296, in4296_1, in4296_2;
    wire c4296;
    assign in4296_1 = {pp97[63]};
    assign in4296_2 = {pp98[62]};
    Full_Adder FA_4296(s4296, c4296, in4296_1, in4296_2, pp96[64]);
    wire[0:0] s4297, in4297_1, in4297_2;
    wire c4297;
    assign in4297_1 = {pp100[60]};
    assign in4297_2 = {pp101[59]};
    Full_Adder FA_4297(s4297, c4297, in4297_1, in4297_2, pp99[61]);
    wire[0:0] s4298, in4298_1, in4298_2;
    wire c4298;
    assign in4298_1 = {pp103[57]};
    assign in4298_2 = {pp104[56]};
    Full_Adder FA_4298(s4298, c4298, in4298_1, in4298_2, pp102[58]);
    wire[0:0] s4299, in4299_1, in4299_2;
    wire c4299;
    assign in4299_1 = {pp106[54]};
    assign in4299_2 = {pp107[53]};
    Full_Adder FA_4299(s4299, c4299, in4299_1, in4299_2, pp105[55]);
    wire[0:0] s4300, in4300_1, in4300_2;
    wire c4300;
    assign in4300_1 = {pp109[51]};
    assign in4300_2 = {pp110[50]};
    Full_Adder FA_4300(s4300, c4300, in4300_1, in4300_2, pp108[52]);
    wire[0:0] s4301, in4301_1, in4301_2;
    wire c4301;
    assign in4301_1 = {pp112[48]};
    assign in4301_2 = {pp113[47]};
    Full_Adder FA_4301(s4301, c4301, in4301_1, in4301_2, pp111[49]);
    wire[0:0] s4302, in4302_1, in4302_2;
    wire c4302;
    assign in4302_1 = {pp115[45]};
    assign in4302_2 = {pp116[44]};
    Full_Adder FA_4302(s4302, c4302, in4302_1, in4302_2, pp114[46]);
    wire[0:0] s4303, in4303_1, in4303_2;
    wire c4303;
    assign in4303_1 = {pp118[42]};
    assign in4303_2 = {pp119[41]};
    Full_Adder FA_4303(s4303, c4303, in4303_1, in4303_2, pp117[43]);
    wire[0:0] s4304, in4304_1, in4304_2;
    wire c4304;
    assign in4304_1 = {pp121[39]};
    assign in4304_2 = {pp122[38]};
    Full_Adder FA_4304(s4304, c4304, in4304_1, in4304_2, pp120[40]);
    wire[0:0] s4305, in4305_1, in4305_2;
    wire c4305;
    assign in4305_1 = {pp124[36]};
    assign in4305_2 = {pp125[35]};
    Full_Adder FA_4305(s4305, c4305, in4305_1, in4305_2, pp123[37]);
    wire[0:0] s4306, in4306_1, in4306_2;
    wire c4306;
    assign in4306_1 = {pp127[33]};
    assign in4306_2 = {c1741};
    Full_Adder FA_4306(s4306, c4306, in4306_1, in4306_2, pp126[34]);
    wire[0:0] s4307, in4307_1, in4307_2;
    wire c4307;
    assign in4307_1 = {c1743};
    assign in4307_2 = {c1744};
    Full_Adder FA_4307(s4307, c4307, in4307_1, in4307_2, c1742);
    wire[0:0] s4308, in4308_1, in4308_2;
    wire c4308;
    assign in4308_1 = {c1746};
    assign in4308_2 = {c1747};
    Full_Adder FA_4308(s4308, c4308, in4308_1, in4308_2, c1745);
    wire[0:0] s4309, in4309_1, in4309_2;
    wire c4309;
    assign in4309_1 = {c1749};
    assign in4309_2 = {c1750};
    Full_Adder FA_4309(s4309, c4309, in4309_1, in4309_2, c1748);
    wire[0:0] s4310, in4310_1, in4310_2;
    wire c4310;
    assign in4310_1 = {s1752[0]};
    assign in4310_2 = {s1753[0]};
    Full_Adder FA_4310(s4310, c4310, in4310_1, in4310_2, c1751);
    wire[0:0] s4311, in4311_1, in4311_2;
    wire c4311;
    assign in4311_1 = {s1755[0]};
    assign in4311_2 = {s1756[0]};
    Full_Adder FA_4311(s4311, c4311, in4311_1, in4311_2, s1754[0]);
    wire[0:0] s4312, in4312_1, in4312_2;
    wire c4312;
    assign in4312_1 = {s1758[0]};
    assign in4312_2 = {s1759[0]};
    Full_Adder FA_4312(s4312, c4312, in4312_1, in4312_2, s1757[0]);
    wire[0:0] s4313, in4313_1, in4313_2;
    wire c4313;
    assign in4313_1 = {pp62[99]};
    assign in4313_2 = {pp63[98]};
    Full_Adder FA_4313(s4313, c4313, in4313_1, in4313_2, pp61[100]);
    wire[0:0] s4314, in4314_1, in4314_2;
    wire c4314;
    assign in4314_1 = {pp65[96]};
    assign in4314_2 = {pp66[95]};
    Full_Adder FA_4314(s4314, c4314, in4314_1, in4314_2, pp64[97]);
    wire[0:0] s4315, in4315_1, in4315_2;
    wire c4315;
    assign in4315_1 = {pp68[93]};
    assign in4315_2 = {pp69[92]};
    Full_Adder FA_4315(s4315, c4315, in4315_1, in4315_2, pp67[94]);
    wire[0:0] s4316, in4316_1, in4316_2;
    wire c4316;
    assign in4316_1 = {pp71[90]};
    assign in4316_2 = {pp72[89]};
    Full_Adder FA_4316(s4316, c4316, in4316_1, in4316_2, pp70[91]);
    wire[0:0] s4317, in4317_1, in4317_2;
    wire c4317;
    assign in4317_1 = {pp74[87]};
    assign in4317_2 = {pp75[86]};
    Full_Adder FA_4317(s4317, c4317, in4317_1, in4317_2, pp73[88]);
    wire[0:0] s4318, in4318_1, in4318_2;
    wire c4318;
    assign in4318_1 = {pp77[84]};
    assign in4318_2 = {pp78[83]};
    Full_Adder FA_4318(s4318, c4318, in4318_1, in4318_2, pp76[85]);
    wire[0:0] s4319, in4319_1, in4319_2;
    wire c4319;
    assign in4319_1 = {pp80[81]};
    assign in4319_2 = {pp81[80]};
    Full_Adder FA_4319(s4319, c4319, in4319_1, in4319_2, pp79[82]);
    wire[0:0] s4320, in4320_1, in4320_2;
    wire c4320;
    assign in4320_1 = {pp83[78]};
    assign in4320_2 = {pp84[77]};
    Full_Adder FA_4320(s4320, c4320, in4320_1, in4320_2, pp82[79]);
    wire[0:0] s4321, in4321_1, in4321_2;
    wire c4321;
    assign in4321_1 = {pp86[75]};
    assign in4321_2 = {pp87[74]};
    Full_Adder FA_4321(s4321, c4321, in4321_1, in4321_2, pp85[76]);
    wire[0:0] s4322, in4322_1, in4322_2;
    wire c4322;
    assign in4322_1 = {pp89[72]};
    assign in4322_2 = {pp90[71]};
    Full_Adder FA_4322(s4322, c4322, in4322_1, in4322_2, pp88[73]);
    wire[0:0] s4323, in4323_1, in4323_2;
    wire c4323;
    assign in4323_1 = {pp92[69]};
    assign in4323_2 = {pp93[68]};
    Full_Adder FA_4323(s4323, c4323, in4323_1, in4323_2, pp91[70]);
    wire[0:0] s4324, in4324_1, in4324_2;
    wire c4324;
    assign in4324_1 = {pp95[66]};
    assign in4324_2 = {pp96[65]};
    Full_Adder FA_4324(s4324, c4324, in4324_1, in4324_2, pp94[67]);
    wire[0:0] s4325, in4325_1, in4325_2;
    wire c4325;
    assign in4325_1 = {pp98[63]};
    assign in4325_2 = {pp99[62]};
    Full_Adder FA_4325(s4325, c4325, in4325_1, in4325_2, pp97[64]);
    wire[0:0] s4326, in4326_1, in4326_2;
    wire c4326;
    assign in4326_1 = {pp101[60]};
    assign in4326_2 = {pp102[59]};
    Full_Adder FA_4326(s4326, c4326, in4326_1, in4326_2, pp100[61]);
    wire[0:0] s4327, in4327_1, in4327_2;
    wire c4327;
    assign in4327_1 = {pp104[57]};
    assign in4327_2 = {pp105[56]};
    Full_Adder FA_4327(s4327, c4327, in4327_1, in4327_2, pp103[58]);
    wire[0:0] s4328, in4328_1, in4328_2;
    wire c4328;
    assign in4328_1 = {pp107[54]};
    assign in4328_2 = {pp108[53]};
    Full_Adder FA_4328(s4328, c4328, in4328_1, in4328_2, pp106[55]);
    wire[0:0] s4329, in4329_1, in4329_2;
    wire c4329;
    assign in4329_1 = {pp110[51]};
    assign in4329_2 = {pp111[50]};
    Full_Adder FA_4329(s4329, c4329, in4329_1, in4329_2, pp109[52]);
    wire[0:0] s4330, in4330_1, in4330_2;
    wire c4330;
    assign in4330_1 = {pp113[48]};
    assign in4330_2 = {pp114[47]};
    Full_Adder FA_4330(s4330, c4330, in4330_1, in4330_2, pp112[49]);
    wire[0:0] s4331, in4331_1, in4331_2;
    wire c4331;
    assign in4331_1 = {pp116[45]};
    assign in4331_2 = {pp117[44]};
    Full_Adder FA_4331(s4331, c4331, in4331_1, in4331_2, pp115[46]);
    wire[0:0] s4332, in4332_1, in4332_2;
    wire c4332;
    assign in4332_1 = {pp119[42]};
    assign in4332_2 = {pp120[41]};
    Full_Adder FA_4332(s4332, c4332, in4332_1, in4332_2, pp118[43]);
    wire[0:0] s4333, in4333_1, in4333_2;
    wire c4333;
    assign in4333_1 = {pp122[39]};
    assign in4333_2 = {pp123[38]};
    Full_Adder FA_4333(s4333, c4333, in4333_1, in4333_2, pp121[40]);
    wire[0:0] s4334, in4334_1, in4334_2;
    wire c4334;
    assign in4334_1 = {pp125[36]};
    assign in4334_2 = {pp126[35]};
    Full_Adder FA_4334(s4334, c4334, in4334_1, in4334_2, pp124[37]);
    wire[0:0] s4335, in4335_1, in4335_2;
    wire c4335;
    assign in4335_1 = {c1752};
    assign in4335_2 = {c1753};
    Full_Adder FA_4335(s4335, c4335, in4335_1, in4335_2, pp127[34]);
    wire[0:0] s4336, in4336_1, in4336_2;
    wire c4336;
    assign in4336_1 = {c1755};
    assign in4336_2 = {c1756};
    Full_Adder FA_4336(s4336, c4336, in4336_1, in4336_2, c1754);
    wire[0:0] s4337, in4337_1, in4337_2;
    wire c4337;
    assign in4337_1 = {c1758};
    assign in4337_2 = {c1759};
    Full_Adder FA_4337(s4337, c4337, in4337_1, in4337_2, c1757);
    wire[0:0] s4338, in4338_1, in4338_2;
    wire c4338;
    assign in4338_1 = {c1761};
    assign in4338_2 = {s1762[0]};
    Full_Adder FA_4338(s4338, c4338, in4338_1, in4338_2, c1760);
    wire[0:0] s4339, in4339_1, in4339_2;
    wire c4339;
    assign in4339_1 = {s1764[0]};
    assign in4339_2 = {s1765[0]};
    Full_Adder FA_4339(s4339, c4339, in4339_1, in4339_2, s1763[0]);
    wire[0:0] s4340, in4340_1, in4340_2;
    wire c4340;
    assign in4340_1 = {s1767[0]};
    assign in4340_2 = {s1768[0]};
    Full_Adder FA_4340(s4340, c4340, in4340_1, in4340_2, s1766[0]);
    wire[0:0] s4341, in4341_1, in4341_2;
    wire c4341;
    assign in4341_1 = {pp60[102]};
    assign in4341_2 = {pp61[101]};
    Full_Adder FA_4341(s4341, c4341, in4341_1, in4341_2, pp59[103]);
    wire[0:0] s4342, in4342_1, in4342_2;
    wire c4342;
    assign in4342_1 = {pp63[99]};
    assign in4342_2 = {pp64[98]};
    Full_Adder FA_4342(s4342, c4342, in4342_1, in4342_2, pp62[100]);
    wire[0:0] s4343, in4343_1, in4343_2;
    wire c4343;
    assign in4343_1 = {pp66[96]};
    assign in4343_2 = {pp67[95]};
    Full_Adder FA_4343(s4343, c4343, in4343_1, in4343_2, pp65[97]);
    wire[0:0] s4344, in4344_1, in4344_2;
    wire c4344;
    assign in4344_1 = {pp69[93]};
    assign in4344_2 = {pp70[92]};
    Full_Adder FA_4344(s4344, c4344, in4344_1, in4344_2, pp68[94]);
    wire[0:0] s4345, in4345_1, in4345_2;
    wire c4345;
    assign in4345_1 = {pp72[90]};
    assign in4345_2 = {pp73[89]};
    Full_Adder FA_4345(s4345, c4345, in4345_1, in4345_2, pp71[91]);
    wire[0:0] s4346, in4346_1, in4346_2;
    wire c4346;
    assign in4346_1 = {pp75[87]};
    assign in4346_2 = {pp76[86]};
    Full_Adder FA_4346(s4346, c4346, in4346_1, in4346_2, pp74[88]);
    wire[0:0] s4347, in4347_1, in4347_2;
    wire c4347;
    assign in4347_1 = {pp78[84]};
    assign in4347_2 = {pp79[83]};
    Full_Adder FA_4347(s4347, c4347, in4347_1, in4347_2, pp77[85]);
    wire[0:0] s4348, in4348_1, in4348_2;
    wire c4348;
    assign in4348_1 = {pp81[81]};
    assign in4348_2 = {pp82[80]};
    Full_Adder FA_4348(s4348, c4348, in4348_1, in4348_2, pp80[82]);
    wire[0:0] s4349, in4349_1, in4349_2;
    wire c4349;
    assign in4349_1 = {pp84[78]};
    assign in4349_2 = {pp85[77]};
    Full_Adder FA_4349(s4349, c4349, in4349_1, in4349_2, pp83[79]);
    wire[0:0] s4350, in4350_1, in4350_2;
    wire c4350;
    assign in4350_1 = {pp87[75]};
    assign in4350_2 = {pp88[74]};
    Full_Adder FA_4350(s4350, c4350, in4350_1, in4350_2, pp86[76]);
    wire[0:0] s4351, in4351_1, in4351_2;
    wire c4351;
    assign in4351_1 = {pp90[72]};
    assign in4351_2 = {pp91[71]};
    Full_Adder FA_4351(s4351, c4351, in4351_1, in4351_2, pp89[73]);
    wire[0:0] s4352, in4352_1, in4352_2;
    wire c4352;
    assign in4352_1 = {pp93[69]};
    assign in4352_2 = {pp94[68]};
    Full_Adder FA_4352(s4352, c4352, in4352_1, in4352_2, pp92[70]);
    wire[0:0] s4353, in4353_1, in4353_2;
    wire c4353;
    assign in4353_1 = {pp96[66]};
    assign in4353_2 = {pp97[65]};
    Full_Adder FA_4353(s4353, c4353, in4353_1, in4353_2, pp95[67]);
    wire[0:0] s4354, in4354_1, in4354_2;
    wire c4354;
    assign in4354_1 = {pp99[63]};
    assign in4354_2 = {pp100[62]};
    Full_Adder FA_4354(s4354, c4354, in4354_1, in4354_2, pp98[64]);
    wire[0:0] s4355, in4355_1, in4355_2;
    wire c4355;
    assign in4355_1 = {pp102[60]};
    assign in4355_2 = {pp103[59]};
    Full_Adder FA_4355(s4355, c4355, in4355_1, in4355_2, pp101[61]);
    wire[0:0] s4356, in4356_1, in4356_2;
    wire c4356;
    assign in4356_1 = {pp105[57]};
    assign in4356_2 = {pp106[56]};
    Full_Adder FA_4356(s4356, c4356, in4356_1, in4356_2, pp104[58]);
    wire[0:0] s4357, in4357_1, in4357_2;
    wire c4357;
    assign in4357_1 = {pp108[54]};
    assign in4357_2 = {pp109[53]};
    Full_Adder FA_4357(s4357, c4357, in4357_1, in4357_2, pp107[55]);
    wire[0:0] s4358, in4358_1, in4358_2;
    wire c4358;
    assign in4358_1 = {pp111[51]};
    assign in4358_2 = {pp112[50]};
    Full_Adder FA_4358(s4358, c4358, in4358_1, in4358_2, pp110[52]);
    wire[0:0] s4359, in4359_1, in4359_2;
    wire c4359;
    assign in4359_1 = {pp114[48]};
    assign in4359_2 = {pp115[47]};
    Full_Adder FA_4359(s4359, c4359, in4359_1, in4359_2, pp113[49]);
    wire[0:0] s4360, in4360_1, in4360_2;
    wire c4360;
    assign in4360_1 = {pp117[45]};
    assign in4360_2 = {pp118[44]};
    Full_Adder FA_4360(s4360, c4360, in4360_1, in4360_2, pp116[46]);
    wire[0:0] s4361, in4361_1, in4361_2;
    wire c4361;
    assign in4361_1 = {pp120[42]};
    assign in4361_2 = {pp121[41]};
    Full_Adder FA_4361(s4361, c4361, in4361_1, in4361_2, pp119[43]);
    wire[0:0] s4362, in4362_1, in4362_2;
    wire c4362;
    assign in4362_1 = {pp123[39]};
    assign in4362_2 = {pp124[38]};
    Full_Adder FA_4362(s4362, c4362, in4362_1, in4362_2, pp122[40]);
    wire[0:0] s4363, in4363_1, in4363_2;
    wire c4363;
    assign in4363_1 = {pp126[36]};
    assign in4363_2 = {pp127[35]};
    Full_Adder FA_4363(s4363, c4363, in4363_1, in4363_2, pp125[37]);
    wire[0:0] s4364, in4364_1, in4364_2;
    wire c4364;
    assign in4364_1 = {c1763};
    assign in4364_2 = {c1764};
    Full_Adder FA_4364(s4364, c4364, in4364_1, in4364_2, c1762);
    wire[0:0] s4365, in4365_1, in4365_2;
    wire c4365;
    assign in4365_1 = {c1766};
    assign in4365_2 = {c1767};
    Full_Adder FA_4365(s4365, c4365, in4365_1, in4365_2, c1765);
    wire[0:0] s4366, in4366_1, in4366_2;
    wire c4366;
    assign in4366_1 = {c1769};
    assign in4366_2 = {c1770};
    Full_Adder FA_4366(s4366, c4366, in4366_1, in4366_2, c1768);
    wire[0:0] s4367, in4367_1, in4367_2;
    wire c4367;
    assign in4367_1 = {s1772[0]};
    assign in4367_2 = {s1773[0]};
    Full_Adder FA_4367(s4367, c4367, in4367_1, in4367_2, s1771[0]);
    wire[0:0] s4368, in4368_1, in4368_2;
    wire c4368;
    assign in4368_1 = {s1775[0]};
    assign in4368_2 = {s1776[0]};
    Full_Adder FA_4368(s4368, c4368, in4368_1, in4368_2, s1774[0]);
    wire[0:0] s4369, in4369_1, in4369_2;
    wire c4369;
    assign in4369_1 = {pp58[105]};
    assign in4369_2 = {pp59[104]};
    Full_Adder FA_4369(s4369, c4369, in4369_1, in4369_2, pp57[106]);
    wire[0:0] s4370, in4370_1, in4370_2;
    wire c4370;
    assign in4370_1 = {pp61[102]};
    assign in4370_2 = {pp62[101]};
    Full_Adder FA_4370(s4370, c4370, in4370_1, in4370_2, pp60[103]);
    wire[0:0] s4371, in4371_1, in4371_2;
    wire c4371;
    assign in4371_1 = {pp64[99]};
    assign in4371_2 = {pp65[98]};
    Full_Adder FA_4371(s4371, c4371, in4371_1, in4371_2, pp63[100]);
    wire[0:0] s4372, in4372_1, in4372_2;
    wire c4372;
    assign in4372_1 = {pp67[96]};
    assign in4372_2 = {pp68[95]};
    Full_Adder FA_4372(s4372, c4372, in4372_1, in4372_2, pp66[97]);
    wire[0:0] s4373, in4373_1, in4373_2;
    wire c4373;
    assign in4373_1 = {pp70[93]};
    assign in4373_2 = {pp71[92]};
    Full_Adder FA_4373(s4373, c4373, in4373_1, in4373_2, pp69[94]);
    wire[0:0] s4374, in4374_1, in4374_2;
    wire c4374;
    assign in4374_1 = {pp73[90]};
    assign in4374_2 = {pp74[89]};
    Full_Adder FA_4374(s4374, c4374, in4374_1, in4374_2, pp72[91]);
    wire[0:0] s4375, in4375_1, in4375_2;
    wire c4375;
    assign in4375_1 = {pp76[87]};
    assign in4375_2 = {pp77[86]};
    Full_Adder FA_4375(s4375, c4375, in4375_1, in4375_2, pp75[88]);
    wire[0:0] s4376, in4376_1, in4376_2;
    wire c4376;
    assign in4376_1 = {pp79[84]};
    assign in4376_2 = {pp80[83]};
    Full_Adder FA_4376(s4376, c4376, in4376_1, in4376_2, pp78[85]);
    wire[0:0] s4377, in4377_1, in4377_2;
    wire c4377;
    assign in4377_1 = {pp82[81]};
    assign in4377_2 = {pp83[80]};
    Full_Adder FA_4377(s4377, c4377, in4377_1, in4377_2, pp81[82]);
    wire[0:0] s4378, in4378_1, in4378_2;
    wire c4378;
    assign in4378_1 = {pp85[78]};
    assign in4378_2 = {pp86[77]};
    Full_Adder FA_4378(s4378, c4378, in4378_1, in4378_2, pp84[79]);
    wire[0:0] s4379, in4379_1, in4379_2;
    wire c4379;
    assign in4379_1 = {pp88[75]};
    assign in4379_2 = {pp89[74]};
    Full_Adder FA_4379(s4379, c4379, in4379_1, in4379_2, pp87[76]);
    wire[0:0] s4380, in4380_1, in4380_2;
    wire c4380;
    assign in4380_1 = {pp91[72]};
    assign in4380_2 = {pp92[71]};
    Full_Adder FA_4380(s4380, c4380, in4380_1, in4380_2, pp90[73]);
    wire[0:0] s4381, in4381_1, in4381_2;
    wire c4381;
    assign in4381_1 = {pp94[69]};
    assign in4381_2 = {pp95[68]};
    Full_Adder FA_4381(s4381, c4381, in4381_1, in4381_2, pp93[70]);
    wire[0:0] s4382, in4382_1, in4382_2;
    wire c4382;
    assign in4382_1 = {pp97[66]};
    assign in4382_2 = {pp98[65]};
    Full_Adder FA_4382(s4382, c4382, in4382_1, in4382_2, pp96[67]);
    wire[0:0] s4383, in4383_1, in4383_2;
    wire c4383;
    assign in4383_1 = {pp100[63]};
    assign in4383_2 = {pp101[62]};
    Full_Adder FA_4383(s4383, c4383, in4383_1, in4383_2, pp99[64]);
    wire[0:0] s4384, in4384_1, in4384_2;
    wire c4384;
    assign in4384_1 = {pp103[60]};
    assign in4384_2 = {pp104[59]};
    Full_Adder FA_4384(s4384, c4384, in4384_1, in4384_2, pp102[61]);
    wire[0:0] s4385, in4385_1, in4385_2;
    wire c4385;
    assign in4385_1 = {pp106[57]};
    assign in4385_2 = {pp107[56]};
    Full_Adder FA_4385(s4385, c4385, in4385_1, in4385_2, pp105[58]);
    wire[0:0] s4386, in4386_1, in4386_2;
    wire c4386;
    assign in4386_1 = {pp109[54]};
    assign in4386_2 = {pp110[53]};
    Full_Adder FA_4386(s4386, c4386, in4386_1, in4386_2, pp108[55]);
    wire[0:0] s4387, in4387_1, in4387_2;
    wire c4387;
    assign in4387_1 = {pp112[51]};
    assign in4387_2 = {pp113[50]};
    Full_Adder FA_4387(s4387, c4387, in4387_1, in4387_2, pp111[52]);
    wire[0:0] s4388, in4388_1, in4388_2;
    wire c4388;
    assign in4388_1 = {pp115[48]};
    assign in4388_2 = {pp116[47]};
    Full_Adder FA_4388(s4388, c4388, in4388_1, in4388_2, pp114[49]);
    wire[0:0] s4389, in4389_1, in4389_2;
    wire c4389;
    assign in4389_1 = {pp118[45]};
    assign in4389_2 = {pp119[44]};
    Full_Adder FA_4389(s4389, c4389, in4389_1, in4389_2, pp117[46]);
    wire[0:0] s4390, in4390_1, in4390_2;
    wire c4390;
    assign in4390_1 = {pp121[42]};
    assign in4390_2 = {pp122[41]};
    Full_Adder FA_4390(s4390, c4390, in4390_1, in4390_2, pp120[43]);
    wire[0:0] s4391, in4391_1, in4391_2;
    wire c4391;
    assign in4391_1 = {pp124[39]};
    assign in4391_2 = {pp125[38]};
    Full_Adder FA_4391(s4391, c4391, in4391_1, in4391_2, pp123[40]);
    wire[0:0] s4392, in4392_1, in4392_2;
    wire c4392;
    assign in4392_1 = {pp127[36]};
    assign in4392_2 = {c1771};
    Full_Adder FA_4392(s4392, c4392, in4392_1, in4392_2, pp126[37]);
    wire[0:0] s4393, in4393_1, in4393_2;
    wire c4393;
    assign in4393_1 = {c1773};
    assign in4393_2 = {c1774};
    Full_Adder FA_4393(s4393, c4393, in4393_1, in4393_2, c1772);
    wire[0:0] s4394, in4394_1, in4394_2;
    wire c4394;
    assign in4394_1 = {c1776};
    assign in4394_2 = {c1777};
    Full_Adder FA_4394(s4394, c4394, in4394_1, in4394_2, c1775);
    wire[0:0] s4395, in4395_1, in4395_2;
    wire c4395;
    assign in4395_1 = {s1779[0]};
    assign in4395_2 = {s1780[0]};
    Full_Adder FA_4395(s4395, c4395, in4395_1, in4395_2, c1778);
    wire[0:0] s4396, in4396_1, in4396_2;
    wire c4396;
    assign in4396_1 = {s1782[0]};
    assign in4396_2 = {s1783[0]};
    Full_Adder FA_4396(s4396, c4396, in4396_1, in4396_2, s1781[0]);
    wire[0:0] s4397, in4397_1, in4397_2;
    wire c4397;
    assign in4397_1 = {pp56[108]};
    assign in4397_2 = {pp57[107]};
    Full_Adder FA_4397(s4397, c4397, in4397_1, in4397_2, pp55[109]);
    wire[0:0] s4398, in4398_1, in4398_2;
    wire c4398;
    assign in4398_1 = {pp59[105]};
    assign in4398_2 = {pp60[104]};
    Full_Adder FA_4398(s4398, c4398, in4398_1, in4398_2, pp58[106]);
    wire[0:0] s4399, in4399_1, in4399_2;
    wire c4399;
    assign in4399_1 = {pp62[102]};
    assign in4399_2 = {pp63[101]};
    Full_Adder FA_4399(s4399, c4399, in4399_1, in4399_2, pp61[103]);
    wire[0:0] s4400, in4400_1, in4400_2;
    wire c4400;
    assign in4400_1 = {pp65[99]};
    assign in4400_2 = {pp66[98]};
    Full_Adder FA_4400(s4400, c4400, in4400_1, in4400_2, pp64[100]);
    wire[0:0] s4401, in4401_1, in4401_2;
    wire c4401;
    assign in4401_1 = {pp68[96]};
    assign in4401_2 = {pp69[95]};
    Full_Adder FA_4401(s4401, c4401, in4401_1, in4401_2, pp67[97]);
    wire[0:0] s4402, in4402_1, in4402_2;
    wire c4402;
    assign in4402_1 = {pp71[93]};
    assign in4402_2 = {pp72[92]};
    Full_Adder FA_4402(s4402, c4402, in4402_1, in4402_2, pp70[94]);
    wire[0:0] s4403, in4403_1, in4403_2;
    wire c4403;
    assign in4403_1 = {pp74[90]};
    assign in4403_2 = {pp75[89]};
    Full_Adder FA_4403(s4403, c4403, in4403_1, in4403_2, pp73[91]);
    wire[0:0] s4404, in4404_1, in4404_2;
    wire c4404;
    assign in4404_1 = {pp77[87]};
    assign in4404_2 = {pp78[86]};
    Full_Adder FA_4404(s4404, c4404, in4404_1, in4404_2, pp76[88]);
    wire[0:0] s4405, in4405_1, in4405_2;
    wire c4405;
    assign in4405_1 = {pp80[84]};
    assign in4405_2 = {pp81[83]};
    Full_Adder FA_4405(s4405, c4405, in4405_1, in4405_2, pp79[85]);
    wire[0:0] s4406, in4406_1, in4406_2;
    wire c4406;
    assign in4406_1 = {pp83[81]};
    assign in4406_2 = {pp84[80]};
    Full_Adder FA_4406(s4406, c4406, in4406_1, in4406_2, pp82[82]);
    wire[0:0] s4407, in4407_1, in4407_2;
    wire c4407;
    assign in4407_1 = {pp86[78]};
    assign in4407_2 = {pp87[77]};
    Full_Adder FA_4407(s4407, c4407, in4407_1, in4407_2, pp85[79]);
    wire[0:0] s4408, in4408_1, in4408_2;
    wire c4408;
    assign in4408_1 = {pp89[75]};
    assign in4408_2 = {pp90[74]};
    Full_Adder FA_4408(s4408, c4408, in4408_1, in4408_2, pp88[76]);
    wire[0:0] s4409, in4409_1, in4409_2;
    wire c4409;
    assign in4409_1 = {pp92[72]};
    assign in4409_2 = {pp93[71]};
    Full_Adder FA_4409(s4409, c4409, in4409_1, in4409_2, pp91[73]);
    wire[0:0] s4410, in4410_1, in4410_2;
    wire c4410;
    assign in4410_1 = {pp95[69]};
    assign in4410_2 = {pp96[68]};
    Full_Adder FA_4410(s4410, c4410, in4410_1, in4410_2, pp94[70]);
    wire[0:0] s4411, in4411_1, in4411_2;
    wire c4411;
    assign in4411_1 = {pp98[66]};
    assign in4411_2 = {pp99[65]};
    Full_Adder FA_4411(s4411, c4411, in4411_1, in4411_2, pp97[67]);
    wire[0:0] s4412, in4412_1, in4412_2;
    wire c4412;
    assign in4412_1 = {pp101[63]};
    assign in4412_2 = {pp102[62]};
    Full_Adder FA_4412(s4412, c4412, in4412_1, in4412_2, pp100[64]);
    wire[0:0] s4413, in4413_1, in4413_2;
    wire c4413;
    assign in4413_1 = {pp104[60]};
    assign in4413_2 = {pp105[59]};
    Full_Adder FA_4413(s4413, c4413, in4413_1, in4413_2, pp103[61]);
    wire[0:0] s4414, in4414_1, in4414_2;
    wire c4414;
    assign in4414_1 = {pp107[57]};
    assign in4414_2 = {pp108[56]};
    Full_Adder FA_4414(s4414, c4414, in4414_1, in4414_2, pp106[58]);
    wire[0:0] s4415, in4415_1, in4415_2;
    wire c4415;
    assign in4415_1 = {pp110[54]};
    assign in4415_2 = {pp111[53]};
    Full_Adder FA_4415(s4415, c4415, in4415_1, in4415_2, pp109[55]);
    wire[0:0] s4416, in4416_1, in4416_2;
    wire c4416;
    assign in4416_1 = {pp113[51]};
    assign in4416_2 = {pp114[50]};
    Full_Adder FA_4416(s4416, c4416, in4416_1, in4416_2, pp112[52]);
    wire[0:0] s4417, in4417_1, in4417_2;
    wire c4417;
    assign in4417_1 = {pp116[48]};
    assign in4417_2 = {pp117[47]};
    Full_Adder FA_4417(s4417, c4417, in4417_1, in4417_2, pp115[49]);
    wire[0:0] s4418, in4418_1, in4418_2;
    wire c4418;
    assign in4418_1 = {pp119[45]};
    assign in4418_2 = {pp120[44]};
    Full_Adder FA_4418(s4418, c4418, in4418_1, in4418_2, pp118[46]);
    wire[0:0] s4419, in4419_1, in4419_2;
    wire c4419;
    assign in4419_1 = {pp122[42]};
    assign in4419_2 = {pp123[41]};
    Full_Adder FA_4419(s4419, c4419, in4419_1, in4419_2, pp121[43]);
    wire[0:0] s4420, in4420_1, in4420_2;
    wire c4420;
    assign in4420_1 = {pp125[39]};
    assign in4420_2 = {pp126[38]};
    Full_Adder FA_4420(s4420, c4420, in4420_1, in4420_2, pp124[40]);
    wire[0:0] s4421, in4421_1, in4421_2;
    wire c4421;
    assign in4421_1 = {c1779};
    assign in4421_2 = {c1780};
    Full_Adder FA_4421(s4421, c4421, in4421_1, in4421_2, pp127[37]);
    wire[0:0] s4422, in4422_1, in4422_2;
    wire c4422;
    assign in4422_1 = {c1782};
    assign in4422_2 = {c1783};
    Full_Adder FA_4422(s4422, c4422, in4422_1, in4422_2, c1781);
    wire[0:0] s4423, in4423_1, in4423_2;
    wire c4423;
    assign in4423_1 = {c1785};
    assign in4423_2 = {s1786[0]};
    Full_Adder FA_4423(s4423, c4423, in4423_1, in4423_2, c1784);
    wire[0:0] s4424, in4424_1, in4424_2;
    wire c4424;
    assign in4424_1 = {s1788[0]};
    assign in4424_2 = {s1789[0]};
    Full_Adder FA_4424(s4424, c4424, in4424_1, in4424_2, s1787[0]);
    wire[0:0] s4425, in4425_1, in4425_2;
    wire c4425;
    assign in4425_1 = {pp54[111]};
    assign in4425_2 = {pp55[110]};
    Full_Adder FA_4425(s4425, c4425, in4425_1, in4425_2, pp53[112]);
    wire[0:0] s4426, in4426_1, in4426_2;
    wire c4426;
    assign in4426_1 = {pp57[108]};
    assign in4426_2 = {pp58[107]};
    Full_Adder FA_4426(s4426, c4426, in4426_1, in4426_2, pp56[109]);
    wire[0:0] s4427, in4427_1, in4427_2;
    wire c4427;
    assign in4427_1 = {pp60[105]};
    assign in4427_2 = {pp61[104]};
    Full_Adder FA_4427(s4427, c4427, in4427_1, in4427_2, pp59[106]);
    wire[0:0] s4428, in4428_1, in4428_2;
    wire c4428;
    assign in4428_1 = {pp63[102]};
    assign in4428_2 = {pp64[101]};
    Full_Adder FA_4428(s4428, c4428, in4428_1, in4428_2, pp62[103]);
    wire[0:0] s4429, in4429_1, in4429_2;
    wire c4429;
    assign in4429_1 = {pp66[99]};
    assign in4429_2 = {pp67[98]};
    Full_Adder FA_4429(s4429, c4429, in4429_1, in4429_2, pp65[100]);
    wire[0:0] s4430, in4430_1, in4430_2;
    wire c4430;
    assign in4430_1 = {pp69[96]};
    assign in4430_2 = {pp70[95]};
    Full_Adder FA_4430(s4430, c4430, in4430_1, in4430_2, pp68[97]);
    wire[0:0] s4431, in4431_1, in4431_2;
    wire c4431;
    assign in4431_1 = {pp72[93]};
    assign in4431_2 = {pp73[92]};
    Full_Adder FA_4431(s4431, c4431, in4431_1, in4431_2, pp71[94]);
    wire[0:0] s4432, in4432_1, in4432_2;
    wire c4432;
    assign in4432_1 = {pp75[90]};
    assign in4432_2 = {pp76[89]};
    Full_Adder FA_4432(s4432, c4432, in4432_1, in4432_2, pp74[91]);
    wire[0:0] s4433, in4433_1, in4433_2;
    wire c4433;
    assign in4433_1 = {pp78[87]};
    assign in4433_2 = {pp79[86]};
    Full_Adder FA_4433(s4433, c4433, in4433_1, in4433_2, pp77[88]);
    wire[0:0] s4434, in4434_1, in4434_2;
    wire c4434;
    assign in4434_1 = {pp81[84]};
    assign in4434_2 = {pp82[83]};
    Full_Adder FA_4434(s4434, c4434, in4434_1, in4434_2, pp80[85]);
    wire[0:0] s4435, in4435_1, in4435_2;
    wire c4435;
    assign in4435_1 = {pp84[81]};
    assign in4435_2 = {pp85[80]};
    Full_Adder FA_4435(s4435, c4435, in4435_1, in4435_2, pp83[82]);
    wire[0:0] s4436, in4436_1, in4436_2;
    wire c4436;
    assign in4436_1 = {pp87[78]};
    assign in4436_2 = {pp88[77]};
    Full_Adder FA_4436(s4436, c4436, in4436_1, in4436_2, pp86[79]);
    wire[0:0] s4437, in4437_1, in4437_2;
    wire c4437;
    assign in4437_1 = {pp90[75]};
    assign in4437_2 = {pp91[74]};
    Full_Adder FA_4437(s4437, c4437, in4437_1, in4437_2, pp89[76]);
    wire[0:0] s4438, in4438_1, in4438_2;
    wire c4438;
    assign in4438_1 = {pp93[72]};
    assign in4438_2 = {pp94[71]};
    Full_Adder FA_4438(s4438, c4438, in4438_1, in4438_2, pp92[73]);
    wire[0:0] s4439, in4439_1, in4439_2;
    wire c4439;
    assign in4439_1 = {pp96[69]};
    assign in4439_2 = {pp97[68]};
    Full_Adder FA_4439(s4439, c4439, in4439_1, in4439_2, pp95[70]);
    wire[0:0] s4440, in4440_1, in4440_2;
    wire c4440;
    assign in4440_1 = {pp99[66]};
    assign in4440_2 = {pp100[65]};
    Full_Adder FA_4440(s4440, c4440, in4440_1, in4440_2, pp98[67]);
    wire[0:0] s4441, in4441_1, in4441_2;
    wire c4441;
    assign in4441_1 = {pp102[63]};
    assign in4441_2 = {pp103[62]};
    Full_Adder FA_4441(s4441, c4441, in4441_1, in4441_2, pp101[64]);
    wire[0:0] s4442, in4442_1, in4442_2;
    wire c4442;
    assign in4442_1 = {pp105[60]};
    assign in4442_2 = {pp106[59]};
    Full_Adder FA_4442(s4442, c4442, in4442_1, in4442_2, pp104[61]);
    wire[0:0] s4443, in4443_1, in4443_2;
    wire c4443;
    assign in4443_1 = {pp108[57]};
    assign in4443_2 = {pp109[56]};
    Full_Adder FA_4443(s4443, c4443, in4443_1, in4443_2, pp107[58]);
    wire[0:0] s4444, in4444_1, in4444_2;
    wire c4444;
    assign in4444_1 = {pp111[54]};
    assign in4444_2 = {pp112[53]};
    Full_Adder FA_4444(s4444, c4444, in4444_1, in4444_2, pp110[55]);
    wire[0:0] s4445, in4445_1, in4445_2;
    wire c4445;
    assign in4445_1 = {pp114[51]};
    assign in4445_2 = {pp115[50]};
    Full_Adder FA_4445(s4445, c4445, in4445_1, in4445_2, pp113[52]);
    wire[0:0] s4446, in4446_1, in4446_2;
    wire c4446;
    assign in4446_1 = {pp117[48]};
    assign in4446_2 = {pp118[47]};
    Full_Adder FA_4446(s4446, c4446, in4446_1, in4446_2, pp116[49]);
    wire[0:0] s4447, in4447_1, in4447_2;
    wire c4447;
    assign in4447_1 = {pp120[45]};
    assign in4447_2 = {pp121[44]};
    Full_Adder FA_4447(s4447, c4447, in4447_1, in4447_2, pp119[46]);
    wire[0:0] s4448, in4448_1, in4448_2;
    wire c4448;
    assign in4448_1 = {pp123[42]};
    assign in4448_2 = {pp124[41]};
    Full_Adder FA_4448(s4448, c4448, in4448_1, in4448_2, pp122[43]);
    wire[0:0] s4449, in4449_1, in4449_2;
    wire c4449;
    assign in4449_1 = {pp126[39]};
    assign in4449_2 = {pp127[38]};
    Full_Adder FA_4449(s4449, c4449, in4449_1, in4449_2, pp125[40]);
    wire[0:0] s4450, in4450_1, in4450_2;
    wire c4450;
    assign in4450_1 = {c1787};
    assign in4450_2 = {c1788};
    Full_Adder FA_4450(s4450, c4450, in4450_1, in4450_2, c1786);
    wire[0:0] s4451, in4451_1, in4451_2;
    wire c4451;
    assign in4451_1 = {c1790};
    assign in4451_2 = {c1791};
    Full_Adder FA_4451(s4451, c4451, in4451_1, in4451_2, c1789);
    wire[0:0] s4452, in4452_1, in4452_2;
    wire c4452;
    assign in4452_1 = {s1793[0]};
    assign in4452_2 = {s1794[0]};
    Full_Adder FA_4452(s4452, c4452, in4452_1, in4452_2, s1792[0]);
    wire[0:0] s4453, in4453_1, in4453_2;
    wire c4453;
    assign in4453_1 = {pp52[114]};
    assign in4453_2 = {pp53[113]};
    Full_Adder FA_4453(s4453, c4453, in4453_1, in4453_2, pp51[115]);
    wire[0:0] s4454, in4454_1, in4454_2;
    wire c4454;
    assign in4454_1 = {pp55[111]};
    assign in4454_2 = {pp56[110]};
    Full_Adder FA_4454(s4454, c4454, in4454_1, in4454_2, pp54[112]);
    wire[0:0] s4455, in4455_1, in4455_2;
    wire c4455;
    assign in4455_1 = {pp58[108]};
    assign in4455_2 = {pp59[107]};
    Full_Adder FA_4455(s4455, c4455, in4455_1, in4455_2, pp57[109]);
    wire[0:0] s4456, in4456_1, in4456_2;
    wire c4456;
    assign in4456_1 = {pp61[105]};
    assign in4456_2 = {pp62[104]};
    Full_Adder FA_4456(s4456, c4456, in4456_1, in4456_2, pp60[106]);
    wire[0:0] s4457, in4457_1, in4457_2;
    wire c4457;
    assign in4457_1 = {pp64[102]};
    assign in4457_2 = {pp65[101]};
    Full_Adder FA_4457(s4457, c4457, in4457_1, in4457_2, pp63[103]);
    wire[0:0] s4458, in4458_1, in4458_2;
    wire c4458;
    assign in4458_1 = {pp67[99]};
    assign in4458_2 = {pp68[98]};
    Full_Adder FA_4458(s4458, c4458, in4458_1, in4458_2, pp66[100]);
    wire[0:0] s4459, in4459_1, in4459_2;
    wire c4459;
    assign in4459_1 = {pp70[96]};
    assign in4459_2 = {pp71[95]};
    Full_Adder FA_4459(s4459, c4459, in4459_1, in4459_2, pp69[97]);
    wire[0:0] s4460, in4460_1, in4460_2;
    wire c4460;
    assign in4460_1 = {pp73[93]};
    assign in4460_2 = {pp74[92]};
    Full_Adder FA_4460(s4460, c4460, in4460_1, in4460_2, pp72[94]);
    wire[0:0] s4461, in4461_1, in4461_2;
    wire c4461;
    assign in4461_1 = {pp76[90]};
    assign in4461_2 = {pp77[89]};
    Full_Adder FA_4461(s4461, c4461, in4461_1, in4461_2, pp75[91]);
    wire[0:0] s4462, in4462_1, in4462_2;
    wire c4462;
    assign in4462_1 = {pp79[87]};
    assign in4462_2 = {pp80[86]};
    Full_Adder FA_4462(s4462, c4462, in4462_1, in4462_2, pp78[88]);
    wire[0:0] s4463, in4463_1, in4463_2;
    wire c4463;
    assign in4463_1 = {pp82[84]};
    assign in4463_2 = {pp83[83]};
    Full_Adder FA_4463(s4463, c4463, in4463_1, in4463_2, pp81[85]);
    wire[0:0] s4464, in4464_1, in4464_2;
    wire c4464;
    assign in4464_1 = {pp85[81]};
    assign in4464_2 = {pp86[80]};
    Full_Adder FA_4464(s4464, c4464, in4464_1, in4464_2, pp84[82]);
    wire[0:0] s4465, in4465_1, in4465_2;
    wire c4465;
    assign in4465_1 = {pp88[78]};
    assign in4465_2 = {pp89[77]};
    Full_Adder FA_4465(s4465, c4465, in4465_1, in4465_2, pp87[79]);
    wire[0:0] s4466, in4466_1, in4466_2;
    wire c4466;
    assign in4466_1 = {pp91[75]};
    assign in4466_2 = {pp92[74]};
    Full_Adder FA_4466(s4466, c4466, in4466_1, in4466_2, pp90[76]);
    wire[0:0] s4467, in4467_1, in4467_2;
    wire c4467;
    assign in4467_1 = {pp94[72]};
    assign in4467_2 = {pp95[71]};
    Full_Adder FA_4467(s4467, c4467, in4467_1, in4467_2, pp93[73]);
    wire[0:0] s4468, in4468_1, in4468_2;
    wire c4468;
    assign in4468_1 = {pp97[69]};
    assign in4468_2 = {pp98[68]};
    Full_Adder FA_4468(s4468, c4468, in4468_1, in4468_2, pp96[70]);
    wire[0:0] s4469, in4469_1, in4469_2;
    wire c4469;
    assign in4469_1 = {pp100[66]};
    assign in4469_2 = {pp101[65]};
    Full_Adder FA_4469(s4469, c4469, in4469_1, in4469_2, pp99[67]);
    wire[0:0] s4470, in4470_1, in4470_2;
    wire c4470;
    assign in4470_1 = {pp103[63]};
    assign in4470_2 = {pp104[62]};
    Full_Adder FA_4470(s4470, c4470, in4470_1, in4470_2, pp102[64]);
    wire[0:0] s4471, in4471_1, in4471_2;
    wire c4471;
    assign in4471_1 = {pp106[60]};
    assign in4471_2 = {pp107[59]};
    Full_Adder FA_4471(s4471, c4471, in4471_1, in4471_2, pp105[61]);
    wire[0:0] s4472, in4472_1, in4472_2;
    wire c4472;
    assign in4472_1 = {pp109[57]};
    assign in4472_2 = {pp110[56]};
    Full_Adder FA_4472(s4472, c4472, in4472_1, in4472_2, pp108[58]);
    wire[0:0] s4473, in4473_1, in4473_2;
    wire c4473;
    assign in4473_1 = {pp112[54]};
    assign in4473_2 = {pp113[53]};
    Full_Adder FA_4473(s4473, c4473, in4473_1, in4473_2, pp111[55]);
    wire[0:0] s4474, in4474_1, in4474_2;
    wire c4474;
    assign in4474_1 = {pp115[51]};
    assign in4474_2 = {pp116[50]};
    Full_Adder FA_4474(s4474, c4474, in4474_1, in4474_2, pp114[52]);
    wire[0:0] s4475, in4475_1, in4475_2;
    wire c4475;
    assign in4475_1 = {pp118[48]};
    assign in4475_2 = {pp119[47]};
    Full_Adder FA_4475(s4475, c4475, in4475_1, in4475_2, pp117[49]);
    wire[0:0] s4476, in4476_1, in4476_2;
    wire c4476;
    assign in4476_1 = {pp121[45]};
    assign in4476_2 = {pp122[44]};
    Full_Adder FA_4476(s4476, c4476, in4476_1, in4476_2, pp120[46]);
    wire[0:0] s4477, in4477_1, in4477_2;
    wire c4477;
    assign in4477_1 = {pp124[42]};
    assign in4477_2 = {pp125[41]};
    Full_Adder FA_4477(s4477, c4477, in4477_1, in4477_2, pp123[43]);
    wire[0:0] s4478, in4478_1, in4478_2;
    wire c4478;
    assign in4478_1 = {pp127[39]};
    assign in4478_2 = {c1792};
    Full_Adder FA_4478(s4478, c4478, in4478_1, in4478_2, pp126[40]);
    wire[0:0] s4479, in4479_1, in4479_2;
    wire c4479;
    assign in4479_1 = {c1794};
    assign in4479_2 = {c1795};
    Full_Adder FA_4479(s4479, c4479, in4479_1, in4479_2, c1793);
    wire[0:0] s4480, in4480_1, in4480_2;
    wire c4480;
    assign in4480_1 = {s1797[0]};
    assign in4480_2 = {s1798[0]};
    Full_Adder FA_4480(s4480, c4480, in4480_1, in4480_2, c1796);
    wire[0:0] s4481, in4481_1, in4481_2;
    wire c4481;
    assign in4481_1 = {pp50[117]};
    assign in4481_2 = {pp51[116]};
    Full_Adder FA_4481(s4481, c4481, in4481_1, in4481_2, pp49[118]);
    wire[0:0] s4482, in4482_1, in4482_2;
    wire c4482;
    assign in4482_1 = {pp53[114]};
    assign in4482_2 = {pp54[113]};
    Full_Adder FA_4482(s4482, c4482, in4482_1, in4482_2, pp52[115]);
    wire[0:0] s4483, in4483_1, in4483_2;
    wire c4483;
    assign in4483_1 = {pp56[111]};
    assign in4483_2 = {pp57[110]};
    Full_Adder FA_4483(s4483, c4483, in4483_1, in4483_2, pp55[112]);
    wire[0:0] s4484, in4484_1, in4484_2;
    wire c4484;
    assign in4484_1 = {pp59[108]};
    assign in4484_2 = {pp60[107]};
    Full_Adder FA_4484(s4484, c4484, in4484_1, in4484_2, pp58[109]);
    wire[0:0] s4485, in4485_1, in4485_2;
    wire c4485;
    assign in4485_1 = {pp62[105]};
    assign in4485_2 = {pp63[104]};
    Full_Adder FA_4485(s4485, c4485, in4485_1, in4485_2, pp61[106]);
    wire[0:0] s4486, in4486_1, in4486_2;
    wire c4486;
    assign in4486_1 = {pp65[102]};
    assign in4486_2 = {pp66[101]};
    Full_Adder FA_4486(s4486, c4486, in4486_1, in4486_2, pp64[103]);
    wire[0:0] s4487, in4487_1, in4487_2;
    wire c4487;
    assign in4487_1 = {pp68[99]};
    assign in4487_2 = {pp69[98]};
    Full_Adder FA_4487(s4487, c4487, in4487_1, in4487_2, pp67[100]);
    wire[0:0] s4488, in4488_1, in4488_2;
    wire c4488;
    assign in4488_1 = {pp71[96]};
    assign in4488_2 = {pp72[95]};
    Full_Adder FA_4488(s4488, c4488, in4488_1, in4488_2, pp70[97]);
    wire[0:0] s4489, in4489_1, in4489_2;
    wire c4489;
    assign in4489_1 = {pp74[93]};
    assign in4489_2 = {pp75[92]};
    Full_Adder FA_4489(s4489, c4489, in4489_1, in4489_2, pp73[94]);
    wire[0:0] s4490, in4490_1, in4490_2;
    wire c4490;
    assign in4490_1 = {pp77[90]};
    assign in4490_2 = {pp78[89]};
    Full_Adder FA_4490(s4490, c4490, in4490_1, in4490_2, pp76[91]);
    wire[0:0] s4491, in4491_1, in4491_2;
    wire c4491;
    assign in4491_1 = {pp80[87]};
    assign in4491_2 = {pp81[86]};
    Full_Adder FA_4491(s4491, c4491, in4491_1, in4491_2, pp79[88]);
    wire[0:0] s4492, in4492_1, in4492_2;
    wire c4492;
    assign in4492_1 = {pp83[84]};
    assign in4492_2 = {pp84[83]};
    Full_Adder FA_4492(s4492, c4492, in4492_1, in4492_2, pp82[85]);
    wire[0:0] s4493, in4493_1, in4493_2;
    wire c4493;
    assign in4493_1 = {pp86[81]};
    assign in4493_2 = {pp87[80]};
    Full_Adder FA_4493(s4493, c4493, in4493_1, in4493_2, pp85[82]);
    wire[0:0] s4494, in4494_1, in4494_2;
    wire c4494;
    assign in4494_1 = {pp89[78]};
    assign in4494_2 = {pp90[77]};
    Full_Adder FA_4494(s4494, c4494, in4494_1, in4494_2, pp88[79]);
    wire[0:0] s4495, in4495_1, in4495_2;
    wire c4495;
    assign in4495_1 = {pp92[75]};
    assign in4495_2 = {pp93[74]};
    Full_Adder FA_4495(s4495, c4495, in4495_1, in4495_2, pp91[76]);
    wire[0:0] s4496, in4496_1, in4496_2;
    wire c4496;
    assign in4496_1 = {pp95[72]};
    assign in4496_2 = {pp96[71]};
    Full_Adder FA_4496(s4496, c4496, in4496_1, in4496_2, pp94[73]);
    wire[0:0] s4497, in4497_1, in4497_2;
    wire c4497;
    assign in4497_1 = {pp98[69]};
    assign in4497_2 = {pp99[68]};
    Full_Adder FA_4497(s4497, c4497, in4497_1, in4497_2, pp97[70]);
    wire[0:0] s4498, in4498_1, in4498_2;
    wire c4498;
    assign in4498_1 = {pp101[66]};
    assign in4498_2 = {pp102[65]};
    Full_Adder FA_4498(s4498, c4498, in4498_1, in4498_2, pp100[67]);
    wire[0:0] s4499, in4499_1, in4499_2;
    wire c4499;
    assign in4499_1 = {pp104[63]};
    assign in4499_2 = {pp105[62]};
    Full_Adder FA_4499(s4499, c4499, in4499_1, in4499_2, pp103[64]);
    wire[0:0] s4500, in4500_1, in4500_2;
    wire c4500;
    assign in4500_1 = {pp107[60]};
    assign in4500_2 = {pp108[59]};
    Full_Adder FA_4500(s4500, c4500, in4500_1, in4500_2, pp106[61]);
    wire[0:0] s4501, in4501_1, in4501_2;
    wire c4501;
    assign in4501_1 = {pp110[57]};
    assign in4501_2 = {pp111[56]};
    Full_Adder FA_4501(s4501, c4501, in4501_1, in4501_2, pp109[58]);
    wire[0:0] s4502, in4502_1, in4502_2;
    wire c4502;
    assign in4502_1 = {pp113[54]};
    assign in4502_2 = {pp114[53]};
    Full_Adder FA_4502(s4502, c4502, in4502_1, in4502_2, pp112[55]);
    wire[0:0] s4503, in4503_1, in4503_2;
    wire c4503;
    assign in4503_1 = {pp116[51]};
    assign in4503_2 = {pp117[50]};
    Full_Adder FA_4503(s4503, c4503, in4503_1, in4503_2, pp115[52]);
    wire[0:0] s4504, in4504_1, in4504_2;
    wire c4504;
    assign in4504_1 = {pp119[48]};
    assign in4504_2 = {pp120[47]};
    Full_Adder FA_4504(s4504, c4504, in4504_1, in4504_2, pp118[49]);
    wire[0:0] s4505, in4505_1, in4505_2;
    wire c4505;
    assign in4505_1 = {pp122[45]};
    assign in4505_2 = {pp123[44]};
    Full_Adder FA_4505(s4505, c4505, in4505_1, in4505_2, pp121[46]);
    wire[0:0] s4506, in4506_1, in4506_2;
    wire c4506;
    assign in4506_1 = {pp125[42]};
    assign in4506_2 = {pp126[41]};
    Full_Adder FA_4506(s4506, c4506, in4506_1, in4506_2, pp124[43]);
    wire[0:0] s4507, in4507_1, in4507_2;
    wire c4507;
    assign in4507_1 = {c1797};
    assign in4507_2 = {c1798};
    Full_Adder FA_4507(s4507, c4507, in4507_1, in4507_2, pp127[40]);
    wire[0:0] s4508, in4508_1, in4508_2;
    wire c4508;
    assign in4508_1 = {c1800};
    assign in4508_2 = {s1801[0]};
    Full_Adder FA_4508(s4508, c4508, in4508_1, in4508_2, c1799);
    wire[0:0] s4509, in4509_1, in4509_2;
    wire c4509;
    assign in4509_1 = {pp48[120]};
    assign in4509_2 = {pp49[119]};
    Full_Adder FA_4509(s4509, c4509, in4509_1, in4509_2, pp47[121]);
    wire[0:0] s4510, in4510_1, in4510_2;
    wire c4510;
    assign in4510_1 = {pp51[117]};
    assign in4510_2 = {pp52[116]};
    Full_Adder FA_4510(s4510, c4510, in4510_1, in4510_2, pp50[118]);
    wire[0:0] s4511, in4511_1, in4511_2;
    wire c4511;
    assign in4511_1 = {pp54[114]};
    assign in4511_2 = {pp55[113]};
    Full_Adder FA_4511(s4511, c4511, in4511_1, in4511_2, pp53[115]);
    wire[0:0] s4512, in4512_1, in4512_2;
    wire c4512;
    assign in4512_1 = {pp57[111]};
    assign in4512_2 = {pp58[110]};
    Full_Adder FA_4512(s4512, c4512, in4512_1, in4512_2, pp56[112]);
    wire[0:0] s4513, in4513_1, in4513_2;
    wire c4513;
    assign in4513_1 = {pp60[108]};
    assign in4513_2 = {pp61[107]};
    Full_Adder FA_4513(s4513, c4513, in4513_1, in4513_2, pp59[109]);
    wire[0:0] s4514, in4514_1, in4514_2;
    wire c4514;
    assign in4514_1 = {pp63[105]};
    assign in4514_2 = {pp64[104]};
    Full_Adder FA_4514(s4514, c4514, in4514_1, in4514_2, pp62[106]);
    wire[0:0] s4515, in4515_1, in4515_2;
    wire c4515;
    assign in4515_1 = {pp66[102]};
    assign in4515_2 = {pp67[101]};
    Full_Adder FA_4515(s4515, c4515, in4515_1, in4515_2, pp65[103]);
    wire[0:0] s4516, in4516_1, in4516_2;
    wire c4516;
    assign in4516_1 = {pp69[99]};
    assign in4516_2 = {pp70[98]};
    Full_Adder FA_4516(s4516, c4516, in4516_1, in4516_2, pp68[100]);
    wire[0:0] s4517, in4517_1, in4517_2;
    wire c4517;
    assign in4517_1 = {pp72[96]};
    assign in4517_2 = {pp73[95]};
    Full_Adder FA_4517(s4517, c4517, in4517_1, in4517_2, pp71[97]);
    wire[0:0] s4518, in4518_1, in4518_2;
    wire c4518;
    assign in4518_1 = {pp75[93]};
    assign in4518_2 = {pp76[92]};
    Full_Adder FA_4518(s4518, c4518, in4518_1, in4518_2, pp74[94]);
    wire[0:0] s4519, in4519_1, in4519_2;
    wire c4519;
    assign in4519_1 = {pp78[90]};
    assign in4519_2 = {pp79[89]};
    Full_Adder FA_4519(s4519, c4519, in4519_1, in4519_2, pp77[91]);
    wire[0:0] s4520, in4520_1, in4520_2;
    wire c4520;
    assign in4520_1 = {pp81[87]};
    assign in4520_2 = {pp82[86]};
    Full_Adder FA_4520(s4520, c4520, in4520_1, in4520_2, pp80[88]);
    wire[0:0] s4521, in4521_1, in4521_2;
    wire c4521;
    assign in4521_1 = {pp84[84]};
    assign in4521_2 = {pp85[83]};
    Full_Adder FA_4521(s4521, c4521, in4521_1, in4521_2, pp83[85]);
    wire[0:0] s4522, in4522_1, in4522_2;
    wire c4522;
    assign in4522_1 = {pp87[81]};
    assign in4522_2 = {pp88[80]};
    Full_Adder FA_4522(s4522, c4522, in4522_1, in4522_2, pp86[82]);
    wire[0:0] s4523, in4523_1, in4523_2;
    wire c4523;
    assign in4523_1 = {pp90[78]};
    assign in4523_2 = {pp91[77]};
    Full_Adder FA_4523(s4523, c4523, in4523_1, in4523_2, pp89[79]);
    wire[0:0] s4524, in4524_1, in4524_2;
    wire c4524;
    assign in4524_1 = {pp93[75]};
    assign in4524_2 = {pp94[74]};
    Full_Adder FA_4524(s4524, c4524, in4524_1, in4524_2, pp92[76]);
    wire[0:0] s4525, in4525_1, in4525_2;
    wire c4525;
    assign in4525_1 = {pp96[72]};
    assign in4525_2 = {pp97[71]};
    Full_Adder FA_4525(s4525, c4525, in4525_1, in4525_2, pp95[73]);
    wire[0:0] s4526, in4526_1, in4526_2;
    wire c4526;
    assign in4526_1 = {pp99[69]};
    assign in4526_2 = {pp100[68]};
    Full_Adder FA_4526(s4526, c4526, in4526_1, in4526_2, pp98[70]);
    wire[0:0] s4527, in4527_1, in4527_2;
    wire c4527;
    assign in4527_1 = {pp102[66]};
    assign in4527_2 = {pp103[65]};
    Full_Adder FA_4527(s4527, c4527, in4527_1, in4527_2, pp101[67]);
    wire[0:0] s4528, in4528_1, in4528_2;
    wire c4528;
    assign in4528_1 = {pp105[63]};
    assign in4528_2 = {pp106[62]};
    Full_Adder FA_4528(s4528, c4528, in4528_1, in4528_2, pp104[64]);
    wire[0:0] s4529, in4529_1, in4529_2;
    wire c4529;
    assign in4529_1 = {pp108[60]};
    assign in4529_2 = {pp109[59]};
    Full_Adder FA_4529(s4529, c4529, in4529_1, in4529_2, pp107[61]);
    wire[0:0] s4530, in4530_1, in4530_2;
    wire c4530;
    assign in4530_1 = {pp111[57]};
    assign in4530_2 = {pp112[56]};
    Full_Adder FA_4530(s4530, c4530, in4530_1, in4530_2, pp110[58]);
    wire[0:0] s4531, in4531_1, in4531_2;
    wire c4531;
    assign in4531_1 = {pp114[54]};
    assign in4531_2 = {pp115[53]};
    Full_Adder FA_4531(s4531, c4531, in4531_1, in4531_2, pp113[55]);
    wire[0:0] s4532, in4532_1, in4532_2;
    wire c4532;
    assign in4532_1 = {pp117[51]};
    assign in4532_2 = {pp118[50]};
    Full_Adder FA_4532(s4532, c4532, in4532_1, in4532_2, pp116[52]);
    wire[0:0] s4533, in4533_1, in4533_2;
    wire c4533;
    assign in4533_1 = {pp120[48]};
    assign in4533_2 = {pp121[47]};
    Full_Adder FA_4533(s4533, c4533, in4533_1, in4533_2, pp119[49]);
    wire[0:0] s4534, in4534_1, in4534_2;
    wire c4534;
    assign in4534_1 = {pp123[45]};
    assign in4534_2 = {pp124[44]};
    Full_Adder FA_4534(s4534, c4534, in4534_1, in4534_2, pp122[46]);
    wire[0:0] s4535, in4535_1, in4535_2;
    wire c4535;
    assign in4535_1 = {pp126[42]};
    assign in4535_2 = {pp127[41]};
    Full_Adder FA_4535(s4535, c4535, in4535_1, in4535_2, pp125[43]);
    wire[0:0] s4536, in4536_1, in4536_2;
    wire c4536;
    assign in4536_1 = {c1802};
    assign in4536_2 = {c1803};
    Full_Adder FA_4536(s4536, c4536, in4536_1, in4536_2, c1801);
    wire[0:0] s4537, in4537_1, in4537_2;
    wire c4537;
    assign in4537_1 = {pp46[123]};
    assign in4537_2 = {pp47[122]};
    Full_Adder FA_4537(s4537, c4537, in4537_1, in4537_2, pp45[124]);
    wire[0:0] s4538, in4538_1, in4538_2;
    wire c4538;
    assign in4538_1 = {pp49[120]};
    assign in4538_2 = {pp50[119]};
    Full_Adder FA_4538(s4538, c4538, in4538_1, in4538_2, pp48[121]);
    wire[0:0] s4539, in4539_1, in4539_2;
    wire c4539;
    assign in4539_1 = {pp52[117]};
    assign in4539_2 = {pp53[116]};
    Full_Adder FA_4539(s4539, c4539, in4539_1, in4539_2, pp51[118]);
    wire[0:0] s4540, in4540_1, in4540_2;
    wire c4540;
    assign in4540_1 = {pp55[114]};
    assign in4540_2 = {pp56[113]};
    Full_Adder FA_4540(s4540, c4540, in4540_1, in4540_2, pp54[115]);
    wire[0:0] s4541, in4541_1, in4541_2;
    wire c4541;
    assign in4541_1 = {pp58[111]};
    assign in4541_2 = {pp59[110]};
    Full_Adder FA_4541(s4541, c4541, in4541_1, in4541_2, pp57[112]);
    wire[0:0] s4542, in4542_1, in4542_2;
    wire c4542;
    assign in4542_1 = {pp61[108]};
    assign in4542_2 = {pp62[107]};
    Full_Adder FA_4542(s4542, c4542, in4542_1, in4542_2, pp60[109]);
    wire[0:0] s4543, in4543_1, in4543_2;
    wire c4543;
    assign in4543_1 = {pp64[105]};
    assign in4543_2 = {pp65[104]};
    Full_Adder FA_4543(s4543, c4543, in4543_1, in4543_2, pp63[106]);
    wire[0:0] s4544, in4544_1, in4544_2;
    wire c4544;
    assign in4544_1 = {pp67[102]};
    assign in4544_2 = {pp68[101]};
    Full_Adder FA_4544(s4544, c4544, in4544_1, in4544_2, pp66[103]);
    wire[0:0] s4545, in4545_1, in4545_2;
    wire c4545;
    assign in4545_1 = {pp70[99]};
    assign in4545_2 = {pp71[98]};
    Full_Adder FA_4545(s4545, c4545, in4545_1, in4545_2, pp69[100]);
    wire[0:0] s4546, in4546_1, in4546_2;
    wire c4546;
    assign in4546_1 = {pp73[96]};
    assign in4546_2 = {pp74[95]};
    Full_Adder FA_4546(s4546, c4546, in4546_1, in4546_2, pp72[97]);
    wire[0:0] s4547, in4547_1, in4547_2;
    wire c4547;
    assign in4547_1 = {pp76[93]};
    assign in4547_2 = {pp77[92]};
    Full_Adder FA_4547(s4547, c4547, in4547_1, in4547_2, pp75[94]);
    wire[0:0] s4548, in4548_1, in4548_2;
    wire c4548;
    assign in4548_1 = {pp79[90]};
    assign in4548_2 = {pp80[89]};
    Full_Adder FA_4548(s4548, c4548, in4548_1, in4548_2, pp78[91]);
    wire[0:0] s4549, in4549_1, in4549_2;
    wire c4549;
    assign in4549_1 = {pp82[87]};
    assign in4549_2 = {pp83[86]};
    Full_Adder FA_4549(s4549, c4549, in4549_1, in4549_2, pp81[88]);
    wire[0:0] s4550, in4550_1, in4550_2;
    wire c4550;
    assign in4550_1 = {pp85[84]};
    assign in4550_2 = {pp86[83]};
    Full_Adder FA_4550(s4550, c4550, in4550_1, in4550_2, pp84[85]);
    wire[0:0] s4551, in4551_1, in4551_2;
    wire c4551;
    assign in4551_1 = {pp88[81]};
    assign in4551_2 = {pp89[80]};
    Full_Adder FA_4551(s4551, c4551, in4551_1, in4551_2, pp87[82]);
    wire[0:0] s4552, in4552_1, in4552_2;
    wire c4552;
    assign in4552_1 = {pp91[78]};
    assign in4552_2 = {pp92[77]};
    Full_Adder FA_4552(s4552, c4552, in4552_1, in4552_2, pp90[79]);
    wire[0:0] s4553, in4553_1, in4553_2;
    wire c4553;
    assign in4553_1 = {pp94[75]};
    assign in4553_2 = {pp95[74]};
    Full_Adder FA_4553(s4553, c4553, in4553_1, in4553_2, pp93[76]);
    wire[0:0] s4554, in4554_1, in4554_2;
    wire c4554;
    assign in4554_1 = {pp97[72]};
    assign in4554_2 = {pp98[71]};
    Full_Adder FA_4554(s4554, c4554, in4554_1, in4554_2, pp96[73]);
    wire[0:0] s4555, in4555_1, in4555_2;
    wire c4555;
    assign in4555_1 = {pp100[69]};
    assign in4555_2 = {pp101[68]};
    Full_Adder FA_4555(s4555, c4555, in4555_1, in4555_2, pp99[70]);
    wire[0:0] s4556, in4556_1, in4556_2;
    wire c4556;
    assign in4556_1 = {pp103[66]};
    assign in4556_2 = {pp104[65]};
    Full_Adder FA_4556(s4556, c4556, in4556_1, in4556_2, pp102[67]);
    wire[0:0] s4557, in4557_1, in4557_2;
    wire c4557;
    assign in4557_1 = {pp106[63]};
    assign in4557_2 = {pp107[62]};
    Full_Adder FA_4557(s4557, c4557, in4557_1, in4557_2, pp105[64]);
    wire[0:0] s4558, in4558_1, in4558_2;
    wire c4558;
    assign in4558_1 = {pp109[60]};
    assign in4558_2 = {pp110[59]};
    Full_Adder FA_4558(s4558, c4558, in4558_1, in4558_2, pp108[61]);
    wire[0:0] s4559, in4559_1, in4559_2;
    wire c4559;
    assign in4559_1 = {pp112[57]};
    assign in4559_2 = {pp113[56]};
    Full_Adder FA_4559(s4559, c4559, in4559_1, in4559_2, pp111[58]);
    wire[0:0] s4560, in4560_1, in4560_2;
    wire c4560;
    assign in4560_1 = {pp115[54]};
    assign in4560_2 = {pp116[53]};
    Full_Adder FA_4560(s4560, c4560, in4560_1, in4560_2, pp114[55]);
    wire[0:0] s4561, in4561_1, in4561_2;
    wire c4561;
    assign in4561_1 = {pp118[51]};
    assign in4561_2 = {pp119[50]};
    Full_Adder FA_4561(s4561, c4561, in4561_1, in4561_2, pp117[52]);
    wire[0:0] s4562, in4562_1, in4562_2;
    wire c4562;
    assign in4562_1 = {pp121[48]};
    assign in4562_2 = {pp122[47]};
    Full_Adder FA_4562(s4562, c4562, in4562_1, in4562_2, pp120[49]);
    wire[0:0] s4563, in4563_1, in4563_2;
    wire c4563;
    assign in4563_1 = {pp124[45]};
    assign in4563_2 = {pp125[44]};
    Full_Adder FA_4563(s4563, c4563, in4563_1, in4563_2, pp123[46]);
    wire[0:0] s4564, in4564_1, in4564_2;
    wire c4564;
    assign in4564_1 = {pp127[42]};
    assign in4564_2 = {c1804};
    Full_Adder FA_4564(s4564, c4564, in4564_1, in4564_2, pp126[43]);
    wire[0:0] s4565, in4565_1, in4565_2;
    wire c4565;
    assign in4565_1 = {pp44[126]};
    assign in4565_2 = {pp45[125]};
    Full_Adder FA_4565(s4565, c4565, in4565_1, in4565_2, pp43[127]);
    wire[0:0] s4566, in4566_1, in4566_2;
    wire c4566;
    assign in4566_1 = {pp47[123]};
    assign in4566_2 = {pp48[122]};
    Full_Adder FA_4566(s4566, c4566, in4566_1, in4566_2, pp46[124]);
    wire[0:0] s4567, in4567_1, in4567_2;
    wire c4567;
    assign in4567_1 = {pp50[120]};
    assign in4567_2 = {pp51[119]};
    Full_Adder FA_4567(s4567, c4567, in4567_1, in4567_2, pp49[121]);
    wire[0:0] s4568, in4568_1, in4568_2;
    wire c4568;
    assign in4568_1 = {pp53[117]};
    assign in4568_2 = {pp54[116]};
    Full_Adder FA_4568(s4568, c4568, in4568_1, in4568_2, pp52[118]);
    wire[0:0] s4569, in4569_1, in4569_2;
    wire c4569;
    assign in4569_1 = {pp56[114]};
    assign in4569_2 = {pp57[113]};
    Full_Adder FA_4569(s4569, c4569, in4569_1, in4569_2, pp55[115]);
    wire[0:0] s4570, in4570_1, in4570_2;
    wire c4570;
    assign in4570_1 = {pp59[111]};
    assign in4570_2 = {pp60[110]};
    Full_Adder FA_4570(s4570, c4570, in4570_1, in4570_2, pp58[112]);
    wire[0:0] s4571, in4571_1, in4571_2;
    wire c4571;
    assign in4571_1 = {pp62[108]};
    assign in4571_2 = {pp63[107]};
    Full_Adder FA_4571(s4571, c4571, in4571_1, in4571_2, pp61[109]);
    wire[0:0] s4572, in4572_1, in4572_2;
    wire c4572;
    assign in4572_1 = {pp65[105]};
    assign in4572_2 = {pp66[104]};
    Full_Adder FA_4572(s4572, c4572, in4572_1, in4572_2, pp64[106]);
    wire[0:0] s4573, in4573_1, in4573_2;
    wire c4573;
    assign in4573_1 = {pp68[102]};
    assign in4573_2 = {pp69[101]};
    Full_Adder FA_4573(s4573, c4573, in4573_1, in4573_2, pp67[103]);
    wire[0:0] s4574, in4574_1, in4574_2;
    wire c4574;
    assign in4574_1 = {pp71[99]};
    assign in4574_2 = {pp72[98]};
    Full_Adder FA_4574(s4574, c4574, in4574_1, in4574_2, pp70[100]);
    wire[0:0] s4575, in4575_1, in4575_2;
    wire c4575;
    assign in4575_1 = {pp74[96]};
    assign in4575_2 = {pp75[95]};
    Full_Adder FA_4575(s4575, c4575, in4575_1, in4575_2, pp73[97]);
    wire[0:0] s4576, in4576_1, in4576_2;
    wire c4576;
    assign in4576_1 = {pp77[93]};
    assign in4576_2 = {pp78[92]};
    Full_Adder FA_4576(s4576, c4576, in4576_1, in4576_2, pp76[94]);
    wire[0:0] s4577, in4577_1, in4577_2;
    wire c4577;
    assign in4577_1 = {pp80[90]};
    assign in4577_2 = {pp81[89]};
    Full_Adder FA_4577(s4577, c4577, in4577_1, in4577_2, pp79[91]);
    wire[0:0] s4578, in4578_1, in4578_2;
    wire c4578;
    assign in4578_1 = {pp83[87]};
    assign in4578_2 = {pp84[86]};
    Full_Adder FA_4578(s4578, c4578, in4578_1, in4578_2, pp82[88]);
    wire[0:0] s4579, in4579_1, in4579_2;
    wire c4579;
    assign in4579_1 = {pp86[84]};
    assign in4579_2 = {pp87[83]};
    Full_Adder FA_4579(s4579, c4579, in4579_1, in4579_2, pp85[85]);
    wire[0:0] s4580, in4580_1, in4580_2;
    wire c4580;
    assign in4580_1 = {pp89[81]};
    assign in4580_2 = {pp90[80]};
    Full_Adder FA_4580(s4580, c4580, in4580_1, in4580_2, pp88[82]);
    wire[0:0] s4581, in4581_1, in4581_2;
    wire c4581;
    assign in4581_1 = {pp92[78]};
    assign in4581_2 = {pp93[77]};
    Full_Adder FA_4581(s4581, c4581, in4581_1, in4581_2, pp91[79]);
    wire[0:0] s4582, in4582_1, in4582_2;
    wire c4582;
    assign in4582_1 = {pp95[75]};
    assign in4582_2 = {pp96[74]};
    Full_Adder FA_4582(s4582, c4582, in4582_1, in4582_2, pp94[76]);
    wire[0:0] s4583, in4583_1, in4583_2;
    wire c4583;
    assign in4583_1 = {pp98[72]};
    assign in4583_2 = {pp99[71]};
    Full_Adder FA_4583(s4583, c4583, in4583_1, in4583_2, pp97[73]);
    wire[0:0] s4584, in4584_1, in4584_2;
    wire c4584;
    assign in4584_1 = {pp101[69]};
    assign in4584_2 = {pp102[68]};
    Full_Adder FA_4584(s4584, c4584, in4584_1, in4584_2, pp100[70]);
    wire[0:0] s4585, in4585_1, in4585_2;
    wire c4585;
    assign in4585_1 = {pp104[66]};
    assign in4585_2 = {pp105[65]};
    Full_Adder FA_4585(s4585, c4585, in4585_1, in4585_2, pp103[67]);
    wire[0:0] s4586, in4586_1, in4586_2;
    wire c4586;
    assign in4586_1 = {pp107[63]};
    assign in4586_2 = {pp108[62]};
    Full_Adder FA_4586(s4586, c4586, in4586_1, in4586_2, pp106[64]);
    wire[0:0] s4587, in4587_1, in4587_2;
    wire c4587;
    assign in4587_1 = {pp110[60]};
    assign in4587_2 = {pp111[59]};
    Full_Adder FA_4587(s4587, c4587, in4587_1, in4587_2, pp109[61]);
    wire[0:0] s4588, in4588_1, in4588_2;
    wire c4588;
    assign in4588_1 = {pp113[57]};
    assign in4588_2 = {pp114[56]};
    Full_Adder FA_4588(s4588, c4588, in4588_1, in4588_2, pp112[58]);
    wire[0:0] s4589, in4589_1, in4589_2;
    wire c4589;
    assign in4589_1 = {pp116[54]};
    assign in4589_2 = {pp117[53]};
    Full_Adder FA_4589(s4589, c4589, in4589_1, in4589_2, pp115[55]);
    wire[0:0] s4590, in4590_1, in4590_2;
    wire c4590;
    assign in4590_1 = {pp119[51]};
    assign in4590_2 = {pp120[50]};
    Full_Adder FA_4590(s4590, c4590, in4590_1, in4590_2, pp118[52]);
    wire[0:0] s4591, in4591_1, in4591_2;
    wire c4591;
    assign in4591_1 = {pp122[48]};
    assign in4591_2 = {pp123[47]};
    Full_Adder FA_4591(s4591, c4591, in4591_1, in4591_2, pp121[49]);
    wire[0:0] s4592, in4592_1, in4592_2;
    wire c4592;
    assign in4592_1 = {pp125[45]};
    assign in4592_2 = {pp126[44]};
    Full_Adder FA_4592(s4592, c4592, in4592_1, in4592_2, pp124[46]);
    wire[0:0] s4593, in4593_1, in4593_2;
    wire c4593;
    assign in4593_1 = {pp45[126]};
    assign in4593_2 = {pp46[125]};
    Full_Adder FA_4593(s4593, c4593, in4593_1, in4593_2, pp44[127]);
    wire[0:0] s4594, in4594_1, in4594_2;
    wire c4594;
    assign in4594_1 = {pp48[123]};
    assign in4594_2 = {pp49[122]};
    Full_Adder FA_4594(s4594, c4594, in4594_1, in4594_2, pp47[124]);
    wire[0:0] s4595, in4595_1, in4595_2;
    wire c4595;
    assign in4595_1 = {pp51[120]};
    assign in4595_2 = {pp52[119]};
    Full_Adder FA_4595(s4595, c4595, in4595_1, in4595_2, pp50[121]);
    wire[0:0] s4596, in4596_1, in4596_2;
    wire c4596;
    assign in4596_1 = {pp54[117]};
    assign in4596_2 = {pp55[116]};
    Full_Adder FA_4596(s4596, c4596, in4596_1, in4596_2, pp53[118]);
    wire[0:0] s4597, in4597_1, in4597_2;
    wire c4597;
    assign in4597_1 = {pp57[114]};
    assign in4597_2 = {pp58[113]};
    Full_Adder FA_4597(s4597, c4597, in4597_1, in4597_2, pp56[115]);
    wire[0:0] s4598, in4598_1, in4598_2;
    wire c4598;
    assign in4598_1 = {pp60[111]};
    assign in4598_2 = {pp61[110]};
    Full_Adder FA_4598(s4598, c4598, in4598_1, in4598_2, pp59[112]);
    wire[0:0] s4599, in4599_1, in4599_2;
    wire c4599;
    assign in4599_1 = {pp63[108]};
    assign in4599_2 = {pp64[107]};
    Full_Adder FA_4599(s4599, c4599, in4599_1, in4599_2, pp62[109]);
    wire[0:0] s4600, in4600_1, in4600_2;
    wire c4600;
    assign in4600_1 = {pp66[105]};
    assign in4600_2 = {pp67[104]};
    Full_Adder FA_4600(s4600, c4600, in4600_1, in4600_2, pp65[106]);
    wire[0:0] s4601, in4601_1, in4601_2;
    wire c4601;
    assign in4601_1 = {pp69[102]};
    assign in4601_2 = {pp70[101]};
    Full_Adder FA_4601(s4601, c4601, in4601_1, in4601_2, pp68[103]);
    wire[0:0] s4602, in4602_1, in4602_2;
    wire c4602;
    assign in4602_1 = {pp72[99]};
    assign in4602_2 = {pp73[98]};
    Full_Adder FA_4602(s4602, c4602, in4602_1, in4602_2, pp71[100]);
    wire[0:0] s4603, in4603_1, in4603_2;
    wire c4603;
    assign in4603_1 = {pp75[96]};
    assign in4603_2 = {pp76[95]};
    Full_Adder FA_4603(s4603, c4603, in4603_1, in4603_2, pp74[97]);
    wire[0:0] s4604, in4604_1, in4604_2;
    wire c4604;
    assign in4604_1 = {pp78[93]};
    assign in4604_2 = {pp79[92]};
    Full_Adder FA_4604(s4604, c4604, in4604_1, in4604_2, pp77[94]);
    wire[0:0] s4605, in4605_1, in4605_2;
    wire c4605;
    assign in4605_1 = {pp81[90]};
    assign in4605_2 = {pp82[89]};
    Full_Adder FA_4605(s4605, c4605, in4605_1, in4605_2, pp80[91]);
    wire[0:0] s4606, in4606_1, in4606_2;
    wire c4606;
    assign in4606_1 = {pp84[87]};
    assign in4606_2 = {pp85[86]};
    Full_Adder FA_4606(s4606, c4606, in4606_1, in4606_2, pp83[88]);
    wire[0:0] s4607, in4607_1, in4607_2;
    wire c4607;
    assign in4607_1 = {pp87[84]};
    assign in4607_2 = {pp88[83]};
    Full_Adder FA_4607(s4607, c4607, in4607_1, in4607_2, pp86[85]);
    wire[0:0] s4608, in4608_1, in4608_2;
    wire c4608;
    assign in4608_1 = {pp90[81]};
    assign in4608_2 = {pp91[80]};
    Full_Adder FA_4608(s4608, c4608, in4608_1, in4608_2, pp89[82]);
    wire[0:0] s4609, in4609_1, in4609_2;
    wire c4609;
    assign in4609_1 = {pp93[78]};
    assign in4609_2 = {pp94[77]};
    Full_Adder FA_4609(s4609, c4609, in4609_1, in4609_2, pp92[79]);
    wire[0:0] s4610, in4610_1, in4610_2;
    wire c4610;
    assign in4610_1 = {pp96[75]};
    assign in4610_2 = {pp97[74]};
    Full_Adder FA_4610(s4610, c4610, in4610_1, in4610_2, pp95[76]);
    wire[0:0] s4611, in4611_1, in4611_2;
    wire c4611;
    assign in4611_1 = {pp99[72]};
    assign in4611_2 = {pp100[71]};
    Full_Adder FA_4611(s4611, c4611, in4611_1, in4611_2, pp98[73]);
    wire[0:0] s4612, in4612_1, in4612_2;
    wire c4612;
    assign in4612_1 = {pp102[69]};
    assign in4612_2 = {pp103[68]};
    Full_Adder FA_4612(s4612, c4612, in4612_1, in4612_2, pp101[70]);
    wire[0:0] s4613, in4613_1, in4613_2;
    wire c4613;
    assign in4613_1 = {pp105[66]};
    assign in4613_2 = {pp106[65]};
    Full_Adder FA_4613(s4613, c4613, in4613_1, in4613_2, pp104[67]);
    wire[0:0] s4614, in4614_1, in4614_2;
    wire c4614;
    assign in4614_1 = {pp108[63]};
    assign in4614_2 = {pp109[62]};
    Full_Adder FA_4614(s4614, c4614, in4614_1, in4614_2, pp107[64]);
    wire[0:0] s4615, in4615_1, in4615_2;
    wire c4615;
    assign in4615_1 = {pp111[60]};
    assign in4615_2 = {pp112[59]};
    Full_Adder FA_4615(s4615, c4615, in4615_1, in4615_2, pp110[61]);
    wire[0:0] s4616, in4616_1, in4616_2;
    wire c4616;
    assign in4616_1 = {pp114[57]};
    assign in4616_2 = {pp115[56]};
    Full_Adder FA_4616(s4616, c4616, in4616_1, in4616_2, pp113[58]);
    wire[0:0] s4617, in4617_1, in4617_2;
    wire c4617;
    assign in4617_1 = {pp117[54]};
    assign in4617_2 = {pp118[53]};
    Full_Adder FA_4617(s4617, c4617, in4617_1, in4617_2, pp116[55]);
    wire[0:0] s4618, in4618_1, in4618_2;
    wire c4618;
    assign in4618_1 = {pp120[51]};
    assign in4618_2 = {pp121[50]};
    Full_Adder FA_4618(s4618, c4618, in4618_1, in4618_2, pp119[52]);
    wire[0:0] s4619, in4619_1, in4619_2;
    wire c4619;
    assign in4619_1 = {pp123[48]};
    assign in4619_2 = {pp124[47]};
    Full_Adder FA_4619(s4619, c4619, in4619_1, in4619_2, pp122[49]);
    wire[0:0] s4620, in4620_1, in4620_2;
    wire c4620;
    assign in4620_1 = {pp46[126]};
    assign in4620_2 = {pp47[125]};
    Full_Adder FA_4620(s4620, c4620, in4620_1, in4620_2, pp45[127]);
    wire[0:0] s4621, in4621_1, in4621_2;
    wire c4621;
    assign in4621_1 = {pp49[123]};
    assign in4621_2 = {pp50[122]};
    Full_Adder FA_4621(s4621, c4621, in4621_1, in4621_2, pp48[124]);
    wire[0:0] s4622, in4622_1, in4622_2;
    wire c4622;
    assign in4622_1 = {pp52[120]};
    assign in4622_2 = {pp53[119]};
    Full_Adder FA_4622(s4622, c4622, in4622_1, in4622_2, pp51[121]);
    wire[0:0] s4623, in4623_1, in4623_2;
    wire c4623;
    assign in4623_1 = {pp55[117]};
    assign in4623_2 = {pp56[116]};
    Full_Adder FA_4623(s4623, c4623, in4623_1, in4623_2, pp54[118]);
    wire[0:0] s4624, in4624_1, in4624_2;
    wire c4624;
    assign in4624_1 = {pp58[114]};
    assign in4624_2 = {pp59[113]};
    Full_Adder FA_4624(s4624, c4624, in4624_1, in4624_2, pp57[115]);
    wire[0:0] s4625, in4625_1, in4625_2;
    wire c4625;
    assign in4625_1 = {pp61[111]};
    assign in4625_2 = {pp62[110]};
    Full_Adder FA_4625(s4625, c4625, in4625_1, in4625_2, pp60[112]);
    wire[0:0] s4626, in4626_1, in4626_2;
    wire c4626;
    assign in4626_1 = {pp64[108]};
    assign in4626_2 = {pp65[107]};
    Full_Adder FA_4626(s4626, c4626, in4626_1, in4626_2, pp63[109]);
    wire[0:0] s4627, in4627_1, in4627_2;
    wire c4627;
    assign in4627_1 = {pp67[105]};
    assign in4627_2 = {pp68[104]};
    Full_Adder FA_4627(s4627, c4627, in4627_1, in4627_2, pp66[106]);
    wire[0:0] s4628, in4628_1, in4628_2;
    wire c4628;
    assign in4628_1 = {pp70[102]};
    assign in4628_2 = {pp71[101]};
    Full_Adder FA_4628(s4628, c4628, in4628_1, in4628_2, pp69[103]);
    wire[0:0] s4629, in4629_1, in4629_2;
    wire c4629;
    assign in4629_1 = {pp73[99]};
    assign in4629_2 = {pp74[98]};
    Full_Adder FA_4629(s4629, c4629, in4629_1, in4629_2, pp72[100]);
    wire[0:0] s4630, in4630_1, in4630_2;
    wire c4630;
    assign in4630_1 = {pp76[96]};
    assign in4630_2 = {pp77[95]};
    Full_Adder FA_4630(s4630, c4630, in4630_1, in4630_2, pp75[97]);
    wire[0:0] s4631, in4631_1, in4631_2;
    wire c4631;
    assign in4631_1 = {pp79[93]};
    assign in4631_2 = {pp80[92]};
    Full_Adder FA_4631(s4631, c4631, in4631_1, in4631_2, pp78[94]);
    wire[0:0] s4632, in4632_1, in4632_2;
    wire c4632;
    assign in4632_1 = {pp82[90]};
    assign in4632_2 = {pp83[89]};
    Full_Adder FA_4632(s4632, c4632, in4632_1, in4632_2, pp81[91]);
    wire[0:0] s4633, in4633_1, in4633_2;
    wire c4633;
    assign in4633_1 = {pp85[87]};
    assign in4633_2 = {pp86[86]};
    Full_Adder FA_4633(s4633, c4633, in4633_1, in4633_2, pp84[88]);
    wire[0:0] s4634, in4634_1, in4634_2;
    wire c4634;
    assign in4634_1 = {pp88[84]};
    assign in4634_2 = {pp89[83]};
    Full_Adder FA_4634(s4634, c4634, in4634_1, in4634_2, pp87[85]);
    wire[0:0] s4635, in4635_1, in4635_2;
    wire c4635;
    assign in4635_1 = {pp91[81]};
    assign in4635_2 = {pp92[80]};
    Full_Adder FA_4635(s4635, c4635, in4635_1, in4635_2, pp90[82]);
    wire[0:0] s4636, in4636_1, in4636_2;
    wire c4636;
    assign in4636_1 = {pp94[78]};
    assign in4636_2 = {pp95[77]};
    Full_Adder FA_4636(s4636, c4636, in4636_1, in4636_2, pp93[79]);
    wire[0:0] s4637, in4637_1, in4637_2;
    wire c4637;
    assign in4637_1 = {pp97[75]};
    assign in4637_2 = {pp98[74]};
    Full_Adder FA_4637(s4637, c4637, in4637_1, in4637_2, pp96[76]);
    wire[0:0] s4638, in4638_1, in4638_2;
    wire c4638;
    assign in4638_1 = {pp100[72]};
    assign in4638_2 = {pp101[71]};
    Full_Adder FA_4638(s4638, c4638, in4638_1, in4638_2, pp99[73]);
    wire[0:0] s4639, in4639_1, in4639_2;
    wire c4639;
    assign in4639_1 = {pp103[69]};
    assign in4639_2 = {pp104[68]};
    Full_Adder FA_4639(s4639, c4639, in4639_1, in4639_2, pp102[70]);
    wire[0:0] s4640, in4640_1, in4640_2;
    wire c4640;
    assign in4640_1 = {pp106[66]};
    assign in4640_2 = {pp107[65]};
    Full_Adder FA_4640(s4640, c4640, in4640_1, in4640_2, pp105[67]);
    wire[0:0] s4641, in4641_1, in4641_2;
    wire c4641;
    assign in4641_1 = {pp109[63]};
    assign in4641_2 = {pp110[62]};
    Full_Adder FA_4641(s4641, c4641, in4641_1, in4641_2, pp108[64]);
    wire[0:0] s4642, in4642_1, in4642_2;
    wire c4642;
    assign in4642_1 = {pp112[60]};
    assign in4642_2 = {pp113[59]};
    Full_Adder FA_4642(s4642, c4642, in4642_1, in4642_2, pp111[61]);
    wire[0:0] s4643, in4643_1, in4643_2;
    wire c4643;
    assign in4643_1 = {pp115[57]};
    assign in4643_2 = {pp116[56]};
    Full_Adder FA_4643(s4643, c4643, in4643_1, in4643_2, pp114[58]);
    wire[0:0] s4644, in4644_1, in4644_2;
    wire c4644;
    assign in4644_1 = {pp118[54]};
    assign in4644_2 = {pp119[53]};
    Full_Adder FA_4644(s4644, c4644, in4644_1, in4644_2, pp117[55]);
    wire[0:0] s4645, in4645_1, in4645_2;
    wire c4645;
    assign in4645_1 = {pp121[51]};
    assign in4645_2 = {pp122[50]};
    Full_Adder FA_4645(s4645, c4645, in4645_1, in4645_2, pp120[52]);
    wire[0:0] s4646, in4646_1, in4646_2;
    wire c4646;
    assign in4646_1 = {pp47[126]};
    assign in4646_2 = {pp48[125]};
    Full_Adder FA_4646(s4646, c4646, in4646_1, in4646_2, pp46[127]);
    wire[0:0] s4647, in4647_1, in4647_2;
    wire c4647;
    assign in4647_1 = {pp50[123]};
    assign in4647_2 = {pp51[122]};
    Full_Adder FA_4647(s4647, c4647, in4647_1, in4647_2, pp49[124]);
    wire[0:0] s4648, in4648_1, in4648_2;
    wire c4648;
    assign in4648_1 = {pp53[120]};
    assign in4648_2 = {pp54[119]};
    Full_Adder FA_4648(s4648, c4648, in4648_1, in4648_2, pp52[121]);
    wire[0:0] s4649, in4649_1, in4649_2;
    wire c4649;
    assign in4649_1 = {pp56[117]};
    assign in4649_2 = {pp57[116]};
    Full_Adder FA_4649(s4649, c4649, in4649_1, in4649_2, pp55[118]);
    wire[0:0] s4650, in4650_1, in4650_2;
    wire c4650;
    assign in4650_1 = {pp59[114]};
    assign in4650_2 = {pp60[113]};
    Full_Adder FA_4650(s4650, c4650, in4650_1, in4650_2, pp58[115]);
    wire[0:0] s4651, in4651_1, in4651_2;
    wire c4651;
    assign in4651_1 = {pp62[111]};
    assign in4651_2 = {pp63[110]};
    Full_Adder FA_4651(s4651, c4651, in4651_1, in4651_2, pp61[112]);
    wire[0:0] s4652, in4652_1, in4652_2;
    wire c4652;
    assign in4652_1 = {pp65[108]};
    assign in4652_2 = {pp66[107]};
    Full_Adder FA_4652(s4652, c4652, in4652_1, in4652_2, pp64[109]);
    wire[0:0] s4653, in4653_1, in4653_2;
    wire c4653;
    assign in4653_1 = {pp68[105]};
    assign in4653_2 = {pp69[104]};
    Full_Adder FA_4653(s4653, c4653, in4653_1, in4653_2, pp67[106]);
    wire[0:0] s4654, in4654_1, in4654_2;
    wire c4654;
    assign in4654_1 = {pp71[102]};
    assign in4654_2 = {pp72[101]};
    Full_Adder FA_4654(s4654, c4654, in4654_1, in4654_2, pp70[103]);
    wire[0:0] s4655, in4655_1, in4655_2;
    wire c4655;
    assign in4655_1 = {pp74[99]};
    assign in4655_2 = {pp75[98]};
    Full_Adder FA_4655(s4655, c4655, in4655_1, in4655_2, pp73[100]);
    wire[0:0] s4656, in4656_1, in4656_2;
    wire c4656;
    assign in4656_1 = {pp77[96]};
    assign in4656_2 = {pp78[95]};
    Full_Adder FA_4656(s4656, c4656, in4656_1, in4656_2, pp76[97]);
    wire[0:0] s4657, in4657_1, in4657_2;
    wire c4657;
    assign in4657_1 = {pp80[93]};
    assign in4657_2 = {pp81[92]};
    Full_Adder FA_4657(s4657, c4657, in4657_1, in4657_2, pp79[94]);
    wire[0:0] s4658, in4658_1, in4658_2;
    wire c4658;
    assign in4658_1 = {pp83[90]};
    assign in4658_2 = {pp84[89]};
    Full_Adder FA_4658(s4658, c4658, in4658_1, in4658_2, pp82[91]);
    wire[0:0] s4659, in4659_1, in4659_2;
    wire c4659;
    assign in4659_1 = {pp86[87]};
    assign in4659_2 = {pp87[86]};
    Full_Adder FA_4659(s4659, c4659, in4659_1, in4659_2, pp85[88]);
    wire[0:0] s4660, in4660_1, in4660_2;
    wire c4660;
    assign in4660_1 = {pp89[84]};
    assign in4660_2 = {pp90[83]};
    Full_Adder FA_4660(s4660, c4660, in4660_1, in4660_2, pp88[85]);
    wire[0:0] s4661, in4661_1, in4661_2;
    wire c4661;
    assign in4661_1 = {pp92[81]};
    assign in4661_2 = {pp93[80]};
    Full_Adder FA_4661(s4661, c4661, in4661_1, in4661_2, pp91[82]);
    wire[0:0] s4662, in4662_1, in4662_2;
    wire c4662;
    assign in4662_1 = {pp95[78]};
    assign in4662_2 = {pp96[77]};
    Full_Adder FA_4662(s4662, c4662, in4662_1, in4662_2, pp94[79]);
    wire[0:0] s4663, in4663_1, in4663_2;
    wire c4663;
    assign in4663_1 = {pp98[75]};
    assign in4663_2 = {pp99[74]};
    Full_Adder FA_4663(s4663, c4663, in4663_1, in4663_2, pp97[76]);
    wire[0:0] s4664, in4664_1, in4664_2;
    wire c4664;
    assign in4664_1 = {pp101[72]};
    assign in4664_2 = {pp102[71]};
    Full_Adder FA_4664(s4664, c4664, in4664_1, in4664_2, pp100[73]);
    wire[0:0] s4665, in4665_1, in4665_2;
    wire c4665;
    assign in4665_1 = {pp104[69]};
    assign in4665_2 = {pp105[68]};
    Full_Adder FA_4665(s4665, c4665, in4665_1, in4665_2, pp103[70]);
    wire[0:0] s4666, in4666_1, in4666_2;
    wire c4666;
    assign in4666_1 = {pp107[66]};
    assign in4666_2 = {pp108[65]};
    Full_Adder FA_4666(s4666, c4666, in4666_1, in4666_2, pp106[67]);
    wire[0:0] s4667, in4667_1, in4667_2;
    wire c4667;
    assign in4667_1 = {pp110[63]};
    assign in4667_2 = {pp111[62]};
    Full_Adder FA_4667(s4667, c4667, in4667_1, in4667_2, pp109[64]);
    wire[0:0] s4668, in4668_1, in4668_2;
    wire c4668;
    assign in4668_1 = {pp113[60]};
    assign in4668_2 = {pp114[59]};
    Full_Adder FA_4668(s4668, c4668, in4668_1, in4668_2, pp112[61]);
    wire[0:0] s4669, in4669_1, in4669_2;
    wire c4669;
    assign in4669_1 = {pp116[57]};
    assign in4669_2 = {pp117[56]};
    Full_Adder FA_4669(s4669, c4669, in4669_1, in4669_2, pp115[58]);
    wire[0:0] s4670, in4670_1, in4670_2;
    wire c4670;
    assign in4670_1 = {pp119[54]};
    assign in4670_2 = {pp120[53]};
    Full_Adder FA_4670(s4670, c4670, in4670_1, in4670_2, pp118[55]);
    wire[0:0] s4671, in4671_1, in4671_2;
    wire c4671;
    assign in4671_1 = {pp48[126]};
    assign in4671_2 = {pp49[125]};
    Full_Adder FA_4671(s4671, c4671, in4671_1, in4671_2, pp47[127]);
    wire[0:0] s4672, in4672_1, in4672_2;
    wire c4672;
    assign in4672_1 = {pp51[123]};
    assign in4672_2 = {pp52[122]};
    Full_Adder FA_4672(s4672, c4672, in4672_1, in4672_2, pp50[124]);
    wire[0:0] s4673, in4673_1, in4673_2;
    wire c4673;
    assign in4673_1 = {pp54[120]};
    assign in4673_2 = {pp55[119]};
    Full_Adder FA_4673(s4673, c4673, in4673_1, in4673_2, pp53[121]);
    wire[0:0] s4674, in4674_1, in4674_2;
    wire c4674;
    assign in4674_1 = {pp57[117]};
    assign in4674_2 = {pp58[116]};
    Full_Adder FA_4674(s4674, c4674, in4674_1, in4674_2, pp56[118]);
    wire[0:0] s4675, in4675_1, in4675_2;
    wire c4675;
    assign in4675_1 = {pp60[114]};
    assign in4675_2 = {pp61[113]};
    Full_Adder FA_4675(s4675, c4675, in4675_1, in4675_2, pp59[115]);
    wire[0:0] s4676, in4676_1, in4676_2;
    wire c4676;
    assign in4676_1 = {pp63[111]};
    assign in4676_2 = {pp64[110]};
    Full_Adder FA_4676(s4676, c4676, in4676_1, in4676_2, pp62[112]);
    wire[0:0] s4677, in4677_1, in4677_2;
    wire c4677;
    assign in4677_1 = {pp66[108]};
    assign in4677_2 = {pp67[107]};
    Full_Adder FA_4677(s4677, c4677, in4677_1, in4677_2, pp65[109]);
    wire[0:0] s4678, in4678_1, in4678_2;
    wire c4678;
    assign in4678_1 = {pp69[105]};
    assign in4678_2 = {pp70[104]};
    Full_Adder FA_4678(s4678, c4678, in4678_1, in4678_2, pp68[106]);
    wire[0:0] s4679, in4679_1, in4679_2;
    wire c4679;
    assign in4679_1 = {pp72[102]};
    assign in4679_2 = {pp73[101]};
    Full_Adder FA_4679(s4679, c4679, in4679_1, in4679_2, pp71[103]);
    wire[0:0] s4680, in4680_1, in4680_2;
    wire c4680;
    assign in4680_1 = {pp75[99]};
    assign in4680_2 = {pp76[98]};
    Full_Adder FA_4680(s4680, c4680, in4680_1, in4680_2, pp74[100]);
    wire[0:0] s4681, in4681_1, in4681_2;
    wire c4681;
    assign in4681_1 = {pp78[96]};
    assign in4681_2 = {pp79[95]};
    Full_Adder FA_4681(s4681, c4681, in4681_1, in4681_2, pp77[97]);
    wire[0:0] s4682, in4682_1, in4682_2;
    wire c4682;
    assign in4682_1 = {pp81[93]};
    assign in4682_2 = {pp82[92]};
    Full_Adder FA_4682(s4682, c4682, in4682_1, in4682_2, pp80[94]);
    wire[0:0] s4683, in4683_1, in4683_2;
    wire c4683;
    assign in4683_1 = {pp84[90]};
    assign in4683_2 = {pp85[89]};
    Full_Adder FA_4683(s4683, c4683, in4683_1, in4683_2, pp83[91]);
    wire[0:0] s4684, in4684_1, in4684_2;
    wire c4684;
    assign in4684_1 = {pp87[87]};
    assign in4684_2 = {pp88[86]};
    Full_Adder FA_4684(s4684, c4684, in4684_1, in4684_2, pp86[88]);
    wire[0:0] s4685, in4685_1, in4685_2;
    wire c4685;
    assign in4685_1 = {pp90[84]};
    assign in4685_2 = {pp91[83]};
    Full_Adder FA_4685(s4685, c4685, in4685_1, in4685_2, pp89[85]);
    wire[0:0] s4686, in4686_1, in4686_2;
    wire c4686;
    assign in4686_1 = {pp93[81]};
    assign in4686_2 = {pp94[80]};
    Full_Adder FA_4686(s4686, c4686, in4686_1, in4686_2, pp92[82]);
    wire[0:0] s4687, in4687_1, in4687_2;
    wire c4687;
    assign in4687_1 = {pp96[78]};
    assign in4687_2 = {pp97[77]};
    Full_Adder FA_4687(s4687, c4687, in4687_1, in4687_2, pp95[79]);
    wire[0:0] s4688, in4688_1, in4688_2;
    wire c4688;
    assign in4688_1 = {pp99[75]};
    assign in4688_2 = {pp100[74]};
    Full_Adder FA_4688(s4688, c4688, in4688_1, in4688_2, pp98[76]);
    wire[0:0] s4689, in4689_1, in4689_2;
    wire c4689;
    assign in4689_1 = {pp102[72]};
    assign in4689_2 = {pp103[71]};
    Full_Adder FA_4689(s4689, c4689, in4689_1, in4689_2, pp101[73]);
    wire[0:0] s4690, in4690_1, in4690_2;
    wire c4690;
    assign in4690_1 = {pp105[69]};
    assign in4690_2 = {pp106[68]};
    Full_Adder FA_4690(s4690, c4690, in4690_1, in4690_2, pp104[70]);
    wire[0:0] s4691, in4691_1, in4691_2;
    wire c4691;
    assign in4691_1 = {pp108[66]};
    assign in4691_2 = {pp109[65]};
    Full_Adder FA_4691(s4691, c4691, in4691_1, in4691_2, pp107[67]);
    wire[0:0] s4692, in4692_1, in4692_2;
    wire c4692;
    assign in4692_1 = {pp111[63]};
    assign in4692_2 = {pp112[62]};
    Full_Adder FA_4692(s4692, c4692, in4692_1, in4692_2, pp110[64]);
    wire[0:0] s4693, in4693_1, in4693_2;
    wire c4693;
    assign in4693_1 = {pp114[60]};
    assign in4693_2 = {pp115[59]};
    Full_Adder FA_4693(s4693, c4693, in4693_1, in4693_2, pp113[61]);
    wire[0:0] s4694, in4694_1, in4694_2;
    wire c4694;
    assign in4694_1 = {pp117[57]};
    assign in4694_2 = {pp118[56]};
    Full_Adder FA_4694(s4694, c4694, in4694_1, in4694_2, pp116[58]);
    wire[0:0] s4695, in4695_1, in4695_2;
    wire c4695;
    assign in4695_1 = {pp49[126]};
    assign in4695_2 = {pp50[125]};
    Full_Adder FA_4695(s4695, c4695, in4695_1, in4695_2, pp48[127]);
    wire[0:0] s4696, in4696_1, in4696_2;
    wire c4696;
    assign in4696_1 = {pp52[123]};
    assign in4696_2 = {pp53[122]};
    Full_Adder FA_4696(s4696, c4696, in4696_1, in4696_2, pp51[124]);
    wire[0:0] s4697, in4697_1, in4697_2;
    wire c4697;
    assign in4697_1 = {pp55[120]};
    assign in4697_2 = {pp56[119]};
    Full_Adder FA_4697(s4697, c4697, in4697_1, in4697_2, pp54[121]);
    wire[0:0] s4698, in4698_1, in4698_2;
    wire c4698;
    assign in4698_1 = {pp58[117]};
    assign in4698_2 = {pp59[116]};
    Full_Adder FA_4698(s4698, c4698, in4698_1, in4698_2, pp57[118]);
    wire[0:0] s4699, in4699_1, in4699_2;
    wire c4699;
    assign in4699_1 = {pp61[114]};
    assign in4699_2 = {pp62[113]};
    Full_Adder FA_4699(s4699, c4699, in4699_1, in4699_2, pp60[115]);
    wire[0:0] s4700, in4700_1, in4700_2;
    wire c4700;
    assign in4700_1 = {pp64[111]};
    assign in4700_2 = {pp65[110]};
    Full_Adder FA_4700(s4700, c4700, in4700_1, in4700_2, pp63[112]);
    wire[0:0] s4701, in4701_1, in4701_2;
    wire c4701;
    assign in4701_1 = {pp67[108]};
    assign in4701_2 = {pp68[107]};
    Full_Adder FA_4701(s4701, c4701, in4701_1, in4701_2, pp66[109]);
    wire[0:0] s4702, in4702_1, in4702_2;
    wire c4702;
    assign in4702_1 = {pp70[105]};
    assign in4702_2 = {pp71[104]};
    Full_Adder FA_4702(s4702, c4702, in4702_1, in4702_2, pp69[106]);
    wire[0:0] s4703, in4703_1, in4703_2;
    wire c4703;
    assign in4703_1 = {pp73[102]};
    assign in4703_2 = {pp74[101]};
    Full_Adder FA_4703(s4703, c4703, in4703_1, in4703_2, pp72[103]);
    wire[0:0] s4704, in4704_1, in4704_2;
    wire c4704;
    assign in4704_1 = {pp76[99]};
    assign in4704_2 = {pp77[98]};
    Full_Adder FA_4704(s4704, c4704, in4704_1, in4704_2, pp75[100]);
    wire[0:0] s4705, in4705_1, in4705_2;
    wire c4705;
    assign in4705_1 = {pp79[96]};
    assign in4705_2 = {pp80[95]};
    Full_Adder FA_4705(s4705, c4705, in4705_1, in4705_2, pp78[97]);
    wire[0:0] s4706, in4706_1, in4706_2;
    wire c4706;
    assign in4706_1 = {pp82[93]};
    assign in4706_2 = {pp83[92]};
    Full_Adder FA_4706(s4706, c4706, in4706_1, in4706_2, pp81[94]);
    wire[0:0] s4707, in4707_1, in4707_2;
    wire c4707;
    assign in4707_1 = {pp85[90]};
    assign in4707_2 = {pp86[89]};
    Full_Adder FA_4707(s4707, c4707, in4707_1, in4707_2, pp84[91]);
    wire[0:0] s4708, in4708_1, in4708_2;
    wire c4708;
    assign in4708_1 = {pp88[87]};
    assign in4708_2 = {pp89[86]};
    Full_Adder FA_4708(s4708, c4708, in4708_1, in4708_2, pp87[88]);
    wire[0:0] s4709, in4709_1, in4709_2;
    wire c4709;
    assign in4709_1 = {pp91[84]};
    assign in4709_2 = {pp92[83]};
    Full_Adder FA_4709(s4709, c4709, in4709_1, in4709_2, pp90[85]);
    wire[0:0] s4710, in4710_1, in4710_2;
    wire c4710;
    assign in4710_1 = {pp94[81]};
    assign in4710_2 = {pp95[80]};
    Full_Adder FA_4710(s4710, c4710, in4710_1, in4710_2, pp93[82]);
    wire[0:0] s4711, in4711_1, in4711_2;
    wire c4711;
    assign in4711_1 = {pp97[78]};
    assign in4711_2 = {pp98[77]};
    Full_Adder FA_4711(s4711, c4711, in4711_1, in4711_2, pp96[79]);
    wire[0:0] s4712, in4712_1, in4712_2;
    wire c4712;
    assign in4712_1 = {pp100[75]};
    assign in4712_2 = {pp101[74]};
    Full_Adder FA_4712(s4712, c4712, in4712_1, in4712_2, pp99[76]);
    wire[0:0] s4713, in4713_1, in4713_2;
    wire c4713;
    assign in4713_1 = {pp103[72]};
    assign in4713_2 = {pp104[71]};
    Full_Adder FA_4713(s4713, c4713, in4713_1, in4713_2, pp102[73]);
    wire[0:0] s4714, in4714_1, in4714_2;
    wire c4714;
    assign in4714_1 = {pp106[69]};
    assign in4714_2 = {pp107[68]};
    Full_Adder FA_4714(s4714, c4714, in4714_1, in4714_2, pp105[70]);
    wire[0:0] s4715, in4715_1, in4715_2;
    wire c4715;
    assign in4715_1 = {pp109[66]};
    assign in4715_2 = {pp110[65]};
    Full_Adder FA_4715(s4715, c4715, in4715_1, in4715_2, pp108[67]);
    wire[0:0] s4716, in4716_1, in4716_2;
    wire c4716;
    assign in4716_1 = {pp112[63]};
    assign in4716_2 = {pp113[62]};
    Full_Adder FA_4716(s4716, c4716, in4716_1, in4716_2, pp111[64]);
    wire[0:0] s4717, in4717_1, in4717_2;
    wire c4717;
    assign in4717_1 = {pp115[60]};
    assign in4717_2 = {pp116[59]};
    Full_Adder FA_4717(s4717, c4717, in4717_1, in4717_2, pp114[61]);
    wire[0:0] s4718, in4718_1, in4718_2;
    wire c4718;
    assign in4718_1 = {pp50[126]};
    assign in4718_2 = {pp51[125]};
    Full_Adder FA_4718(s4718, c4718, in4718_1, in4718_2, pp49[127]);
    wire[0:0] s4719, in4719_1, in4719_2;
    wire c4719;
    assign in4719_1 = {pp53[123]};
    assign in4719_2 = {pp54[122]};
    Full_Adder FA_4719(s4719, c4719, in4719_1, in4719_2, pp52[124]);
    wire[0:0] s4720, in4720_1, in4720_2;
    wire c4720;
    assign in4720_1 = {pp56[120]};
    assign in4720_2 = {pp57[119]};
    Full_Adder FA_4720(s4720, c4720, in4720_1, in4720_2, pp55[121]);
    wire[0:0] s4721, in4721_1, in4721_2;
    wire c4721;
    assign in4721_1 = {pp59[117]};
    assign in4721_2 = {pp60[116]};
    Full_Adder FA_4721(s4721, c4721, in4721_1, in4721_2, pp58[118]);
    wire[0:0] s4722, in4722_1, in4722_2;
    wire c4722;
    assign in4722_1 = {pp62[114]};
    assign in4722_2 = {pp63[113]};
    Full_Adder FA_4722(s4722, c4722, in4722_1, in4722_2, pp61[115]);
    wire[0:0] s4723, in4723_1, in4723_2;
    wire c4723;
    assign in4723_1 = {pp65[111]};
    assign in4723_2 = {pp66[110]};
    Full_Adder FA_4723(s4723, c4723, in4723_1, in4723_2, pp64[112]);
    wire[0:0] s4724, in4724_1, in4724_2;
    wire c4724;
    assign in4724_1 = {pp68[108]};
    assign in4724_2 = {pp69[107]};
    Full_Adder FA_4724(s4724, c4724, in4724_1, in4724_2, pp67[109]);
    wire[0:0] s4725, in4725_1, in4725_2;
    wire c4725;
    assign in4725_1 = {pp71[105]};
    assign in4725_2 = {pp72[104]};
    Full_Adder FA_4725(s4725, c4725, in4725_1, in4725_2, pp70[106]);
    wire[0:0] s4726, in4726_1, in4726_2;
    wire c4726;
    assign in4726_1 = {pp74[102]};
    assign in4726_2 = {pp75[101]};
    Full_Adder FA_4726(s4726, c4726, in4726_1, in4726_2, pp73[103]);
    wire[0:0] s4727, in4727_1, in4727_2;
    wire c4727;
    assign in4727_1 = {pp77[99]};
    assign in4727_2 = {pp78[98]};
    Full_Adder FA_4727(s4727, c4727, in4727_1, in4727_2, pp76[100]);
    wire[0:0] s4728, in4728_1, in4728_2;
    wire c4728;
    assign in4728_1 = {pp80[96]};
    assign in4728_2 = {pp81[95]};
    Full_Adder FA_4728(s4728, c4728, in4728_1, in4728_2, pp79[97]);
    wire[0:0] s4729, in4729_1, in4729_2;
    wire c4729;
    assign in4729_1 = {pp83[93]};
    assign in4729_2 = {pp84[92]};
    Full_Adder FA_4729(s4729, c4729, in4729_1, in4729_2, pp82[94]);
    wire[0:0] s4730, in4730_1, in4730_2;
    wire c4730;
    assign in4730_1 = {pp86[90]};
    assign in4730_2 = {pp87[89]};
    Full_Adder FA_4730(s4730, c4730, in4730_1, in4730_2, pp85[91]);
    wire[0:0] s4731, in4731_1, in4731_2;
    wire c4731;
    assign in4731_1 = {pp89[87]};
    assign in4731_2 = {pp90[86]};
    Full_Adder FA_4731(s4731, c4731, in4731_1, in4731_2, pp88[88]);
    wire[0:0] s4732, in4732_1, in4732_2;
    wire c4732;
    assign in4732_1 = {pp92[84]};
    assign in4732_2 = {pp93[83]};
    Full_Adder FA_4732(s4732, c4732, in4732_1, in4732_2, pp91[85]);
    wire[0:0] s4733, in4733_1, in4733_2;
    wire c4733;
    assign in4733_1 = {pp95[81]};
    assign in4733_2 = {pp96[80]};
    Full_Adder FA_4733(s4733, c4733, in4733_1, in4733_2, pp94[82]);
    wire[0:0] s4734, in4734_1, in4734_2;
    wire c4734;
    assign in4734_1 = {pp98[78]};
    assign in4734_2 = {pp99[77]};
    Full_Adder FA_4734(s4734, c4734, in4734_1, in4734_2, pp97[79]);
    wire[0:0] s4735, in4735_1, in4735_2;
    wire c4735;
    assign in4735_1 = {pp101[75]};
    assign in4735_2 = {pp102[74]};
    Full_Adder FA_4735(s4735, c4735, in4735_1, in4735_2, pp100[76]);
    wire[0:0] s4736, in4736_1, in4736_2;
    wire c4736;
    assign in4736_1 = {pp104[72]};
    assign in4736_2 = {pp105[71]};
    Full_Adder FA_4736(s4736, c4736, in4736_1, in4736_2, pp103[73]);
    wire[0:0] s4737, in4737_1, in4737_2;
    wire c4737;
    assign in4737_1 = {pp107[69]};
    assign in4737_2 = {pp108[68]};
    Full_Adder FA_4737(s4737, c4737, in4737_1, in4737_2, pp106[70]);
    wire[0:0] s4738, in4738_1, in4738_2;
    wire c4738;
    assign in4738_1 = {pp110[66]};
    assign in4738_2 = {pp111[65]};
    Full_Adder FA_4738(s4738, c4738, in4738_1, in4738_2, pp109[67]);
    wire[0:0] s4739, in4739_1, in4739_2;
    wire c4739;
    assign in4739_1 = {pp113[63]};
    assign in4739_2 = {pp114[62]};
    Full_Adder FA_4739(s4739, c4739, in4739_1, in4739_2, pp112[64]);
    wire[0:0] s4740, in4740_1, in4740_2;
    wire c4740;
    assign in4740_1 = {pp51[126]};
    assign in4740_2 = {pp52[125]};
    Full_Adder FA_4740(s4740, c4740, in4740_1, in4740_2, pp50[127]);
    wire[0:0] s4741, in4741_1, in4741_2;
    wire c4741;
    assign in4741_1 = {pp54[123]};
    assign in4741_2 = {pp55[122]};
    Full_Adder FA_4741(s4741, c4741, in4741_1, in4741_2, pp53[124]);
    wire[0:0] s4742, in4742_1, in4742_2;
    wire c4742;
    assign in4742_1 = {pp57[120]};
    assign in4742_2 = {pp58[119]};
    Full_Adder FA_4742(s4742, c4742, in4742_1, in4742_2, pp56[121]);
    wire[0:0] s4743, in4743_1, in4743_2;
    wire c4743;
    assign in4743_1 = {pp60[117]};
    assign in4743_2 = {pp61[116]};
    Full_Adder FA_4743(s4743, c4743, in4743_1, in4743_2, pp59[118]);
    wire[0:0] s4744, in4744_1, in4744_2;
    wire c4744;
    assign in4744_1 = {pp63[114]};
    assign in4744_2 = {pp64[113]};
    Full_Adder FA_4744(s4744, c4744, in4744_1, in4744_2, pp62[115]);
    wire[0:0] s4745, in4745_1, in4745_2;
    wire c4745;
    assign in4745_1 = {pp66[111]};
    assign in4745_2 = {pp67[110]};
    Full_Adder FA_4745(s4745, c4745, in4745_1, in4745_2, pp65[112]);
    wire[0:0] s4746, in4746_1, in4746_2;
    wire c4746;
    assign in4746_1 = {pp69[108]};
    assign in4746_2 = {pp70[107]};
    Full_Adder FA_4746(s4746, c4746, in4746_1, in4746_2, pp68[109]);
    wire[0:0] s4747, in4747_1, in4747_2;
    wire c4747;
    assign in4747_1 = {pp72[105]};
    assign in4747_2 = {pp73[104]};
    Full_Adder FA_4747(s4747, c4747, in4747_1, in4747_2, pp71[106]);
    wire[0:0] s4748, in4748_1, in4748_2;
    wire c4748;
    assign in4748_1 = {pp75[102]};
    assign in4748_2 = {pp76[101]};
    Full_Adder FA_4748(s4748, c4748, in4748_1, in4748_2, pp74[103]);
    wire[0:0] s4749, in4749_1, in4749_2;
    wire c4749;
    assign in4749_1 = {pp78[99]};
    assign in4749_2 = {pp79[98]};
    Full_Adder FA_4749(s4749, c4749, in4749_1, in4749_2, pp77[100]);
    wire[0:0] s4750, in4750_1, in4750_2;
    wire c4750;
    assign in4750_1 = {pp81[96]};
    assign in4750_2 = {pp82[95]};
    Full_Adder FA_4750(s4750, c4750, in4750_1, in4750_2, pp80[97]);
    wire[0:0] s4751, in4751_1, in4751_2;
    wire c4751;
    assign in4751_1 = {pp84[93]};
    assign in4751_2 = {pp85[92]};
    Full_Adder FA_4751(s4751, c4751, in4751_1, in4751_2, pp83[94]);
    wire[0:0] s4752, in4752_1, in4752_2;
    wire c4752;
    assign in4752_1 = {pp87[90]};
    assign in4752_2 = {pp88[89]};
    Full_Adder FA_4752(s4752, c4752, in4752_1, in4752_2, pp86[91]);
    wire[0:0] s4753, in4753_1, in4753_2;
    wire c4753;
    assign in4753_1 = {pp90[87]};
    assign in4753_2 = {pp91[86]};
    Full_Adder FA_4753(s4753, c4753, in4753_1, in4753_2, pp89[88]);
    wire[0:0] s4754, in4754_1, in4754_2;
    wire c4754;
    assign in4754_1 = {pp93[84]};
    assign in4754_2 = {pp94[83]};
    Full_Adder FA_4754(s4754, c4754, in4754_1, in4754_2, pp92[85]);
    wire[0:0] s4755, in4755_1, in4755_2;
    wire c4755;
    assign in4755_1 = {pp96[81]};
    assign in4755_2 = {pp97[80]};
    Full_Adder FA_4755(s4755, c4755, in4755_1, in4755_2, pp95[82]);
    wire[0:0] s4756, in4756_1, in4756_2;
    wire c4756;
    assign in4756_1 = {pp99[78]};
    assign in4756_2 = {pp100[77]};
    Full_Adder FA_4756(s4756, c4756, in4756_1, in4756_2, pp98[79]);
    wire[0:0] s4757, in4757_1, in4757_2;
    wire c4757;
    assign in4757_1 = {pp102[75]};
    assign in4757_2 = {pp103[74]};
    Full_Adder FA_4757(s4757, c4757, in4757_1, in4757_2, pp101[76]);
    wire[0:0] s4758, in4758_1, in4758_2;
    wire c4758;
    assign in4758_1 = {pp105[72]};
    assign in4758_2 = {pp106[71]};
    Full_Adder FA_4758(s4758, c4758, in4758_1, in4758_2, pp104[73]);
    wire[0:0] s4759, in4759_1, in4759_2;
    wire c4759;
    assign in4759_1 = {pp108[69]};
    assign in4759_2 = {pp109[68]};
    Full_Adder FA_4759(s4759, c4759, in4759_1, in4759_2, pp107[70]);
    wire[0:0] s4760, in4760_1, in4760_2;
    wire c4760;
    assign in4760_1 = {pp111[66]};
    assign in4760_2 = {pp112[65]};
    Full_Adder FA_4760(s4760, c4760, in4760_1, in4760_2, pp110[67]);
    wire[0:0] s4761, in4761_1, in4761_2;
    wire c4761;
    assign in4761_1 = {pp52[126]};
    assign in4761_2 = {pp53[125]};
    Full_Adder FA_4761(s4761, c4761, in4761_1, in4761_2, pp51[127]);
    wire[0:0] s4762, in4762_1, in4762_2;
    wire c4762;
    assign in4762_1 = {pp55[123]};
    assign in4762_2 = {pp56[122]};
    Full_Adder FA_4762(s4762, c4762, in4762_1, in4762_2, pp54[124]);
    wire[0:0] s4763, in4763_1, in4763_2;
    wire c4763;
    assign in4763_1 = {pp58[120]};
    assign in4763_2 = {pp59[119]};
    Full_Adder FA_4763(s4763, c4763, in4763_1, in4763_2, pp57[121]);
    wire[0:0] s4764, in4764_1, in4764_2;
    wire c4764;
    assign in4764_1 = {pp61[117]};
    assign in4764_2 = {pp62[116]};
    Full_Adder FA_4764(s4764, c4764, in4764_1, in4764_2, pp60[118]);
    wire[0:0] s4765, in4765_1, in4765_2;
    wire c4765;
    assign in4765_1 = {pp64[114]};
    assign in4765_2 = {pp65[113]};
    Full_Adder FA_4765(s4765, c4765, in4765_1, in4765_2, pp63[115]);
    wire[0:0] s4766, in4766_1, in4766_2;
    wire c4766;
    assign in4766_1 = {pp67[111]};
    assign in4766_2 = {pp68[110]};
    Full_Adder FA_4766(s4766, c4766, in4766_1, in4766_2, pp66[112]);
    wire[0:0] s4767, in4767_1, in4767_2;
    wire c4767;
    assign in4767_1 = {pp70[108]};
    assign in4767_2 = {pp71[107]};
    Full_Adder FA_4767(s4767, c4767, in4767_1, in4767_2, pp69[109]);
    wire[0:0] s4768, in4768_1, in4768_2;
    wire c4768;
    assign in4768_1 = {pp73[105]};
    assign in4768_2 = {pp74[104]};
    Full_Adder FA_4768(s4768, c4768, in4768_1, in4768_2, pp72[106]);
    wire[0:0] s4769, in4769_1, in4769_2;
    wire c4769;
    assign in4769_1 = {pp76[102]};
    assign in4769_2 = {pp77[101]};
    Full_Adder FA_4769(s4769, c4769, in4769_1, in4769_2, pp75[103]);
    wire[0:0] s4770, in4770_1, in4770_2;
    wire c4770;
    assign in4770_1 = {pp79[99]};
    assign in4770_2 = {pp80[98]};
    Full_Adder FA_4770(s4770, c4770, in4770_1, in4770_2, pp78[100]);
    wire[0:0] s4771, in4771_1, in4771_2;
    wire c4771;
    assign in4771_1 = {pp82[96]};
    assign in4771_2 = {pp83[95]};
    Full_Adder FA_4771(s4771, c4771, in4771_1, in4771_2, pp81[97]);
    wire[0:0] s4772, in4772_1, in4772_2;
    wire c4772;
    assign in4772_1 = {pp85[93]};
    assign in4772_2 = {pp86[92]};
    Full_Adder FA_4772(s4772, c4772, in4772_1, in4772_2, pp84[94]);
    wire[0:0] s4773, in4773_1, in4773_2;
    wire c4773;
    assign in4773_1 = {pp88[90]};
    assign in4773_2 = {pp89[89]};
    Full_Adder FA_4773(s4773, c4773, in4773_1, in4773_2, pp87[91]);
    wire[0:0] s4774, in4774_1, in4774_2;
    wire c4774;
    assign in4774_1 = {pp91[87]};
    assign in4774_2 = {pp92[86]};
    Full_Adder FA_4774(s4774, c4774, in4774_1, in4774_2, pp90[88]);
    wire[0:0] s4775, in4775_1, in4775_2;
    wire c4775;
    assign in4775_1 = {pp94[84]};
    assign in4775_2 = {pp95[83]};
    Full_Adder FA_4775(s4775, c4775, in4775_1, in4775_2, pp93[85]);
    wire[0:0] s4776, in4776_1, in4776_2;
    wire c4776;
    assign in4776_1 = {pp97[81]};
    assign in4776_2 = {pp98[80]};
    Full_Adder FA_4776(s4776, c4776, in4776_1, in4776_2, pp96[82]);
    wire[0:0] s4777, in4777_1, in4777_2;
    wire c4777;
    assign in4777_1 = {pp100[78]};
    assign in4777_2 = {pp101[77]};
    Full_Adder FA_4777(s4777, c4777, in4777_1, in4777_2, pp99[79]);
    wire[0:0] s4778, in4778_1, in4778_2;
    wire c4778;
    assign in4778_1 = {pp103[75]};
    assign in4778_2 = {pp104[74]};
    Full_Adder FA_4778(s4778, c4778, in4778_1, in4778_2, pp102[76]);
    wire[0:0] s4779, in4779_1, in4779_2;
    wire c4779;
    assign in4779_1 = {pp106[72]};
    assign in4779_2 = {pp107[71]};
    Full_Adder FA_4779(s4779, c4779, in4779_1, in4779_2, pp105[73]);
    wire[0:0] s4780, in4780_1, in4780_2;
    wire c4780;
    assign in4780_1 = {pp109[69]};
    assign in4780_2 = {pp110[68]};
    Full_Adder FA_4780(s4780, c4780, in4780_1, in4780_2, pp108[70]);
    wire[0:0] s4781, in4781_1, in4781_2;
    wire c4781;
    assign in4781_1 = {pp53[126]};
    assign in4781_2 = {pp54[125]};
    Full_Adder FA_4781(s4781, c4781, in4781_1, in4781_2, pp52[127]);
    wire[0:0] s4782, in4782_1, in4782_2;
    wire c4782;
    assign in4782_1 = {pp56[123]};
    assign in4782_2 = {pp57[122]};
    Full_Adder FA_4782(s4782, c4782, in4782_1, in4782_2, pp55[124]);
    wire[0:0] s4783, in4783_1, in4783_2;
    wire c4783;
    assign in4783_1 = {pp59[120]};
    assign in4783_2 = {pp60[119]};
    Full_Adder FA_4783(s4783, c4783, in4783_1, in4783_2, pp58[121]);
    wire[0:0] s4784, in4784_1, in4784_2;
    wire c4784;
    assign in4784_1 = {pp62[117]};
    assign in4784_2 = {pp63[116]};
    Full_Adder FA_4784(s4784, c4784, in4784_1, in4784_2, pp61[118]);
    wire[0:0] s4785, in4785_1, in4785_2;
    wire c4785;
    assign in4785_1 = {pp65[114]};
    assign in4785_2 = {pp66[113]};
    Full_Adder FA_4785(s4785, c4785, in4785_1, in4785_2, pp64[115]);
    wire[0:0] s4786, in4786_1, in4786_2;
    wire c4786;
    assign in4786_1 = {pp68[111]};
    assign in4786_2 = {pp69[110]};
    Full_Adder FA_4786(s4786, c4786, in4786_1, in4786_2, pp67[112]);
    wire[0:0] s4787, in4787_1, in4787_2;
    wire c4787;
    assign in4787_1 = {pp71[108]};
    assign in4787_2 = {pp72[107]};
    Full_Adder FA_4787(s4787, c4787, in4787_1, in4787_2, pp70[109]);
    wire[0:0] s4788, in4788_1, in4788_2;
    wire c4788;
    assign in4788_1 = {pp74[105]};
    assign in4788_2 = {pp75[104]};
    Full_Adder FA_4788(s4788, c4788, in4788_1, in4788_2, pp73[106]);
    wire[0:0] s4789, in4789_1, in4789_2;
    wire c4789;
    assign in4789_1 = {pp77[102]};
    assign in4789_2 = {pp78[101]};
    Full_Adder FA_4789(s4789, c4789, in4789_1, in4789_2, pp76[103]);
    wire[0:0] s4790, in4790_1, in4790_2;
    wire c4790;
    assign in4790_1 = {pp80[99]};
    assign in4790_2 = {pp81[98]};
    Full_Adder FA_4790(s4790, c4790, in4790_1, in4790_2, pp79[100]);
    wire[0:0] s4791, in4791_1, in4791_2;
    wire c4791;
    assign in4791_1 = {pp83[96]};
    assign in4791_2 = {pp84[95]};
    Full_Adder FA_4791(s4791, c4791, in4791_1, in4791_2, pp82[97]);
    wire[0:0] s4792, in4792_1, in4792_2;
    wire c4792;
    assign in4792_1 = {pp86[93]};
    assign in4792_2 = {pp87[92]};
    Full_Adder FA_4792(s4792, c4792, in4792_1, in4792_2, pp85[94]);
    wire[0:0] s4793, in4793_1, in4793_2;
    wire c4793;
    assign in4793_1 = {pp89[90]};
    assign in4793_2 = {pp90[89]};
    Full_Adder FA_4793(s4793, c4793, in4793_1, in4793_2, pp88[91]);
    wire[0:0] s4794, in4794_1, in4794_2;
    wire c4794;
    assign in4794_1 = {pp92[87]};
    assign in4794_2 = {pp93[86]};
    Full_Adder FA_4794(s4794, c4794, in4794_1, in4794_2, pp91[88]);
    wire[0:0] s4795, in4795_1, in4795_2;
    wire c4795;
    assign in4795_1 = {pp95[84]};
    assign in4795_2 = {pp96[83]};
    Full_Adder FA_4795(s4795, c4795, in4795_1, in4795_2, pp94[85]);
    wire[0:0] s4796, in4796_1, in4796_2;
    wire c4796;
    assign in4796_1 = {pp98[81]};
    assign in4796_2 = {pp99[80]};
    Full_Adder FA_4796(s4796, c4796, in4796_1, in4796_2, pp97[82]);
    wire[0:0] s4797, in4797_1, in4797_2;
    wire c4797;
    assign in4797_1 = {pp101[78]};
    assign in4797_2 = {pp102[77]};
    Full_Adder FA_4797(s4797, c4797, in4797_1, in4797_2, pp100[79]);
    wire[0:0] s4798, in4798_1, in4798_2;
    wire c4798;
    assign in4798_1 = {pp104[75]};
    assign in4798_2 = {pp105[74]};
    Full_Adder FA_4798(s4798, c4798, in4798_1, in4798_2, pp103[76]);
    wire[0:0] s4799, in4799_1, in4799_2;
    wire c4799;
    assign in4799_1 = {pp107[72]};
    assign in4799_2 = {pp108[71]};
    Full_Adder FA_4799(s4799, c4799, in4799_1, in4799_2, pp106[73]);
    wire[0:0] s4800, in4800_1, in4800_2;
    wire c4800;
    assign in4800_1 = {pp54[126]};
    assign in4800_2 = {pp55[125]};
    Full_Adder FA_4800(s4800, c4800, in4800_1, in4800_2, pp53[127]);
    wire[0:0] s4801, in4801_1, in4801_2;
    wire c4801;
    assign in4801_1 = {pp57[123]};
    assign in4801_2 = {pp58[122]};
    Full_Adder FA_4801(s4801, c4801, in4801_1, in4801_2, pp56[124]);
    wire[0:0] s4802, in4802_1, in4802_2;
    wire c4802;
    assign in4802_1 = {pp60[120]};
    assign in4802_2 = {pp61[119]};
    Full_Adder FA_4802(s4802, c4802, in4802_1, in4802_2, pp59[121]);
    wire[0:0] s4803, in4803_1, in4803_2;
    wire c4803;
    assign in4803_1 = {pp63[117]};
    assign in4803_2 = {pp64[116]};
    Full_Adder FA_4803(s4803, c4803, in4803_1, in4803_2, pp62[118]);
    wire[0:0] s4804, in4804_1, in4804_2;
    wire c4804;
    assign in4804_1 = {pp66[114]};
    assign in4804_2 = {pp67[113]};
    Full_Adder FA_4804(s4804, c4804, in4804_1, in4804_2, pp65[115]);
    wire[0:0] s4805, in4805_1, in4805_2;
    wire c4805;
    assign in4805_1 = {pp69[111]};
    assign in4805_2 = {pp70[110]};
    Full_Adder FA_4805(s4805, c4805, in4805_1, in4805_2, pp68[112]);
    wire[0:0] s4806, in4806_1, in4806_2;
    wire c4806;
    assign in4806_1 = {pp72[108]};
    assign in4806_2 = {pp73[107]};
    Full_Adder FA_4806(s4806, c4806, in4806_1, in4806_2, pp71[109]);
    wire[0:0] s4807, in4807_1, in4807_2;
    wire c4807;
    assign in4807_1 = {pp75[105]};
    assign in4807_2 = {pp76[104]};
    Full_Adder FA_4807(s4807, c4807, in4807_1, in4807_2, pp74[106]);
    wire[0:0] s4808, in4808_1, in4808_2;
    wire c4808;
    assign in4808_1 = {pp78[102]};
    assign in4808_2 = {pp79[101]};
    Full_Adder FA_4808(s4808, c4808, in4808_1, in4808_2, pp77[103]);
    wire[0:0] s4809, in4809_1, in4809_2;
    wire c4809;
    assign in4809_1 = {pp81[99]};
    assign in4809_2 = {pp82[98]};
    Full_Adder FA_4809(s4809, c4809, in4809_1, in4809_2, pp80[100]);
    wire[0:0] s4810, in4810_1, in4810_2;
    wire c4810;
    assign in4810_1 = {pp84[96]};
    assign in4810_2 = {pp85[95]};
    Full_Adder FA_4810(s4810, c4810, in4810_1, in4810_2, pp83[97]);
    wire[0:0] s4811, in4811_1, in4811_2;
    wire c4811;
    assign in4811_1 = {pp87[93]};
    assign in4811_2 = {pp88[92]};
    Full_Adder FA_4811(s4811, c4811, in4811_1, in4811_2, pp86[94]);
    wire[0:0] s4812, in4812_1, in4812_2;
    wire c4812;
    assign in4812_1 = {pp90[90]};
    assign in4812_2 = {pp91[89]};
    Full_Adder FA_4812(s4812, c4812, in4812_1, in4812_2, pp89[91]);
    wire[0:0] s4813, in4813_1, in4813_2;
    wire c4813;
    assign in4813_1 = {pp93[87]};
    assign in4813_2 = {pp94[86]};
    Full_Adder FA_4813(s4813, c4813, in4813_1, in4813_2, pp92[88]);
    wire[0:0] s4814, in4814_1, in4814_2;
    wire c4814;
    assign in4814_1 = {pp96[84]};
    assign in4814_2 = {pp97[83]};
    Full_Adder FA_4814(s4814, c4814, in4814_1, in4814_2, pp95[85]);
    wire[0:0] s4815, in4815_1, in4815_2;
    wire c4815;
    assign in4815_1 = {pp99[81]};
    assign in4815_2 = {pp100[80]};
    Full_Adder FA_4815(s4815, c4815, in4815_1, in4815_2, pp98[82]);
    wire[0:0] s4816, in4816_1, in4816_2;
    wire c4816;
    assign in4816_1 = {pp102[78]};
    assign in4816_2 = {pp103[77]};
    Full_Adder FA_4816(s4816, c4816, in4816_1, in4816_2, pp101[79]);
    wire[0:0] s4817, in4817_1, in4817_2;
    wire c4817;
    assign in4817_1 = {pp105[75]};
    assign in4817_2 = {pp106[74]};
    Full_Adder FA_4817(s4817, c4817, in4817_1, in4817_2, pp104[76]);
    wire[0:0] s4818, in4818_1, in4818_2;
    wire c4818;
    assign in4818_1 = {pp55[126]};
    assign in4818_2 = {pp56[125]};
    Full_Adder FA_4818(s4818, c4818, in4818_1, in4818_2, pp54[127]);
    wire[0:0] s4819, in4819_1, in4819_2;
    wire c4819;
    assign in4819_1 = {pp58[123]};
    assign in4819_2 = {pp59[122]};
    Full_Adder FA_4819(s4819, c4819, in4819_1, in4819_2, pp57[124]);
    wire[0:0] s4820, in4820_1, in4820_2;
    wire c4820;
    assign in4820_1 = {pp61[120]};
    assign in4820_2 = {pp62[119]};
    Full_Adder FA_4820(s4820, c4820, in4820_1, in4820_2, pp60[121]);
    wire[0:0] s4821, in4821_1, in4821_2;
    wire c4821;
    assign in4821_1 = {pp64[117]};
    assign in4821_2 = {pp65[116]};
    Full_Adder FA_4821(s4821, c4821, in4821_1, in4821_2, pp63[118]);
    wire[0:0] s4822, in4822_1, in4822_2;
    wire c4822;
    assign in4822_1 = {pp67[114]};
    assign in4822_2 = {pp68[113]};
    Full_Adder FA_4822(s4822, c4822, in4822_1, in4822_2, pp66[115]);
    wire[0:0] s4823, in4823_1, in4823_2;
    wire c4823;
    assign in4823_1 = {pp70[111]};
    assign in4823_2 = {pp71[110]};
    Full_Adder FA_4823(s4823, c4823, in4823_1, in4823_2, pp69[112]);
    wire[0:0] s4824, in4824_1, in4824_2;
    wire c4824;
    assign in4824_1 = {pp73[108]};
    assign in4824_2 = {pp74[107]};
    Full_Adder FA_4824(s4824, c4824, in4824_1, in4824_2, pp72[109]);
    wire[0:0] s4825, in4825_1, in4825_2;
    wire c4825;
    assign in4825_1 = {pp76[105]};
    assign in4825_2 = {pp77[104]};
    Full_Adder FA_4825(s4825, c4825, in4825_1, in4825_2, pp75[106]);
    wire[0:0] s4826, in4826_1, in4826_2;
    wire c4826;
    assign in4826_1 = {pp79[102]};
    assign in4826_2 = {pp80[101]};
    Full_Adder FA_4826(s4826, c4826, in4826_1, in4826_2, pp78[103]);
    wire[0:0] s4827, in4827_1, in4827_2;
    wire c4827;
    assign in4827_1 = {pp82[99]};
    assign in4827_2 = {pp83[98]};
    Full_Adder FA_4827(s4827, c4827, in4827_1, in4827_2, pp81[100]);
    wire[0:0] s4828, in4828_1, in4828_2;
    wire c4828;
    assign in4828_1 = {pp85[96]};
    assign in4828_2 = {pp86[95]};
    Full_Adder FA_4828(s4828, c4828, in4828_1, in4828_2, pp84[97]);
    wire[0:0] s4829, in4829_1, in4829_2;
    wire c4829;
    assign in4829_1 = {pp88[93]};
    assign in4829_2 = {pp89[92]};
    Full_Adder FA_4829(s4829, c4829, in4829_1, in4829_2, pp87[94]);
    wire[0:0] s4830, in4830_1, in4830_2;
    wire c4830;
    assign in4830_1 = {pp91[90]};
    assign in4830_2 = {pp92[89]};
    Full_Adder FA_4830(s4830, c4830, in4830_1, in4830_2, pp90[91]);
    wire[0:0] s4831, in4831_1, in4831_2;
    wire c4831;
    assign in4831_1 = {pp94[87]};
    assign in4831_2 = {pp95[86]};
    Full_Adder FA_4831(s4831, c4831, in4831_1, in4831_2, pp93[88]);
    wire[0:0] s4832, in4832_1, in4832_2;
    wire c4832;
    assign in4832_1 = {pp97[84]};
    assign in4832_2 = {pp98[83]};
    Full_Adder FA_4832(s4832, c4832, in4832_1, in4832_2, pp96[85]);
    wire[0:0] s4833, in4833_1, in4833_2;
    wire c4833;
    assign in4833_1 = {pp100[81]};
    assign in4833_2 = {pp101[80]};
    Full_Adder FA_4833(s4833, c4833, in4833_1, in4833_2, pp99[82]);
    wire[0:0] s4834, in4834_1, in4834_2;
    wire c4834;
    assign in4834_1 = {pp103[78]};
    assign in4834_2 = {pp104[77]};
    Full_Adder FA_4834(s4834, c4834, in4834_1, in4834_2, pp102[79]);
    wire[0:0] s4835, in4835_1, in4835_2;
    wire c4835;
    assign in4835_1 = {pp56[126]};
    assign in4835_2 = {pp57[125]};
    Full_Adder FA_4835(s4835, c4835, in4835_1, in4835_2, pp55[127]);
    wire[0:0] s4836, in4836_1, in4836_2;
    wire c4836;
    assign in4836_1 = {pp59[123]};
    assign in4836_2 = {pp60[122]};
    Full_Adder FA_4836(s4836, c4836, in4836_1, in4836_2, pp58[124]);
    wire[0:0] s4837, in4837_1, in4837_2;
    wire c4837;
    assign in4837_1 = {pp62[120]};
    assign in4837_2 = {pp63[119]};
    Full_Adder FA_4837(s4837, c4837, in4837_1, in4837_2, pp61[121]);
    wire[0:0] s4838, in4838_1, in4838_2;
    wire c4838;
    assign in4838_1 = {pp65[117]};
    assign in4838_2 = {pp66[116]};
    Full_Adder FA_4838(s4838, c4838, in4838_1, in4838_2, pp64[118]);
    wire[0:0] s4839, in4839_1, in4839_2;
    wire c4839;
    assign in4839_1 = {pp68[114]};
    assign in4839_2 = {pp69[113]};
    Full_Adder FA_4839(s4839, c4839, in4839_1, in4839_2, pp67[115]);
    wire[0:0] s4840, in4840_1, in4840_2;
    wire c4840;
    assign in4840_1 = {pp71[111]};
    assign in4840_2 = {pp72[110]};
    Full_Adder FA_4840(s4840, c4840, in4840_1, in4840_2, pp70[112]);
    wire[0:0] s4841, in4841_1, in4841_2;
    wire c4841;
    assign in4841_1 = {pp74[108]};
    assign in4841_2 = {pp75[107]};
    Full_Adder FA_4841(s4841, c4841, in4841_1, in4841_2, pp73[109]);
    wire[0:0] s4842, in4842_1, in4842_2;
    wire c4842;
    assign in4842_1 = {pp77[105]};
    assign in4842_2 = {pp78[104]};
    Full_Adder FA_4842(s4842, c4842, in4842_1, in4842_2, pp76[106]);
    wire[0:0] s4843, in4843_1, in4843_2;
    wire c4843;
    assign in4843_1 = {pp80[102]};
    assign in4843_2 = {pp81[101]};
    Full_Adder FA_4843(s4843, c4843, in4843_1, in4843_2, pp79[103]);
    wire[0:0] s4844, in4844_1, in4844_2;
    wire c4844;
    assign in4844_1 = {pp83[99]};
    assign in4844_2 = {pp84[98]};
    Full_Adder FA_4844(s4844, c4844, in4844_1, in4844_2, pp82[100]);
    wire[0:0] s4845, in4845_1, in4845_2;
    wire c4845;
    assign in4845_1 = {pp86[96]};
    assign in4845_2 = {pp87[95]};
    Full_Adder FA_4845(s4845, c4845, in4845_1, in4845_2, pp85[97]);
    wire[0:0] s4846, in4846_1, in4846_2;
    wire c4846;
    assign in4846_1 = {pp89[93]};
    assign in4846_2 = {pp90[92]};
    Full_Adder FA_4846(s4846, c4846, in4846_1, in4846_2, pp88[94]);
    wire[0:0] s4847, in4847_1, in4847_2;
    wire c4847;
    assign in4847_1 = {pp92[90]};
    assign in4847_2 = {pp93[89]};
    Full_Adder FA_4847(s4847, c4847, in4847_1, in4847_2, pp91[91]);
    wire[0:0] s4848, in4848_1, in4848_2;
    wire c4848;
    assign in4848_1 = {pp95[87]};
    assign in4848_2 = {pp96[86]};
    Full_Adder FA_4848(s4848, c4848, in4848_1, in4848_2, pp94[88]);
    wire[0:0] s4849, in4849_1, in4849_2;
    wire c4849;
    assign in4849_1 = {pp98[84]};
    assign in4849_2 = {pp99[83]};
    Full_Adder FA_4849(s4849, c4849, in4849_1, in4849_2, pp97[85]);
    wire[0:0] s4850, in4850_1, in4850_2;
    wire c4850;
    assign in4850_1 = {pp101[81]};
    assign in4850_2 = {pp102[80]};
    Full_Adder FA_4850(s4850, c4850, in4850_1, in4850_2, pp100[82]);
    wire[0:0] s4851, in4851_1, in4851_2;
    wire c4851;
    assign in4851_1 = {pp57[126]};
    assign in4851_2 = {pp58[125]};
    Full_Adder FA_4851(s4851, c4851, in4851_1, in4851_2, pp56[127]);
    wire[0:0] s4852, in4852_1, in4852_2;
    wire c4852;
    assign in4852_1 = {pp60[123]};
    assign in4852_2 = {pp61[122]};
    Full_Adder FA_4852(s4852, c4852, in4852_1, in4852_2, pp59[124]);
    wire[0:0] s4853, in4853_1, in4853_2;
    wire c4853;
    assign in4853_1 = {pp63[120]};
    assign in4853_2 = {pp64[119]};
    Full_Adder FA_4853(s4853, c4853, in4853_1, in4853_2, pp62[121]);
    wire[0:0] s4854, in4854_1, in4854_2;
    wire c4854;
    assign in4854_1 = {pp66[117]};
    assign in4854_2 = {pp67[116]};
    Full_Adder FA_4854(s4854, c4854, in4854_1, in4854_2, pp65[118]);
    wire[0:0] s4855, in4855_1, in4855_2;
    wire c4855;
    assign in4855_1 = {pp69[114]};
    assign in4855_2 = {pp70[113]};
    Full_Adder FA_4855(s4855, c4855, in4855_1, in4855_2, pp68[115]);
    wire[0:0] s4856, in4856_1, in4856_2;
    wire c4856;
    assign in4856_1 = {pp72[111]};
    assign in4856_2 = {pp73[110]};
    Full_Adder FA_4856(s4856, c4856, in4856_1, in4856_2, pp71[112]);
    wire[0:0] s4857, in4857_1, in4857_2;
    wire c4857;
    assign in4857_1 = {pp75[108]};
    assign in4857_2 = {pp76[107]};
    Full_Adder FA_4857(s4857, c4857, in4857_1, in4857_2, pp74[109]);
    wire[0:0] s4858, in4858_1, in4858_2;
    wire c4858;
    assign in4858_1 = {pp78[105]};
    assign in4858_2 = {pp79[104]};
    Full_Adder FA_4858(s4858, c4858, in4858_1, in4858_2, pp77[106]);
    wire[0:0] s4859, in4859_1, in4859_2;
    wire c4859;
    assign in4859_1 = {pp81[102]};
    assign in4859_2 = {pp82[101]};
    Full_Adder FA_4859(s4859, c4859, in4859_1, in4859_2, pp80[103]);
    wire[0:0] s4860, in4860_1, in4860_2;
    wire c4860;
    assign in4860_1 = {pp84[99]};
    assign in4860_2 = {pp85[98]};
    Full_Adder FA_4860(s4860, c4860, in4860_1, in4860_2, pp83[100]);
    wire[0:0] s4861, in4861_1, in4861_2;
    wire c4861;
    assign in4861_1 = {pp87[96]};
    assign in4861_2 = {pp88[95]};
    Full_Adder FA_4861(s4861, c4861, in4861_1, in4861_2, pp86[97]);
    wire[0:0] s4862, in4862_1, in4862_2;
    wire c4862;
    assign in4862_1 = {pp90[93]};
    assign in4862_2 = {pp91[92]};
    Full_Adder FA_4862(s4862, c4862, in4862_1, in4862_2, pp89[94]);
    wire[0:0] s4863, in4863_1, in4863_2;
    wire c4863;
    assign in4863_1 = {pp93[90]};
    assign in4863_2 = {pp94[89]};
    Full_Adder FA_4863(s4863, c4863, in4863_1, in4863_2, pp92[91]);
    wire[0:0] s4864, in4864_1, in4864_2;
    wire c4864;
    assign in4864_1 = {pp96[87]};
    assign in4864_2 = {pp97[86]};
    Full_Adder FA_4864(s4864, c4864, in4864_1, in4864_2, pp95[88]);
    wire[0:0] s4865, in4865_1, in4865_2;
    wire c4865;
    assign in4865_1 = {pp99[84]};
    assign in4865_2 = {pp100[83]};
    Full_Adder FA_4865(s4865, c4865, in4865_1, in4865_2, pp98[85]);
    wire[0:0] s4866, in4866_1, in4866_2;
    wire c4866;
    assign in4866_1 = {pp58[126]};
    assign in4866_2 = {pp59[125]};
    Full_Adder FA_4866(s4866, c4866, in4866_1, in4866_2, pp57[127]);
    wire[0:0] s4867, in4867_1, in4867_2;
    wire c4867;
    assign in4867_1 = {pp61[123]};
    assign in4867_2 = {pp62[122]};
    Full_Adder FA_4867(s4867, c4867, in4867_1, in4867_2, pp60[124]);
    wire[0:0] s4868, in4868_1, in4868_2;
    wire c4868;
    assign in4868_1 = {pp64[120]};
    assign in4868_2 = {pp65[119]};
    Full_Adder FA_4868(s4868, c4868, in4868_1, in4868_2, pp63[121]);
    wire[0:0] s4869, in4869_1, in4869_2;
    wire c4869;
    assign in4869_1 = {pp67[117]};
    assign in4869_2 = {pp68[116]};
    Full_Adder FA_4869(s4869, c4869, in4869_1, in4869_2, pp66[118]);
    wire[0:0] s4870, in4870_1, in4870_2;
    wire c4870;
    assign in4870_1 = {pp70[114]};
    assign in4870_2 = {pp71[113]};
    Full_Adder FA_4870(s4870, c4870, in4870_1, in4870_2, pp69[115]);
    wire[0:0] s4871, in4871_1, in4871_2;
    wire c4871;
    assign in4871_1 = {pp73[111]};
    assign in4871_2 = {pp74[110]};
    Full_Adder FA_4871(s4871, c4871, in4871_1, in4871_2, pp72[112]);
    wire[0:0] s4872, in4872_1, in4872_2;
    wire c4872;
    assign in4872_1 = {pp76[108]};
    assign in4872_2 = {pp77[107]};
    Full_Adder FA_4872(s4872, c4872, in4872_1, in4872_2, pp75[109]);
    wire[0:0] s4873, in4873_1, in4873_2;
    wire c4873;
    assign in4873_1 = {pp79[105]};
    assign in4873_2 = {pp80[104]};
    Full_Adder FA_4873(s4873, c4873, in4873_1, in4873_2, pp78[106]);
    wire[0:0] s4874, in4874_1, in4874_2;
    wire c4874;
    assign in4874_1 = {pp82[102]};
    assign in4874_2 = {pp83[101]};
    Full_Adder FA_4874(s4874, c4874, in4874_1, in4874_2, pp81[103]);
    wire[0:0] s4875, in4875_1, in4875_2;
    wire c4875;
    assign in4875_1 = {pp85[99]};
    assign in4875_2 = {pp86[98]};
    Full_Adder FA_4875(s4875, c4875, in4875_1, in4875_2, pp84[100]);
    wire[0:0] s4876, in4876_1, in4876_2;
    wire c4876;
    assign in4876_1 = {pp88[96]};
    assign in4876_2 = {pp89[95]};
    Full_Adder FA_4876(s4876, c4876, in4876_1, in4876_2, pp87[97]);
    wire[0:0] s4877, in4877_1, in4877_2;
    wire c4877;
    assign in4877_1 = {pp91[93]};
    assign in4877_2 = {pp92[92]};
    Full_Adder FA_4877(s4877, c4877, in4877_1, in4877_2, pp90[94]);
    wire[0:0] s4878, in4878_1, in4878_2;
    wire c4878;
    assign in4878_1 = {pp94[90]};
    assign in4878_2 = {pp95[89]};
    Full_Adder FA_4878(s4878, c4878, in4878_1, in4878_2, pp93[91]);
    wire[0:0] s4879, in4879_1, in4879_2;
    wire c4879;
    assign in4879_1 = {pp97[87]};
    assign in4879_2 = {pp98[86]};
    Full_Adder FA_4879(s4879, c4879, in4879_1, in4879_2, pp96[88]);
    wire[0:0] s4880, in4880_1, in4880_2;
    wire c4880;
    assign in4880_1 = {pp59[126]};
    assign in4880_2 = {pp60[125]};
    Full_Adder FA_4880(s4880, c4880, in4880_1, in4880_2, pp58[127]);
    wire[0:0] s4881, in4881_1, in4881_2;
    wire c4881;
    assign in4881_1 = {pp62[123]};
    assign in4881_2 = {pp63[122]};
    Full_Adder FA_4881(s4881, c4881, in4881_1, in4881_2, pp61[124]);
    wire[0:0] s4882, in4882_1, in4882_2;
    wire c4882;
    assign in4882_1 = {pp65[120]};
    assign in4882_2 = {pp66[119]};
    Full_Adder FA_4882(s4882, c4882, in4882_1, in4882_2, pp64[121]);
    wire[0:0] s4883, in4883_1, in4883_2;
    wire c4883;
    assign in4883_1 = {pp68[117]};
    assign in4883_2 = {pp69[116]};
    Full_Adder FA_4883(s4883, c4883, in4883_1, in4883_2, pp67[118]);
    wire[0:0] s4884, in4884_1, in4884_2;
    wire c4884;
    assign in4884_1 = {pp71[114]};
    assign in4884_2 = {pp72[113]};
    Full_Adder FA_4884(s4884, c4884, in4884_1, in4884_2, pp70[115]);
    wire[0:0] s4885, in4885_1, in4885_2;
    wire c4885;
    assign in4885_1 = {pp74[111]};
    assign in4885_2 = {pp75[110]};
    Full_Adder FA_4885(s4885, c4885, in4885_1, in4885_2, pp73[112]);
    wire[0:0] s4886, in4886_1, in4886_2;
    wire c4886;
    assign in4886_1 = {pp77[108]};
    assign in4886_2 = {pp78[107]};
    Full_Adder FA_4886(s4886, c4886, in4886_1, in4886_2, pp76[109]);
    wire[0:0] s4887, in4887_1, in4887_2;
    wire c4887;
    assign in4887_1 = {pp80[105]};
    assign in4887_2 = {pp81[104]};
    Full_Adder FA_4887(s4887, c4887, in4887_1, in4887_2, pp79[106]);
    wire[0:0] s4888, in4888_1, in4888_2;
    wire c4888;
    assign in4888_1 = {pp83[102]};
    assign in4888_2 = {pp84[101]};
    Full_Adder FA_4888(s4888, c4888, in4888_1, in4888_2, pp82[103]);
    wire[0:0] s4889, in4889_1, in4889_2;
    wire c4889;
    assign in4889_1 = {pp86[99]};
    assign in4889_2 = {pp87[98]};
    Full_Adder FA_4889(s4889, c4889, in4889_1, in4889_2, pp85[100]);
    wire[0:0] s4890, in4890_1, in4890_2;
    wire c4890;
    assign in4890_1 = {pp89[96]};
    assign in4890_2 = {pp90[95]};
    Full_Adder FA_4890(s4890, c4890, in4890_1, in4890_2, pp88[97]);
    wire[0:0] s4891, in4891_1, in4891_2;
    wire c4891;
    assign in4891_1 = {pp92[93]};
    assign in4891_2 = {pp93[92]};
    Full_Adder FA_4891(s4891, c4891, in4891_1, in4891_2, pp91[94]);
    wire[0:0] s4892, in4892_1, in4892_2;
    wire c4892;
    assign in4892_1 = {pp95[90]};
    assign in4892_2 = {pp96[89]};
    Full_Adder FA_4892(s4892, c4892, in4892_1, in4892_2, pp94[91]);
    wire[0:0] s4893, in4893_1, in4893_2;
    wire c4893;
    assign in4893_1 = {pp60[126]};
    assign in4893_2 = {pp61[125]};
    Full_Adder FA_4893(s4893, c4893, in4893_1, in4893_2, pp59[127]);
    wire[0:0] s4894, in4894_1, in4894_2;
    wire c4894;
    assign in4894_1 = {pp63[123]};
    assign in4894_2 = {pp64[122]};
    Full_Adder FA_4894(s4894, c4894, in4894_1, in4894_2, pp62[124]);
    wire[0:0] s4895, in4895_1, in4895_2;
    wire c4895;
    assign in4895_1 = {pp66[120]};
    assign in4895_2 = {pp67[119]};
    Full_Adder FA_4895(s4895, c4895, in4895_1, in4895_2, pp65[121]);
    wire[0:0] s4896, in4896_1, in4896_2;
    wire c4896;
    assign in4896_1 = {pp69[117]};
    assign in4896_2 = {pp70[116]};
    Full_Adder FA_4896(s4896, c4896, in4896_1, in4896_2, pp68[118]);
    wire[0:0] s4897, in4897_1, in4897_2;
    wire c4897;
    assign in4897_1 = {pp72[114]};
    assign in4897_2 = {pp73[113]};
    Full_Adder FA_4897(s4897, c4897, in4897_1, in4897_2, pp71[115]);
    wire[0:0] s4898, in4898_1, in4898_2;
    wire c4898;
    assign in4898_1 = {pp75[111]};
    assign in4898_2 = {pp76[110]};
    Full_Adder FA_4898(s4898, c4898, in4898_1, in4898_2, pp74[112]);
    wire[0:0] s4899, in4899_1, in4899_2;
    wire c4899;
    assign in4899_1 = {pp78[108]};
    assign in4899_2 = {pp79[107]};
    Full_Adder FA_4899(s4899, c4899, in4899_1, in4899_2, pp77[109]);
    wire[0:0] s4900, in4900_1, in4900_2;
    wire c4900;
    assign in4900_1 = {pp81[105]};
    assign in4900_2 = {pp82[104]};
    Full_Adder FA_4900(s4900, c4900, in4900_1, in4900_2, pp80[106]);
    wire[0:0] s4901, in4901_1, in4901_2;
    wire c4901;
    assign in4901_1 = {pp84[102]};
    assign in4901_2 = {pp85[101]};
    Full_Adder FA_4901(s4901, c4901, in4901_1, in4901_2, pp83[103]);
    wire[0:0] s4902, in4902_1, in4902_2;
    wire c4902;
    assign in4902_1 = {pp87[99]};
    assign in4902_2 = {pp88[98]};
    Full_Adder FA_4902(s4902, c4902, in4902_1, in4902_2, pp86[100]);
    wire[0:0] s4903, in4903_1, in4903_2;
    wire c4903;
    assign in4903_1 = {pp90[96]};
    assign in4903_2 = {pp91[95]};
    Full_Adder FA_4903(s4903, c4903, in4903_1, in4903_2, pp89[97]);
    wire[0:0] s4904, in4904_1, in4904_2;
    wire c4904;
    assign in4904_1 = {pp93[93]};
    assign in4904_2 = {pp94[92]};
    Full_Adder FA_4904(s4904, c4904, in4904_1, in4904_2, pp92[94]);
    wire[0:0] s4905, in4905_1, in4905_2;
    wire c4905;
    assign in4905_1 = {pp61[126]};
    assign in4905_2 = {pp62[125]};
    Full_Adder FA_4905(s4905, c4905, in4905_1, in4905_2, pp60[127]);
    wire[0:0] s4906, in4906_1, in4906_2;
    wire c4906;
    assign in4906_1 = {pp64[123]};
    assign in4906_2 = {pp65[122]};
    Full_Adder FA_4906(s4906, c4906, in4906_1, in4906_2, pp63[124]);
    wire[0:0] s4907, in4907_1, in4907_2;
    wire c4907;
    assign in4907_1 = {pp67[120]};
    assign in4907_2 = {pp68[119]};
    Full_Adder FA_4907(s4907, c4907, in4907_1, in4907_2, pp66[121]);
    wire[0:0] s4908, in4908_1, in4908_2;
    wire c4908;
    assign in4908_1 = {pp70[117]};
    assign in4908_2 = {pp71[116]};
    Full_Adder FA_4908(s4908, c4908, in4908_1, in4908_2, pp69[118]);
    wire[0:0] s4909, in4909_1, in4909_2;
    wire c4909;
    assign in4909_1 = {pp73[114]};
    assign in4909_2 = {pp74[113]};
    Full_Adder FA_4909(s4909, c4909, in4909_1, in4909_2, pp72[115]);
    wire[0:0] s4910, in4910_1, in4910_2;
    wire c4910;
    assign in4910_1 = {pp76[111]};
    assign in4910_2 = {pp77[110]};
    Full_Adder FA_4910(s4910, c4910, in4910_1, in4910_2, pp75[112]);
    wire[0:0] s4911, in4911_1, in4911_2;
    wire c4911;
    assign in4911_1 = {pp79[108]};
    assign in4911_2 = {pp80[107]};
    Full_Adder FA_4911(s4911, c4911, in4911_1, in4911_2, pp78[109]);
    wire[0:0] s4912, in4912_1, in4912_2;
    wire c4912;
    assign in4912_1 = {pp82[105]};
    assign in4912_2 = {pp83[104]};
    Full_Adder FA_4912(s4912, c4912, in4912_1, in4912_2, pp81[106]);
    wire[0:0] s4913, in4913_1, in4913_2;
    wire c4913;
    assign in4913_1 = {pp85[102]};
    assign in4913_2 = {pp86[101]};
    Full_Adder FA_4913(s4913, c4913, in4913_1, in4913_2, pp84[103]);
    wire[0:0] s4914, in4914_1, in4914_2;
    wire c4914;
    assign in4914_1 = {pp88[99]};
    assign in4914_2 = {pp89[98]};
    Full_Adder FA_4914(s4914, c4914, in4914_1, in4914_2, pp87[100]);
    wire[0:0] s4915, in4915_1, in4915_2;
    wire c4915;
    assign in4915_1 = {pp91[96]};
    assign in4915_2 = {pp92[95]};
    Full_Adder FA_4915(s4915, c4915, in4915_1, in4915_2, pp90[97]);
    wire[0:0] s4916, in4916_1, in4916_2;
    wire c4916;
    assign in4916_1 = {pp62[126]};
    assign in4916_2 = {pp63[125]};
    Full_Adder FA_4916(s4916, c4916, in4916_1, in4916_2, pp61[127]);
    wire[0:0] s4917, in4917_1, in4917_2;
    wire c4917;
    assign in4917_1 = {pp65[123]};
    assign in4917_2 = {pp66[122]};
    Full_Adder FA_4917(s4917, c4917, in4917_1, in4917_2, pp64[124]);
    wire[0:0] s4918, in4918_1, in4918_2;
    wire c4918;
    assign in4918_1 = {pp68[120]};
    assign in4918_2 = {pp69[119]};
    Full_Adder FA_4918(s4918, c4918, in4918_1, in4918_2, pp67[121]);
    wire[0:0] s4919, in4919_1, in4919_2;
    wire c4919;
    assign in4919_1 = {pp71[117]};
    assign in4919_2 = {pp72[116]};
    Full_Adder FA_4919(s4919, c4919, in4919_1, in4919_2, pp70[118]);
    wire[0:0] s4920, in4920_1, in4920_2;
    wire c4920;
    assign in4920_1 = {pp74[114]};
    assign in4920_2 = {pp75[113]};
    Full_Adder FA_4920(s4920, c4920, in4920_1, in4920_2, pp73[115]);
    wire[0:0] s4921, in4921_1, in4921_2;
    wire c4921;
    assign in4921_1 = {pp77[111]};
    assign in4921_2 = {pp78[110]};
    Full_Adder FA_4921(s4921, c4921, in4921_1, in4921_2, pp76[112]);
    wire[0:0] s4922, in4922_1, in4922_2;
    wire c4922;
    assign in4922_1 = {pp80[108]};
    assign in4922_2 = {pp81[107]};
    Full_Adder FA_4922(s4922, c4922, in4922_1, in4922_2, pp79[109]);
    wire[0:0] s4923, in4923_1, in4923_2;
    wire c4923;
    assign in4923_1 = {pp83[105]};
    assign in4923_2 = {pp84[104]};
    Full_Adder FA_4923(s4923, c4923, in4923_1, in4923_2, pp82[106]);
    wire[0:0] s4924, in4924_1, in4924_2;
    wire c4924;
    assign in4924_1 = {pp86[102]};
    assign in4924_2 = {pp87[101]};
    Full_Adder FA_4924(s4924, c4924, in4924_1, in4924_2, pp85[103]);
    wire[0:0] s4925, in4925_1, in4925_2;
    wire c4925;
    assign in4925_1 = {pp89[99]};
    assign in4925_2 = {pp90[98]};
    Full_Adder FA_4925(s4925, c4925, in4925_1, in4925_2, pp88[100]);
    wire[0:0] s4926, in4926_1, in4926_2;
    wire c4926;
    assign in4926_1 = {pp63[126]};
    assign in4926_2 = {pp64[125]};
    Full_Adder FA_4926(s4926, c4926, in4926_1, in4926_2, pp62[127]);
    wire[0:0] s4927, in4927_1, in4927_2;
    wire c4927;
    assign in4927_1 = {pp66[123]};
    assign in4927_2 = {pp67[122]};
    Full_Adder FA_4927(s4927, c4927, in4927_1, in4927_2, pp65[124]);
    wire[0:0] s4928, in4928_1, in4928_2;
    wire c4928;
    assign in4928_1 = {pp69[120]};
    assign in4928_2 = {pp70[119]};
    Full_Adder FA_4928(s4928, c4928, in4928_1, in4928_2, pp68[121]);
    wire[0:0] s4929, in4929_1, in4929_2;
    wire c4929;
    assign in4929_1 = {pp72[117]};
    assign in4929_2 = {pp73[116]};
    Full_Adder FA_4929(s4929, c4929, in4929_1, in4929_2, pp71[118]);
    wire[0:0] s4930, in4930_1, in4930_2;
    wire c4930;
    assign in4930_1 = {pp75[114]};
    assign in4930_2 = {pp76[113]};
    Full_Adder FA_4930(s4930, c4930, in4930_1, in4930_2, pp74[115]);
    wire[0:0] s4931, in4931_1, in4931_2;
    wire c4931;
    assign in4931_1 = {pp78[111]};
    assign in4931_2 = {pp79[110]};
    Full_Adder FA_4931(s4931, c4931, in4931_1, in4931_2, pp77[112]);
    wire[0:0] s4932, in4932_1, in4932_2;
    wire c4932;
    assign in4932_1 = {pp81[108]};
    assign in4932_2 = {pp82[107]};
    Full_Adder FA_4932(s4932, c4932, in4932_1, in4932_2, pp80[109]);
    wire[0:0] s4933, in4933_1, in4933_2;
    wire c4933;
    assign in4933_1 = {pp84[105]};
    assign in4933_2 = {pp85[104]};
    Full_Adder FA_4933(s4933, c4933, in4933_1, in4933_2, pp83[106]);
    wire[0:0] s4934, in4934_1, in4934_2;
    wire c4934;
    assign in4934_1 = {pp87[102]};
    assign in4934_2 = {pp88[101]};
    Full_Adder FA_4934(s4934, c4934, in4934_1, in4934_2, pp86[103]);
    wire[0:0] s4935, in4935_1, in4935_2;
    wire c4935;
    assign in4935_1 = {pp64[126]};
    assign in4935_2 = {pp65[125]};
    Full_Adder FA_4935(s4935, c4935, in4935_1, in4935_2, pp63[127]);
    wire[0:0] s4936, in4936_1, in4936_2;
    wire c4936;
    assign in4936_1 = {pp67[123]};
    assign in4936_2 = {pp68[122]};
    Full_Adder FA_4936(s4936, c4936, in4936_1, in4936_2, pp66[124]);
    wire[0:0] s4937, in4937_1, in4937_2;
    wire c4937;
    assign in4937_1 = {pp70[120]};
    assign in4937_2 = {pp71[119]};
    Full_Adder FA_4937(s4937, c4937, in4937_1, in4937_2, pp69[121]);
    wire[0:0] s4938, in4938_1, in4938_2;
    wire c4938;
    assign in4938_1 = {pp73[117]};
    assign in4938_2 = {pp74[116]};
    Full_Adder FA_4938(s4938, c4938, in4938_1, in4938_2, pp72[118]);
    wire[0:0] s4939, in4939_1, in4939_2;
    wire c4939;
    assign in4939_1 = {pp76[114]};
    assign in4939_2 = {pp77[113]};
    Full_Adder FA_4939(s4939, c4939, in4939_1, in4939_2, pp75[115]);
    wire[0:0] s4940, in4940_1, in4940_2;
    wire c4940;
    assign in4940_1 = {pp79[111]};
    assign in4940_2 = {pp80[110]};
    Full_Adder FA_4940(s4940, c4940, in4940_1, in4940_2, pp78[112]);
    wire[0:0] s4941, in4941_1, in4941_2;
    wire c4941;
    assign in4941_1 = {pp82[108]};
    assign in4941_2 = {pp83[107]};
    Full_Adder FA_4941(s4941, c4941, in4941_1, in4941_2, pp81[109]);
    wire[0:0] s4942, in4942_1, in4942_2;
    wire c4942;
    assign in4942_1 = {pp85[105]};
    assign in4942_2 = {pp86[104]};
    Full_Adder FA_4942(s4942, c4942, in4942_1, in4942_2, pp84[106]);
    wire[0:0] s4943, in4943_1, in4943_2;
    wire c4943;
    assign in4943_1 = {pp65[126]};
    assign in4943_2 = {pp66[125]};
    Full_Adder FA_4943(s4943, c4943, in4943_1, in4943_2, pp64[127]);
    wire[0:0] s4944, in4944_1, in4944_2;
    wire c4944;
    assign in4944_1 = {pp68[123]};
    assign in4944_2 = {pp69[122]};
    Full_Adder FA_4944(s4944, c4944, in4944_1, in4944_2, pp67[124]);
    wire[0:0] s4945, in4945_1, in4945_2;
    wire c4945;
    assign in4945_1 = {pp71[120]};
    assign in4945_2 = {pp72[119]};
    Full_Adder FA_4945(s4945, c4945, in4945_1, in4945_2, pp70[121]);
    wire[0:0] s4946, in4946_1, in4946_2;
    wire c4946;
    assign in4946_1 = {pp74[117]};
    assign in4946_2 = {pp75[116]};
    Full_Adder FA_4946(s4946, c4946, in4946_1, in4946_2, pp73[118]);
    wire[0:0] s4947, in4947_1, in4947_2;
    wire c4947;
    assign in4947_1 = {pp77[114]};
    assign in4947_2 = {pp78[113]};
    Full_Adder FA_4947(s4947, c4947, in4947_1, in4947_2, pp76[115]);
    wire[0:0] s4948, in4948_1, in4948_2;
    wire c4948;
    assign in4948_1 = {pp80[111]};
    assign in4948_2 = {pp81[110]};
    Full_Adder FA_4948(s4948, c4948, in4948_1, in4948_2, pp79[112]);
    wire[0:0] s4949, in4949_1, in4949_2;
    wire c4949;
    assign in4949_1 = {pp83[108]};
    assign in4949_2 = {pp84[107]};
    Full_Adder FA_4949(s4949, c4949, in4949_1, in4949_2, pp82[109]);
    wire[0:0] s4950, in4950_1, in4950_2;
    wire c4950;
    assign in4950_1 = {pp66[126]};
    assign in4950_2 = {pp67[125]};
    Full_Adder FA_4950(s4950, c4950, in4950_1, in4950_2, pp65[127]);
    wire[0:0] s4951, in4951_1, in4951_2;
    wire c4951;
    assign in4951_1 = {pp69[123]};
    assign in4951_2 = {pp70[122]};
    Full_Adder FA_4951(s4951, c4951, in4951_1, in4951_2, pp68[124]);
    wire[0:0] s4952, in4952_1, in4952_2;
    wire c4952;
    assign in4952_1 = {pp72[120]};
    assign in4952_2 = {pp73[119]};
    Full_Adder FA_4952(s4952, c4952, in4952_1, in4952_2, pp71[121]);
    wire[0:0] s4953, in4953_1, in4953_2;
    wire c4953;
    assign in4953_1 = {pp75[117]};
    assign in4953_2 = {pp76[116]};
    Full_Adder FA_4953(s4953, c4953, in4953_1, in4953_2, pp74[118]);
    wire[0:0] s4954, in4954_1, in4954_2;
    wire c4954;
    assign in4954_1 = {pp78[114]};
    assign in4954_2 = {pp79[113]};
    Full_Adder FA_4954(s4954, c4954, in4954_1, in4954_2, pp77[115]);
    wire[0:0] s4955, in4955_1, in4955_2;
    wire c4955;
    assign in4955_1 = {pp81[111]};
    assign in4955_2 = {pp82[110]};
    Full_Adder FA_4955(s4955, c4955, in4955_1, in4955_2, pp80[112]);
    wire[0:0] s4956, in4956_1, in4956_2;
    wire c4956;
    assign in4956_1 = {pp67[126]};
    assign in4956_2 = {pp68[125]};
    Full_Adder FA_4956(s4956, c4956, in4956_1, in4956_2, pp66[127]);
    wire[0:0] s4957, in4957_1, in4957_2;
    wire c4957;
    assign in4957_1 = {pp70[123]};
    assign in4957_2 = {pp71[122]};
    Full_Adder FA_4957(s4957, c4957, in4957_1, in4957_2, pp69[124]);
    wire[0:0] s4958, in4958_1, in4958_2;
    wire c4958;
    assign in4958_1 = {pp73[120]};
    assign in4958_2 = {pp74[119]};
    Full_Adder FA_4958(s4958, c4958, in4958_1, in4958_2, pp72[121]);
    wire[0:0] s4959, in4959_1, in4959_2;
    wire c4959;
    assign in4959_1 = {pp76[117]};
    assign in4959_2 = {pp77[116]};
    Full_Adder FA_4959(s4959, c4959, in4959_1, in4959_2, pp75[118]);
    wire[0:0] s4960, in4960_1, in4960_2;
    wire c4960;
    assign in4960_1 = {pp79[114]};
    assign in4960_2 = {pp80[113]};
    Full_Adder FA_4960(s4960, c4960, in4960_1, in4960_2, pp78[115]);
    wire[0:0] s4961, in4961_1, in4961_2;
    wire c4961;
    assign in4961_1 = {pp68[126]};
    assign in4961_2 = {pp69[125]};
    Full_Adder FA_4961(s4961, c4961, in4961_1, in4961_2, pp67[127]);
    wire[0:0] s4962, in4962_1, in4962_2;
    wire c4962;
    assign in4962_1 = {pp71[123]};
    assign in4962_2 = {pp72[122]};
    Full_Adder FA_4962(s4962, c4962, in4962_1, in4962_2, pp70[124]);
    wire[0:0] s4963, in4963_1, in4963_2;
    wire c4963;
    assign in4963_1 = {pp74[120]};
    assign in4963_2 = {pp75[119]};
    Full_Adder FA_4963(s4963, c4963, in4963_1, in4963_2, pp73[121]);
    wire[0:0] s4964, in4964_1, in4964_2;
    wire c4964;
    assign in4964_1 = {pp77[117]};
    assign in4964_2 = {pp78[116]};
    Full_Adder FA_4964(s4964, c4964, in4964_1, in4964_2, pp76[118]);
    wire[0:0] s4965, in4965_1, in4965_2;
    wire c4965;
    assign in4965_1 = {pp69[126]};
    assign in4965_2 = {pp70[125]};
    Full_Adder FA_4965(s4965, c4965, in4965_1, in4965_2, pp68[127]);
    wire[0:0] s4966, in4966_1, in4966_2;
    wire c4966;
    assign in4966_1 = {pp72[123]};
    assign in4966_2 = {pp73[122]};
    Full_Adder FA_4966(s4966, c4966, in4966_1, in4966_2, pp71[124]);
    wire[0:0] s4967, in4967_1, in4967_2;
    wire c4967;
    assign in4967_1 = {pp75[120]};
    assign in4967_2 = {pp76[119]};
    Full_Adder FA_4967(s4967, c4967, in4967_1, in4967_2, pp74[121]);
    wire[0:0] s4968, in4968_1, in4968_2;
    wire c4968;
    assign in4968_1 = {pp70[126]};
    assign in4968_2 = {pp71[125]};
    Full_Adder FA_4968(s4968, c4968, in4968_1, in4968_2, pp69[127]);
    wire[0:0] s4969, in4969_1, in4969_2;
    wire c4969;
    assign in4969_1 = {pp73[123]};
    assign in4969_2 = {pp74[122]};
    Full_Adder FA_4969(s4969, c4969, in4969_1, in4969_2, pp72[124]);
    wire[0:0] s4970, in4970_1, in4970_2;
    wire c4970;
    assign in4970_1 = {pp71[126]};
    assign in4970_2 = {pp72[125]};
    Full_Adder FA_4970(s4970, c4970, in4970_1, in4970_2, pp70[127]);

    /*Stage 3*/
    wire[0:0] s4971, in4971_1, in4971_2;
    wire c4971;
    assign in4971_1 = {pp0[39]};
    assign in4971_2 = {pp1[38]};
    Half_Adder HA_4971(s4971, c4971, in4971_1, in4971_2);
    wire[0:0] s4972, in4972_1, in4972_2;
    wire c4972;
    assign in4972_1 = {pp1[39]};
    assign in4972_2 = {pp2[38]};
    Full_Adder FA_4972(s4972, c4972, in4972_1, in4972_2, pp0[40]);
    wire[0:0] s4973, in4973_1, in4973_2;
    wire c4973;
    assign in4973_1 = {pp3[37]};
    assign in4973_2 = {pp4[36]};
    Half_Adder HA_4973(s4973, c4973, in4973_1, in4973_2);
    wire[0:0] s4974, in4974_1, in4974_2;
    wire c4974;
    assign in4974_1 = {pp1[40]};
    assign in4974_2 = {pp2[39]};
    Full_Adder FA_4974(s4974, c4974, in4974_1, in4974_2, pp0[41]);
    wire[0:0] s4975, in4975_1, in4975_2;
    wire c4975;
    assign in4975_1 = {pp4[37]};
    assign in4975_2 = {pp5[36]};
    Full_Adder FA_4975(s4975, c4975, in4975_1, in4975_2, pp3[38]);
    wire[0:0] s4976, in4976_1, in4976_2;
    wire c4976;
    assign in4976_1 = {pp6[35]};
    assign in4976_2 = {pp7[34]};
    Half_Adder HA_4976(s4976, c4976, in4976_1, in4976_2);
    wire[0:0] s4977, in4977_1, in4977_2;
    wire c4977;
    assign in4977_1 = {pp1[41]};
    assign in4977_2 = {pp2[40]};
    Full_Adder FA_4977(s4977, c4977, in4977_1, in4977_2, pp0[42]);
    wire[0:0] s4978, in4978_1, in4978_2;
    wire c4978;
    assign in4978_1 = {pp4[38]};
    assign in4978_2 = {pp5[37]};
    Full_Adder FA_4978(s4978, c4978, in4978_1, in4978_2, pp3[39]);
    wire[0:0] s4979, in4979_1, in4979_2;
    wire c4979;
    assign in4979_1 = {pp7[35]};
    assign in4979_2 = {pp8[34]};
    Full_Adder FA_4979(s4979, c4979, in4979_1, in4979_2, pp6[36]);
    wire[0:0] s4980, in4980_1, in4980_2;
    wire c4980;
    assign in4980_1 = {pp9[33]};
    assign in4980_2 = {pp10[32]};
    Half_Adder HA_4980(s4980, c4980, in4980_1, in4980_2);
    wire[0:0] s4981, in4981_1, in4981_2;
    wire c4981;
    assign in4981_1 = {pp1[42]};
    assign in4981_2 = {pp2[41]};
    Full_Adder FA_4981(s4981, c4981, in4981_1, in4981_2, pp0[43]);
    wire[0:0] s4982, in4982_1, in4982_2;
    wire c4982;
    assign in4982_1 = {pp4[39]};
    assign in4982_2 = {pp5[38]};
    Full_Adder FA_4982(s4982, c4982, in4982_1, in4982_2, pp3[40]);
    wire[0:0] s4983, in4983_1, in4983_2;
    wire c4983;
    assign in4983_1 = {pp7[36]};
    assign in4983_2 = {pp8[35]};
    Full_Adder FA_4983(s4983, c4983, in4983_1, in4983_2, pp6[37]);
    wire[0:0] s4984, in4984_1, in4984_2;
    wire c4984;
    assign in4984_1 = {pp10[33]};
    assign in4984_2 = {pp11[32]};
    Full_Adder FA_4984(s4984, c4984, in4984_1, in4984_2, pp9[34]);
    wire[0:0] s4985, in4985_1, in4985_2;
    wire c4985;
    assign in4985_1 = {pp12[31]};
    assign in4985_2 = {pp13[30]};
    Half_Adder HA_4985(s4985, c4985, in4985_1, in4985_2);
    wire[0:0] s4986, in4986_1, in4986_2;
    wire c4986;
    assign in4986_1 = {pp1[43]};
    assign in4986_2 = {pp2[42]};
    Full_Adder FA_4986(s4986, c4986, in4986_1, in4986_2, pp0[44]);
    wire[0:0] s4987, in4987_1, in4987_2;
    wire c4987;
    assign in4987_1 = {pp4[40]};
    assign in4987_2 = {pp5[39]};
    Full_Adder FA_4987(s4987, c4987, in4987_1, in4987_2, pp3[41]);
    wire[0:0] s4988, in4988_1, in4988_2;
    wire c4988;
    assign in4988_1 = {pp7[37]};
    assign in4988_2 = {pp8[36]};
    Full_Adder FA_4988(s4988, c4988, in4988_1, in4988_2, pp6[38]);
    wire[0:0] s4989, in4989_1, in4989_2;
    wire c4989;
    assign in4989_1 = {pp10[34]};
    assign in4989_2 = {pp11[33]};
    Full_Adder FA_4989(s4989, c4989, in4989_1, in4989_2, pp9[35]);
    wire[0:0] s4990, in4990_1, in4990_2;
    wire c4990;
    assign in4990_1 = {pp13[31]};
    assign in4990_2 = {pp14[30]};
    Full_Adder FA_4990(s4990, c4990, in4990_1, in4990_2, pp12[32]);
    wire[0:0] s4991, in4991_1, in4991_2;
    wire c4991;
    assign in4991_1 = {pp15[29]};
    assign in4991_2 = {pp16[28]};
    Half_Adder HA_4991(s4991, c4991, in4991_1, in4991_2);
    wire[0:0] s4992, in4992_1, in4992_2;
    wire c4992;
    assign in4992_1 = {pp1[44]};
    assign in4992_2 = {pp2[43]};
    Full_Adder FA_4992(s4992, c4992, in4992_1, in4992_2, pp0[45]);
    wire[0:0] s4993, in4993_1, in4993_2;
    wire c4993;
    assign in4993_1 = {pp4[41]};
    assign in4993_2 = {pp5[40]};
    Full_Adder FA_4993(s4993, c4993, in4993_1, in4993_2, pp3[42]);
    wire[0:0] s4994, in4994_1, in4994_2;
    wire c4994;
    assign in4994_1 = {pp7[38]};
    assign in4994_2 = {pp8[37]};
    Full_Adder FA_4994(s4994, c4994, in4994_1, in4994_2, pp6[39]);
    wire[0:0] s4995, in4995_1, in4995_2;
    wire c4995;
    assign in4995_1 = {pp10[35]};
    assign in4995_2 = {pp11[34]};
    Full_Adder FA_4995(s4995, c4995, in4995_1, in4995_2, pp9[36]);
    wire[0:0] s4996, in4996_1, in4996_2;
    wire c4996;
    assign in4996_1 = {pp13[32]};
    assign in4996_2 = {pp14[31]};
    Full_Adder FA_4996(s4996, c4996, in4996_1, in4996_2, pp12[33]);
    wire[0:0] s4997, in4997_1, in4997_2;
    wire c4997;
    assign in4997_1 = {pp16[29]};
    assign in4997_2 = {pp17[28]};
    Full_Adder FA_4997(s4997, c4997, in4997_1, in4997_2, pp15[30]);
    wire[0:0] s4998, in4998_1, in4998_2;
    wire c4998;
    assign in4998_1 = {pp18[27]};
    assign in4998_2 = {pp19[26]};
    Half_Adder HA_4998(s4998, c4998, in4998_1, in4998_2);
    wire[0:0] s4999, in4999_1, in4999_2;
    wire c4999;
    assign in4999_1 = {pp1[45]};
    assign in4999_2 = {pp2[44]};
    Full_Adder FA_4999(s4999, c4999, in4999_1, in4999_2, pp0[46]);
    wire[0:0] s5000, in5000_1, in5000_2;
    wire c5000;
    assign in5000_1 = {pp4[42]};
    assign in5000_2 = {pp5[41]};
    Full_Adder FA_5000(s5000, c5000, in5000_1, in5000_2, pp3[43]);
    wire[0:0] s5001, in5001_1, in5001_2;
    wire c5001;
    assign in5001_1 = {pp7[39]};
    assign in5001_2 = {pp8[38]};
    Full_Adder FA_5001(s5001, c5001, in5001_1, in5001_2, pp6[40]);
    wire[0:0] s5002, in5002_1, in5002_2;
    wire c5002;
    assign in5002_1 = {pp10[36]};
    assign in5002_2 = {pp11[35]};
    Full_Adder FA_5002(s5002, c5002, in5002_1, in5002_2, pp9[37]);
    wire[0:0] s5003, in5003_1, in5003_2;
    wire c5003;
    assign in5003_1 = {pp13[33]};
    assign in5003_2 = {pp14[32]};
    Full_Adder FA_5003(s5003, c5003, in5003_1, in5003_2, pp12[34]);
    wire[0:0] s5004, in5004_1, in5004_2;
    wire c5004;
    assign in5004_1 = {pp16[30]};
    assign in5004_2 = {pp17[29]};
    Full_Adder FA_5004(s5004, c5004, in5004_1, in5004_2, pp15[31]);
    wire[0:0] s5005, in5005_1, in5005_2;
    wire c5005;
    assign in5005_1 = {pp19[27]};
    assign in5005_2 = {pp20[26]};
    Full_Adder FA_5005(s5005, c5005, in5005_1, in5005_2, pp18[28]);
    wire[0:0] s5006, in5006_1, in5006_2;
    wire c5006;
    assign in5006_1 = {pp21[25]};
    assign in5006_2 = {pp22[24]};
    Half_Adder HA_5006(s5006, c5006, in5006_1, in5006_2);
    wire[0:0] s5007, in5007_1, in5007_2;
    wire c5007;
    assign in5007_1 = {pp1[46]};
    assign in5007_2 = {pp2[45]};
    Full_Adder FA_5007(s5007, c5007, in5007_1, in5007_2, pp0[47]);
    wire[0:0] s5008, in5008_1, in5008_2;
    wire c5008;
    assign in5008_1 = {pp4[43]};
    assign in5008_2 = {pp5[42]};
    Full_Adder FA_5008(s5008, c5008, in5008_1, in5008_2, pp3[44]);
    wire[0:0] s5009, in5009_1, in5009_2;
    wire c5009;
    assign in5009_1 = {pp7[40]};
    assign in5009_2 = {pp8[39]};
    Full_Adder FA_5009(s5009, c5009, in5009_1, in5009_2, pp6[41]);
    wire[0:0] s5010, in5010_1, in5010_2;
    wire c5010;
    assign in5010_1 = {pp10[37]};
    assign in5010_2 = {pp11[36]};
    Full_Adder FA_5010(s5010, c5010, in5010_1, in5010_2, pp9[38]);
    wire[0:0] s5011, in5011_1, in5011_2;
    wire c5011;
    assign in5011_1 = {pp13[34]};
    assign in5011_2 = {pp14[33]};
    Full_Adder FA_5011(s5011, c5011, in5011_1, in5011_2, pp12[35]);
    wire[0:0] s5012, in5012_1, in5012_2;
    wire c5012;
    assign in5012_1 = {pp16[31]};
    assign in5012_2 = {pp17[30]};
    Full_Adder FA_5012(s5012, c5012, in5012_1, in5012_2, pp15[32]);
    wire[0:0] s5013, in5013_1, in5013_2;
    wire c5013;
    assign in5013_1 = {pp19[28]};
    assign in5013_2 = {pp20[27]};
    Full_Adder FA_5013(s5013, c5013, in5013_1, in5013_2, pp18[29]);
    wire[0:0] s5014, in5014_1, in5014_2;
    wire c5014;
    assign in5014_1 = {pp22[25]};
    assign in5014_2 = {pp23[24]};
    Full_Adder FA_5014(s5014, c5014, in5014_1, in5014_2, pp21[26]);
    wire[0:0] s5015, in5015_1, in5015_2;
    wire c5015;
    assign in5015_1 = {pp24[23]};
    assign in5015_2 = {pp25[22]};
    Half_Adder HA_5015(s5015, c5015, in5015_1, in5015_2);
    wire[0:0] s5016, in5016_1, in5016_2;
    wire c5016;
    assign in5016_1 = {pp1[47]};
    assign in5016_2 = {pp2[46]};
    Full_Adder FA_5016(s5016, c5016, in5016_1, in5016_2, pp0[48]);
    wire[0:0] s5017, in5017_1, in5017_2;
    wire c5017;
    assign in5017_1 = {pp4[44]};
    assign in5017_2 = {pp5[43]};
    Full_Adder FA_5017(s5017, c5017, in5017_1, in5017_2, pp3[45]);
    wire[0:0] s5018, in5018_1, in5018_2;
    wire c5018;
    assign in5018_1 = {pp7[41]};
    assign in5018_2 = {pp8[40]};
    Full_Adder FA_5018(s5018, c5018, in5018_1, in5018_2, pp6[42]);
    wire[0:0] s5019, in5019_1, in5019_2;
    wire c5019;
    assign in5019_1 = {pp10[38]};
    assign in5019_2 = {pp11[37]};
    Full_Adder FA_5019(s5019, c5019, in5019_1, in5019_2, pp9[39]);
    wire[0:0] s5020, in5020_1, in5020_2;
    wire c5020;
    assign in5020_1 = {pp13[35]};
    assign in5020_2 = {pp14[34]};
    Full_Adder FA_5020(s5020, c5020, in5020_1, in5020_2, pp12[36]);
    wire[0:0] s5021, in5021_1, in5021_2;
    wire c5021;
    assign in5021_1 = {pp16[32]};
    assign in5021_2 = {pp17[31]};
    Full_Adder FA_5021(s5021, c5021, in5021_1, in5021_2, pp15[33]);
    wire[0:0] s5022, in5022_1, in5022_2;
    wire c5022;
    assign in5022_1 = {pp19[29]};
    assign in5022_2 = {pp20[28]};
    Full_Adder FA_5022(s5022, c5022, in5022_1, in5022_2, pp18[30]);
    wire[0:0] s5023, in5023_1, in5023_2;
    wire c5023;
    assign in5023_1 = {pp22[26]};
    assign in5023_2 = {pp23[25]};
    Full_Adder FA_5023(s5023, c5023, in5023_1, in5023_2, pp21[27]);
    wire[0:0] s5024, in5024_1, in5024_2;
    wire c5024;
    assign in5024_1 = {pp25[23]};
    assign in5024_2 = {pp26[22]};
    Full_Adder FA_5024(s5024, c5024, in5024_1, in5024_2, pp24[24]);
    wire[0:0] s5025, in5025_1, in5025_2;
    wire c5025;
    assign in5025_1 = {pp27[21]};
    assign in5025_2 = {pp28[20]};
    Half_Adder HA_5025(s5025, c5025, in5025_1, in5025_2);
    wire[0:0] s5026, in5026_1, in5026_2;
    wire c5026;
    assign in5026_1 = {pp1[48]};
    assign in5026_2 = {pp2[47]};
    Full_Adder FA_5026(s5026, c5026, in5026_1, in5026_2, pp0[49]);
    wire[0:0] s5027, in5027_1, in5027_2;
    wire c5027;
    assign in5027_1 = {pp4[45]};
    assign in5027_2 = {pp5[44]};
    Full_Adder FA_5027(s5027, c5027, in5027_1, in5027_2, pp3[46]);
    wire[0:0] s5028, in5028_1, in5028_2;
    wire c5028;
    assign in5028_1 = {pp7[42]};
    assign in5028_2 = {pp8[41]};
    Full_Adder FA_5028(s5028, c5028, in5028_1, in5028_2, pp6[43]);
    wire[0:0] s5029, in5029_1, in5029_2;
    wire c5029;
    assign in5029_1 = {pp10[39]};
    assign in5029_2 = {pp11[38]};
    Full_Adder FA_5029(s5029, c5029, in5029_1, in5029_2, pp9[40]);
    wire[0:0] s5030, in5030_1, in5030_2;
    wire c5030;
    assign in5030_1 = {pp13[36]};
    assign in5030_2 = {pp14[35]};
    Full_Adder FA_5030(s5030, c5030, in5030_1, in5030_2, pp12[37]);
    wire[0:0] s5031, in5031_1, in5031_2;
    wire c5031;
    assign in5031_1 = {pp16[33]};
    assign in5031_2 = {pp17[32]};
    Full_Adder FA_5031(s5031, c5031, in5031_1, in5031_2, pp15[34]);
    wire[0:0] s5032, in5032_1, in5032_2;
    wire c5032;
    assign in5032_1 = {pp19[30]};
    assign in5032_2 = {pp20[29]};
    Full_Adder FA_5032(s5032, c5032, in5032_1, in5032_2, pp18[31]);
    wire[0:0] s5033, in5033_1, in5033_2;
    wire c5033;
    assign in5033_1 = {pp22[27]};
    assign in5033_2 = {pp23[26]};
    Full_Adder FA_5033(s5033, c5033, in5033_1, in5033_2, pp21[28]);
    wire[0:0] s5034, in5034_1, in5034_2;
    wire c5034;
    assign in5034_1 = {pp25[24]};
    assign in5034_2 = {pp26[23]};
    Full_Adder FA_5034(s5034, c5034, in5034_1, in5034_2, pp24[25]);
    wire[0:0] s5035, in5035_1, in5035_2;
    wire c5035;
    assign in5035_1 = {pp28[21]};
    assign in5035_2 = {pp29[20]};
    Full_Adder FA_5035(s5035, c5035, in5035_1, in5035_2, pp27[22]);
    wire[0:0] s5036, in5036_1, in5036_2;
    wire c5036;
    assign in5036_1 = {pp30[19]};
    assign in5036_2 = {pp31[18]};
    Half_Adder HA_5036(s5036, c5036, in5036_1, in5036_2);
    wire[0:0] s5037, in5037_1, in5037_2;
    wire c5037;
    assign in5037_1 = {pp1[49]};
    assign in5037_2 = {pp2[48]};
    Full_Adder FA_5037(s5037, c5037, in5037_1, in5037_2, pp0[50]);
    wire[0:0] s5038, in5038_1, in5038_2;
    wire c5038;
    assign in5038_1 = {pp4[46]};
    assign in5038_2 = {pp5[45]};
    Full_Adder FA_5038(s5038, c5038, in5038_1, in5038_2, pp3[47]);
    wire[0:0] s5039, in5039_1, in5039_2;
    wire c5039;
    assign in5039_1 = {pp7[43]};
    assign in5039_2 = {pp8[42]};
    Full_Adder FA_5039(s5039, c5039, in5039_1, in5039_2, pp6[44]);
    wire[0:0] s5040, in5040_1, in5040_2;
    wire c5040;
    assign in5040_1 = {pp10[40]};
    assign in5040_2 = {pp11[39]};
    Full_Adder FA_5040(s5040, c5040, in5040_1, in5040_2, pp9[41]);
    wire[0:0] s5041, in5041_1, in5041_2;
    wire c5041;
    assign in5041_1 = {pp13[37]};
    assign in5041_2 = {pp14[36]};
    Full_Adder FA_5041(s5041, c5041, in5041_1, in5041_2, pp12[38]);
    wire[0:0] s5042, in5042_1, in5042_2;
    wire c5042;
    assign in5042_1 = {pp16[34]};
    assign in5042_2 = {pp17[33]};
    Full_Adder FA_5042(s5042, c5042, in5042_1, in5042_2, pp15[35]);
    wire[0:0] s5043, in5043_1, in5043_2;
    wire c5043;
    assign in5043_1 = {pp19[31]};
    assign in5043_2 = {pp20[30]};
    Full_Adder FA_5043(s5043, c5043, in5043_1, in5043_2, pp18[32]);
    wire[0:0] s5044, in5044_1, in5044_2;
    wire c5044;
    assign in5044_1 = {pp22[28]};
    assign in5044_2 = {pp23[27]};
    Full_Adder FA_5044(s5044, c5044, in5044_1, in5044_2, pp21[29]);
    wire[0:0] s5045, in5045_1, in5045_2;
    wire c5045;
    assign in5045_1 = {pp25[25]};
    assign in5045_2 = {pp26[24]};
    Full_Adder FA_5045(s5045, c5045, in5045_1, in5045_2, pp24[26]);
    wire[0:0] s5046, in5046_1, in5046_2;
    wire c5046;
    assign in5046_1 = {pp28[22]};
    assign in5046_2 = {pp29[21]};
    Full_Adder FA_5046(s5046, c5046, in5046_1, in5046_2, pp27[23]);
    wire[0:0] s5047, in5047_1, in5047_2;
    wire c5047;
    assign in5047_1 = {pp31[19]};
    assign in5047_2 = {pp32[18]};
    Full_Adder FA_5047(s5047, c5047, in5047_1, in5047_2, pp30[20]);
    wire[0:0] s5048, in5048_1, in5048_2;
    wire c5048;
    assign in5048_1 = {pp33[17]};
    assign in5048_2 = {pp34[16]};
    Half_Adder HA_5048(s5048, c5048, in5048_1, in5048_2);
    wire[0:0] s5049, in5049_1, in5049_2;
    wire c5049;
    assign in5049_1 = {pp1[50]};
    assign in5049_2 = {pp2[49]};
    Full_Adder FA_5049(s5049, c5049, in5049_1, in5049_2, pp0[51]);
    wire[0:0] s5050, in5050_1, in5050_2;
    wire c5050;
    assign in5050_1 = {pp4[47]};
    assign in5050_2 = {pp5[46]};
    Full_Adder FA_5050(s5050, c5050, in5050_1, in5050_2, pp3[48]);
    wire[0:0] s5051, in5051_1, in5051_2;
    wire c5051;
    assign in5051_1 = {pp7[44]};
    assign in5051_2 = {pp8[43]};
    Full_Adder FA_5051(s5051, c5051, in5051_1, in5051_2, pp6[45]);
    wire[0:0] s5052, in5052_1, in5052_2;
    wire c5052;
    assign in5052_1 = {pp10[41]};
    assign in5052_2 = {pp11[40]};
    Full_Adder FA_5052(s5052, c5052, in5052_1, in5052_2, pp9[42]);
    wire[0:0] s5053, in5053_1, in5053_2;
    wire c5053;
    assign in5053_1 = {pp13[38]};
    assign in5053_2 = {pp14[37]};
    Full_Adder FA_5053(s5053, c5053, in5053_1, in5053_2, pp12[39]);
    wire[0:0] s5054, in5054_1, in5054_2;
    wire c5054;
    assign in5054_1 = {pp16[35]};
    assign in5054_2 = {pp17[34]};
    Full_Adder FA_5054(s5054, c5054, in5054_1, in5054_2, pp15[36]);
    wire[0:0] s5055, in5055_1, in5055_2;
    wire c5055;
    assign in5055_1 = {pp19[32]};
    assign in5055_2 = {pp20[31]};
    Full_Adder FA_5055(s5055, c5055, in5055_1, in5055_2, pp18[33]);
    wire[0:0] s5056, in5056_1, in5056_2;
    wire c5056;
    assign in5056_1 = {pp22[29]};
    assign in5056_2 = {pp23[28]};
    Full_Adder FA_5056(s5056, c5056, in5056_1, in5056_2, pp21[30]);
    wire[0:0] s5057, in5057_1, in5057_2;
    wire c5057;
    assign in5057_1 = {pp25[26]};
    assign in5057_2 = {pp26[25]};
    Full_Adder FA_5057(s5057, c5057, in5057_1, in5057_2, pp24[27]);
    wire[0:0] s5058, in5058_1, in5058_2;
    wire c5058;
    assign in5058_1 = {pp28[23]};
    assign in5058_2 = {pp29[22]};
    Full_Adder FA_5058(s5058, c5058, in5058_1, in5058_2, pp27[24]);
    wire[0:0] s5059, in5059_1, in5059_2;
    wire c5059;
    assign in5059_1 = {pp31[20]};
    assign in5059_2 = {pp32[19]};
    Full_Adder FA_5059(s5059, c5059, in5059_1, in5059_2, pp30[21]);
    wire[0:0] s5060, in5060_1, in5060_2;
    wire c5060;
    assign in5060_1 = {pp34[17]};
    assign in5060_2 = {pp35[16]};
    Full_Adder FA_5060(s5060, c5060, in5060_1, in5060_2, pp33[18]);
    wire[0:0] s5061, in5061_1, in5061_2;
    wire c5061;
    assign in5061_1 = {pp36[15]};
    assign in5061_2 = {pp37[14]};
    Half_Adder HA_5061(s5061, c5061, in5061_1, in5061_2);
    wire[0:0] s5062, in5062_1, in5062_2;
    wire c5062;
    assign in5062_1 = {pp1[51]};
    assign in5062_2 = {pp2[50]};
    Full_Adder FA_5062(s5062, c5062, in5062_1, in5062_2, pp0[52]);
    wire[0:0] s5063, in5063_1, in5063_2;
    wire c5063;
    assign in5063_1 = {pp4[48]};
    assign in5063_2 = {pp5[47]};
    Full_Adder FA_5063(s5063, c5063, in5063_1, in5063_2, pp3[49]);
    wire[0:0] s5064, in5064_1, in5064_2;
    wire c5064;
    assign in5064_1 = {pp7[45]};
    assign in5064_2 = {pp8[44]};
    Full_Adder FA_5064(s5064, c5064, in5064_1, in5064_2, pp6[46]);
    wire[0:0] s5065, in5065_1, in5065_2;
    wire c5065;
    assign in5065_1 = {pp10[42]};
    assign in5065_2 = {pp11[41]};
    Full_Adder FA_5065(s5065, c5065, in5065_1, in5065_2, pp9[43]);
    wire[0:0] s5066, in5066_1, in5066_2;
    wire c5066;
    assign in5066_1 = {pp13[39]};
    assign in5066_2 = {pp14[38]};
    Full_Adder FA_5066(s5066, c5066, in5066_1, in5066_2, pp12[40]);
    wire[0:0] s5067, in5067_1, in5067_2;
    wire c5067;
    assign in5067_1 = {pp16[36]};
    assign in5067_2 = {pp17[35]};
    Full_Adder FA_5067(s5067, c5067, in5067_1, in5067_2, pp15[37]);
    wire[0:0] s5068, in5068_1, in5068_2;
    wire c5068;
    assign in5068_1 = {pp19[33]};
    assign in5068_2 = {pp20[32]};
    Full_Adder FA_5068(s5068, c5068, in5068_1, in5068_2, pp18[34]);
    wire[0:0] s5069, in5069_1, in5069_2;
    wire c5069;
    assign in5069_1 = {pp22[30]};
    assign in5069_2 = {pp23[29]};
    Full_Adder FA_5069(s5069, c5069, in5069_1, in5069_2, pp21[31]);
    wire[0:0] s5070, in5070_1, in5070_2;
    wire c5070;
    assign in5070_1 = {pp25[27]};
    assign in5070_2 = {pp26[26]};
    Full_Adder FA_5070(s5070, c5070, in5070_1, in5070_2, pp24[28]);
    wire[0:0] s5071, in5071_1, in5071_2;
    wire c5071;
    assign in5071_1 = {pp28[24]};
    assign in5071_2 = {pp29[23]};
    Full_Adder FA_5071(s5071, c5071, in5071_1, in5071_2, pp27[25]);
    wire[0:0] s5072, in5072_1, in5072_2;
    wire c5072;
    assign in5072_1 = {pp31[21]};
    assign in5072_2 = {pp32[20]};
    Full_Adder FA_5072(s5072, c5072, in5072_1, in5072_2, pp30[22]);
    wire[0:0] s5073, in5073_1, in5073_2;
    wire c5073;
    assign in5073_1 = {pp34[18]};
    assign in5073_2 = {pp35[17]};
    Full_Adder FA_5073(s5073, c5073, in5073_1, in5073_2, pp33[19]);
    wire[0:0] s5074, in5074_1, in5074_2;
    wire c5074;
    assign in5074_1 = {pp37[15]};
    assign in5074_2 = {pp38[14]};
    Full_Adder FA_5074(s5074, c5074, in5074_1, in5074_2, pp36[16]);
    wire[0:0] s5075, in5075_1, in5075_2;
    wire c5075;
    assign in5075_1 = {pp39[13]};
    assign in5075_2 = {pp40[12]};
    Half_Adder HA_5075(s5075, c5075, in5075_1, in5075_2);
    wire[0:0] s5076, in5076_1, in5076_2;
    wire c5076;
    assign in5076_1 = {pp1[52]};
    assign in5076_2 = {pp2[51]};
    Full_Adder FA_5076(s5076, c5076, in5076_1, in5076_2, pp0[53]);
    wire[0:0] s5077, in5077_1, in5077_2;
    wire c5077;
    assign in5077_1 = {pp4[49]};
    assign in5077_2 = {pp5[48]};
    Full_Adder FA_5077(s5077, c5077, in5077_1, in5077_2, pp3[50]);
    wire[0:0] s5078, in5078_1, in5078_2;
    wire c5078;
    assign in5078_1 = {pp7[46]};
    assign in5078_2 = {pp8[45]};
    Full_Adder FA_5078(s5078, c5078, in5078_1, in5078_2, pp6[47]);
    wire[0:0] s5079, in5079_1, in5079_2;
    wire c5079;
    assign in5079_1 = {pp10[43]};
    assign in5079_2 = {pp11[42]};
    Full_Adder FA_5079(s5079, c5079, in5079_1, in5079_2, pp9[44]);
    wire[0:0] s5080, in5080_1, in5080_2;
    wire c5080;
    assign in5080_1 = {pp13[40]};
    assign in5080_2 = {pp14[39]};
    Full_Adder FA_5080(s5080, c5080, in5080_1, in5080_2, pp12[41]);
    wire[0:0] s5081, in5081_1, in5081_2;
    wire c5081;
    assign in5081_1 = {pp16[37]};
    assign in5081_2 = {pp17[36]};
    Full_Adder FA_5081(s5081, c5081, in5081_1, in5081_2, pp15[38]);
    wire[0:0] s5082, in5082_1, in5082_2;
    wire c5082;
    assign in5082_1 = {pp19[34]};
    assign in5082_2 = {pp20[33]};
    Full_Adder FA_5082(s5082, c5082, in5082_1, in5082_2, pp18[35]);
    wire[0:0] s5083, in5083_1, in5083_2;
    wire c5083;
    assign in5083_1 = {pp22[31]};
    assign in5083_2 = {pp23[30]};
    Full_Adder FA_5083(s5083, c5083, in5083_1, in5083_2, pp21[32]);
    wire[0:0] s5084, in5084_1, in5084_2;
    wire c5084;
    assign in5084_1 = {pp25[28]};
    assign in5084_2 = {pp26[27]};
    Full_Adder FA_5084(s5084, c5084, in5084_1, in5084_2, pp24[29]);
    wire[0:0] s5085, in5085_1, in5085_2;
    wire c5085;
    assign in5085_1 = {pp28[25]};
    assign in5085_2 = {pp29[24]};
    Full_Adder FA_5085(s5085, c5085, in5085_1, in5085_2, pp27[26]);
    wire[0:0] s5086, in5086_1, in5086_2;
    wire c5086;
    assign in5086_1 = {pp31[22]};
    assign in5086_2 = {pp32[21]};
    Full_Adder FA_5086(s5086, c5086, in5086_1, in5086_2, pp30[23]);
    wire[0:0] s5087, in5087_1, in5087_2;
    wire c5087;
    assign in5087_1 = {pp34[19]};
    assign in5087_2 = {pp35[18]};
    Full_Adder FA_5087(s5087, c5087, in5087_1, in5087_2, pp33[20]);
    wire[0:0] s5088, in5088_1, in5088_2;
    wire c5088;
    assign in5088_1 = {pp37[16]};
    assign in5088_2 = {pp38[15]};
    Full_Adder FA_5088(s5088, c5088, in5088_1, in5088_2, pp36[17]);
    wire[0:0] s5089, in5089_1, in5089_2;
    wire c5089;
    assign in5089_1 = {pp40[13]};
    assign in5089_2 = {pp41[12]};
    Full_Adder FA_5089(s5089, c5089, in5089_1, in5089_2, pp39[14]);
    wire[0:0] s5090, in5090_1, in5090_2;
    wire c5090;
    assign in5090_1 = {pp42[11]};
    assign in5090_2 = {pp43[10]};
    Half_Adder HA_5090(s5090, c5090, in5090_1, in5090_2);
    wire[0:0] s5091, in5091_1, in5091_2;
    wire c5091;
    assign in5091_1 = {pp1[53]};
    assign in5091_2 = {pp2[52]};
    Full_Adder FA_5091(s5091, c5091, in5091_1, in5091_2, pp0[54]);
    wire[0:0] s5092, in5092_1, in5092_2;
    wire c5092;
    assign in5092_1 = {pp4[50]};
    assign in5092_2 = {pp5[49]};
    Full_Adder FA_5092(s5092, c5092, in5092_1, in5092_2, pp3[51]);
    wire[0:0] s5093, in5093_1, in5093_2;
    wire c5093;
    assign in5093_1 = {pp7[47]};
    assign in5093_2 = {pp8[46]};
    Full_Adder FA_5093(s5093, c5093, in5093_1, in5093_2, pp6[48]);
    wire[0:0] s5094, in5094_1, in5094_2;
    wire c5094;
    assign in5094_1 = {pp10[44]};
    assign in5094_2 = {pp11[43]};
    Full_Adder FA_5094(s5094, c5094, in5094_1, in5094_2, pp9[45]);
    wire[0:0] s5095, in5095_1, in5095_2;
    wire c5095;
    assign in5095_1 = {pp13[41]};
    assign in5095_2 = {pp14[40]};
    Full_Adder FA_5095(s5095, c5095, in5095_1, in5095_2, pp12[42]);
    wire[0:0] s5096, in5096_1, in5096_2;
    wire c5096;
    assign in5096_1 = {pp16[38]};
    assign in5096_2 = {pp17[37]};
    Full_Adder FA_5096(s5096, c5096, in5096_1, in5096_2, pp15[39]);
    wire[0:0] s5097, in5097_1, in5097_2;
    wire c5097;
    assign in5097_1 = {pp19[35]};
    assign in5097_2 = {pp20[34]};
    Full_Adder FA_5097(s5097, c5097, in5097_1, in5097_2, pp18[36]);
    wire[0:0] s5098, in5098_1, in5098_2;
    wire c5098;
    assign in5098_1 = {pp22[32]};
    assign in5098_2 = {pp23[31]};
    Full_Adder FA_5098(s5098, c5098, in5098_1, in5098_2, pp21[33]);
    wire[0:0] s5099, in5099_1, in5099_2;
    wire c5099;
    assign in5099_1 = {pp25[29]};
    assign in5099_2 = {pp26[28]};
    Full_Adder FA_5099(s5099, c5099, in5099_1, in5099_2, pp24[30]);
    wire[0:0] s5100, in5100_1, in5100_2;
    wire c5100;
    assign in5100_1 = {pp28[26]};
    assign in5100_2 = {pp29[25]};
    Full_Adder FA_5100(s5100, c5100, in5100_1, in5100_2, pp27[27]);
    wire[0:0] s5101, in5101_1, in5101_2;
    wire c5101;
    assign in5101_1 = {pp31[23]};
    assign in5101_2 = {pp32[22]};
    Full_Adder FA_5101(s5101, c5101, in5101_1, in5101_2, pp30[24]);
    wire[0:0] s5102, in5102_1, in5102_2;
    wire c5102;
    assign in5102_1 = {pp34[20]};
    assign in5102_2 = {pp35[19]};
    Full_Adder FA_5102(s5102, c5102, in5102_1, in5102_2, pp33[21]);
    wire[0:0] s5103, in5103_1, in5103_2;
    wire c5103;
    assign in5103_1 = {pp37[17]};
    assign in5103_2 = {pp38[16]};
    Full_Adder FA_5103(s5103, c5103, in5103_1, in5103_2, pp36[18]);
    wire[0:0] s5104, in5104_1, in5104_2;
    wire c5104;
    assign in5104_1 = {pp40[14]};
    assign in5104_2 = {pp41[13]};
    Full_Adder FA_5104(s5104, c5104, in5104_1, in5104_2, pp39[15]);
    wire[0:0] s5105, in5105_1, in5105_2;
    wire c5105;
    assign in5105_1 = {pp43[11]};
    assign in5105_2 = {pp44[10]};
    Full_Adder FA_5105(s5105, c5105, in5105_1, in5105_2, pp42[12]);
    wire[0:0] s5106, in5106_1, in5106_2;
    wire c5106;
    assign in5106_1 = {pp45[9]};
    assign in5106_2 = {pp46[8]};
    Half_Adder HA_5106(s5106, c5106, in5106_1, in5106_2);
    wire[0:0] s5107, in5107_1, in5107_2;
    wire c5107;
    assign in5107_1 = {pp1[54]};
    assign in5107_2 = {pp2[53]};
    Full_Adder FA_5107(s5107, c5107, in5107_1, in5107_2, pp0[55]);
    wire[0:0] s5108, in5108_1, in5108_2;
    wire c5108;
    assign in5108_1 = {pp4[51]};
    assign in5108_2 = {pp5[50]};
    Full_Adder FA_5108(s5108, c5108, in5108_1, in5108_2, pp3[52]);
    wire[0:0] s5109, in5109_1, in5109_2;
    wire c5109;
    assign in5109_1 = {pp7[48]};
    assign in5109_2 = {pp8[47]};
    Full_Adder FA_5109(s5109, c5109, in5109_1, in5109_2, pp6[49]);
    wire[0:0] s5110, in5110_1, in5110_2;
    wire c5110;
    assign in5110_1 = {pp10[45]};
    assign in5110_2 = {pp11[44]};
    Full_Adder FA_5110(s5110, c5110, in5110_1, in5110_2, pp9[46]);
    wire[0:0] s5111, in5111_1, in5111_2;
    wire c5111;
    assign in5111_1 = {pp13[42]};
    assign in5111_2 = {pp14[41]};
    Full_Adder FA_5111(s5111, c5111, in5111_1, in5111_2, pp12[43]);
    wire[0:0] s5112, in5112_1, in5112_2;
    wire c5112;
    assign in5112_1 = {pp16[39]};
    assign in5112_2 = {pp17[38]};
    Full_Adder FA_5112(s5112, c5112, in5112_1, in5112_2, pp15[40]);
    wire[0:0] s5113, in5113_1, in5113_2;
    wire c5113;
    assign in5113_1 = {pp19[36]};
    assign in5113_2 = {pp20[35]};
    Full_Adder FA_5113(s5113, c5113, in5113_1, in5113_2, pp18[37]);
    wire[0:0] s5114, in5114_1, in5114_2;
    wire c5114;
    assign in5114_1 = {pp22[33]};
    assign in5114_2 = {pp23[32]};
    Full_Adder FA_5114(s5114, c5114, in5114_1, in5114_2, pp21[34]);
    wire[0:0] s5115, in5115_1, in5115_2;
    wire c5115;
    assign in5115_1 = {pp25[30]};
    assign in5115_2 = {pp26[29]};
    Full_Adder FA_5115(s5115, c5115, in5115_1, in5115_2, pp24[31]);
    wire[0:0] s5116, in5116_1, in5116_2;
    wire c5116;
    assign in5116_1 = {pp28[27]};
    assign in5116_2 = {pp29[26]};
    Full_Adder FA_5116(s5116, c5116, in5116_1, in5116_2, pp27[28]);
    wire[0:0] s5117, in5117_1, in5117_2;
    wire c5117;
    assign in5117_1 = {pp31[24]};
    assign in5117_2 = {pp32[23]};
    Full_Adder FA_5117(s5117, c5117, in5117_1, in5117_2, pp30[25]);
    wire[0:0] s5118, in5118_1, in5118_2;
    wire c5118;
    assign in5118_1 = {pp34[21]};
    assign in5118_2 = {pp35[20]};
    Full_Adder FA_5118(s5118, c5118, in5118_1, in5118_2, pp33[22]);
    wire[0:0] s5119, in5119_1, in5119_2;
    wire c5119;
    assign in5119_1 = {pp37[18]};
    assign in5119_2 = {pp38[17]};
    Full_Adder FA_5119(s5119, c5119, in5119_1, in5119_2, pp36[19]);
    wire[0:0] s5120, in5120_1, in5120_2;
    wire c5120;
    assign in5120_1 = {pp40[15]};
    assign in5120_2 = {pp41[14]};
    Full_Adder FA_5120(s5120, c5120, in5120_1, in5120_2, pp39[16]);
    wire[0:0] s5121, in5121_1, in5121_2;
    wire c5121;
    assign in5121_1 = {pp43[12]};
    assign in5121_2 = {pp44[11]};
    Full_Adder FA_5121(s5121, c5121, in5121_1, in5121_2, pp42[13]);
    wire[0:0] s5122, in5122_1, in5122_2;
    wire c5122;
    assign in5122_1 = {pp46[9]};
    assign in5122_2 = {pp47[8]};
    Full_Adder FA_5122(s5122, c5122, in5122_1, in5122_2, pp45[10]);
    wire[0:0] s5123, in5123_1, in5123_2;
    wire c5123;
    assign in5123_1 = {pp48[7]};
    assign in5123_2 = {pp49[6]};
    Half_Adder HA_5123(s5123, c5123, in5123_1, in5123_2);
    wire[0:0] s5124, in5124_1, in5124_2;
    wire c5124;
    assign in5124_1 = {pp1[55]};
    assign in5124_2 = {pp2[54]};
    Full_Adder FA_5124(s5124, c5124, in5124_1, in5124_2, pp0[56]);
    wire[0:0] s5125, in5125_1, in5125_2;
    wire c5125;
    assign in5125_1 = {pp4[52]};
    assign in5125_2 = {pp5[51]};
    Full_Adder FA_5125(s5125, c5125, in5125_1, in5125_2, pp3[53]);
    wire[0:0] s5126, in5126_1, in5126_2;
    wire c5126;
    assign in5126_1 = {pp7[49]};
    assign in5126_2 = {pp8[48]};
    Full_Adder FA_5126(s5126, c5126, in5126_1, in5126_2, pp6[50]);
    wire[0:0] s5127, in5127_1, in5127_2;
    wire c5127;
    assign in5127_1 = {pp10[46]};
    assign in5127_2 = {pp11[45]};
    Full_Adder FA_5127(s5127, c5127, in5127_1, in5127_2, pp9[47]);
    wire[0:0] s5128, in5128_1, in5128_2;
    wire c5128;
    assign in5128_1 = {pp13[43]};
    assign in5128_2 = {pp14[42]};
    Full_Adder FA_5128(s5128, c5128, in5128_1, in5128_2, pp12[44]);
    wire[0:0] s5129, in5129_1, in5129_2;
    wire c5129;
    assign in5129_1 = {pp16[40]};
    assign in5129_2 = {pp17[39]};
    Full_Adder FA_5129(s5129, c5129, in5129_1, in5129_2, pp15[41]);
    wire[0:0] s5130, in5130_1, in5130_2;
    wire c5130;
    assign in5130_1 = {pp19[37]};
    assign in5130_2 = {pp20[36]};
    Full_Adder FA_5130(s5130, c5130, in5130_1, in5130_2, pp18[38]);
    wire[0:0] s5131, in5131_1, in5131_2;
    wire c5131;
    assign in5131_1 = {pp22[34]};
    assign in5131_2 = {pp23[33]};
    Full_Adder FA_5131(s5131, c5131, in5131_1, in5131_2, pp21[35]);
    wire[0:0] s5132, in5132_1, in5132_2;
    wire c5132;
    assign in5132_1 = {pp25[31]};
    assign in5132_2 = {pp26[30]};
    Full_Adder FA_5132(s5132, c5132, in5132_1, in5132_2, pp24[32]);
    wire[0:0] s5133, in5133_1, in5133_2;
    wire c5133;
    assign in5133_1 = {pp28[28]};
    assign in5133_2 = {pp29[27]};
    Full_Adder FA_5133(s5133, c5133, in5133_1, in5133_2, pp27[29]);
    wire[0:0] s5134, in5134_1, in5134_2;
    wire c5134;
    assign in5134_1 = {pp31[25]};
    assign in5134_2 = {pp32[24]};
    Full_Adder FA_5134(s5134, c5134, in5134_1, in5134_2, pp30[26]);
    wire[0:0] s5135, in5135_1, in5135_2;
    wire c5135;
    assign in5135_1 = {pp34[22]};
    assign in5135_2 = {pp35[21]};
    Full_Adder FA_5135(s5135, c5135, in5135_1, in5135_2, pp33[23]);
    wire[0:0] s5136, in5136_1, in5136_2;
    wire c5136;
    assign in5136_1 = {pp37[19]};
    assign in5136_2 = {pp38[18]};
    Full_Adder FA_5136(s5136, c5136, in5136_1, in5136_2, pp36[20]);
    wire[0:0] s5137, in5137_1, in5137_2;
    wire c5137;
    assign in5137_1 = {pp40[16]};
    assign in5137_2 = {pp41[15]};
    Full_Adder FA_5137(s5137, c5137, in5137_1, in5137_2, pp39[17]);
    wire[0:0] s5138, in5138_1, in5138_2;
    wire c5138;
    assign in5138_1 = {pp43[13]};
    assign in5138_2 = {pp44[12]};
    Full_Adder FA_5138(s5138, c5138, in5138_1, in5138_2, pp42[14]);
    wire[0:0] s5139, in5139_1, in5139_2;
    wire c5139;
    assign in5139_1 = {pp46[10]};
    assign in5139_2 = {pp47[9]};
    Full_Adder FA_5139(s5139, c5139, in5139_1, in5139_2, pp45[11]);
    wire[0:0] s5140, in5140_1, in5140_2;
    wire c5140;
    assign in5140_1 = {pp49[7]};
    assign in5140_2 = {pp50[6]};
    Full_Adder FA_5140(s5140, c5140, in5140_1, in5140_2, pp48[8]);
    wire[0:0] s5141, in5141_1, in5141_2;
    wire c5141;
    assign in5141_1 = {pp51[5]};
    assign in5141_2 = {pp52[4]};
    Half_Adder HA_5141(s5141, c5141, in5141_1, in5141_2);
    wire[0:0] s5142, in5142_1, in5142_2;
    wire c5142;
    assign in5142_1 = {pp1[56]};
    assign in5142_2 = {pp2[55]};
    Full_Adder FA_5142(s5142, c5142, in5142_1, in5142_2, pp0[57]);
    wire[0:0] s5143, in5143_1, in5143_2;
    wire c5143;
    assign in5143_1 = {pp4[53]};
    assign in5143_2 = {pp5[52]};
    Full_Adder FA_5143(s5143, c5143, in5143_1, in5143_2, pp3[54]);
    wire[0:0] s5144, in5144_1, in5144_2;
    wire c5144;
    assign in5144_1 = {pp7[50]};
    assign in5144_2 = {pp8[49]};
    Full_Adder FA_5144(s5144, c5144, in5144_1, in5144_2, pp6[51]);
    wire[0:0] s5145, in5145_1, in5145_2;
    wire c5145;
    assign in5145_1 = {pp10[47]};
    assign in5145_2 = {pp11[46]};
    Full_Adder FA_5145(s5145, c5145, in5145_1, in5145_2, pp9[48]);
    wire[0:0] s5146, in5146_1, in5146_2;
    wire c5146;
    assign in5146_1 = {pp13[44]};
    assign in5146_2 = {pp14[43]};
    Full_Adder FA_5146(s5146, c5146, in5146_1, in5146_2, pp12[45]);
    wire[0:0] s5147, in5147_1, in5147_2;
    wire c5147;
    assign in5147_1 = {pp16[41]};
    assign in5147_2 = {pp17[40]};
    Full_Adder FA_5147(s5147, c5147, in5147_1, in5147_2, pp15[42]);
    wire[0:0] s5148, in5148_1, in5148_2;
    wire c5148;
    assign in5148_1 = {pp19[38]};
    assign in5148_2 = {pp20[37]};
    Full_Adder FA_5148(s5148, c5148, in5148_1, in5148_2, pp18[39]);
    wire[0:0] s5149, in5149_1, in5149_2;
    wire c5149;
    assign in5149_1 = {pp22[35]};
    assign in5149_2 = {pp23[34]};
    Full_Adder FA_5149(s5149, c5149, in5149_1, in5149_2, pp21[36]);
    wire[0:0] s5150, in5150_1, in5150_2;
    wire c5150;
    assign in5150_1 = {pp25[32]};
    assign in5150_2 = {pp26[31]};
    Full_Adder FA_5150(s5150, c5150, in5150_1, in5150_2, pp24[33]);
    wire[0:0] s5151, in5151_1, in5151_2;
    wire c5151;
    assign in5151_1 = {pp28[29]};
    assign in5151_2 = {pp29[28]};
    Full_Adder FA_5151(s5151, c5151, in5151_1, in5151_2, pp27[30]);
    wire[0:0] s5152, in5152_1, in5152_2;
    wire c5152;
    assign in5152_1 = {pp31[26]};
    assign in5152_2 = {pp32[25]};
    Full_Adder FA_5152(s5152, c5152, in5152_1, in5152_2, pp30[27]);
    wire[0:0] s5153, in5153_1, in5153_2;
    wire c5153;
    assign in5153_1 = {pp34[23]};
    assign in5153_2 = {pp35[22]};
    Full_Adder FA_5153(s5153, c5153, in5153_1, in5153_2, pp33[24]);
    wire[0:0] s5154, in5154_1, in5154_2;
    wire c5154;
    assign in5154_1 = {pp37[20]};
    assign in5154_2 = {pp38[19]};
    Full_Adder FA_5154(s5154, c5154, in5154_1, in5154_2, pp36[21]);
    wire[0:0] s5155, in5155_1, in5155_2;
    wire c5155;
    assign in5155_1 = {pp40[17]};
    assign in5155_2 = {pp41[16]};
    Full_Adder FA_5155(s5155, c5155, in5155_1, in5155_2, pp39[18]);
    wire[0:0] s5156, in5156_1, in5156_2;
    wire c5156;
    assign in5156_1 = {pp43[14]};
    assign in5156_2 = {pp44[13]};
    Full_Adder FA_5156(s5156, c5156, in5156_1, in5156_2, pp42[15]);
    wire[0:0] s5157, in5157_1, in5157_2;
    wire c5157;
    assign in5157_1 = {pp46[11]};
    assign in5157_2 = {pp47[10]};
    Full_Adder FA_5157(s5157, c5157, in5157_1, in5157_2, pp45[12]);
    wire[0:0] s5158, in5158_1, in5158_2;
    wire c5158;
    assign in5158_1 = {pp49[8]};
    assign in5158_2 = {pp50[7]};
    Full_Adder FA_5158(s5158, c5158, in5158_1, in5158_2, pp48[9]);
    wire[0:0] s5159, in5159_1, in5159_2;
    wire c5159;
    assign in5159_1 = {pp52[5]};
    assign in5159_2 = {pp53[4]};
    Full_Adder FA_5159(s5159, c5159, in5159_1, in5159_2, pp51[6]);
    wire[0:0] s5160, in5160_1, in5160_2;
    wire c5160;
    assign in5160_1 = {pp54[3]};
    assign in5160_2 = {pp55[2]};
    Half_Adder HA_5160(s5160, c5160, in5160_1, in5160_2);
    wire[0:0] s5161, in5161_1, in5161_2;
    wire c5161;
    assign in5161_1 = {pp3[55]};
    assign in5161_2 = {pp4[54]};
    Full_Adder FA_5161(s5161, c5161, in5161_1, in5161_2, pp2[56]);
    wire[0:0] s5162, in5162_1, in5162_2;
    wire c5162;
    assign in5162_1 = {pp6[52]};
    assign in5162_2 = {pp7[51]};
    Full_Adder FA_5162(s5162, c5162, in5162_1, in5162_2, pp5[53]);
    wire[0:0] s5163, in5163_1, in5163_2;
    wire c5163;
    assign in5163_1 = {pp9[49]};
    assign in5163_2 = {pp10[48]};
    Full_Adder FA_5163(s5163, c5163, in5163_1, in5163_2, pp8[50]);
    wire[0:0] s5164, in5164_1, in5164_2;
    wire c5164;
    assign in5164_1 = {pp12[46]};
    assign in5164_2 = {pp13[45]};
    Full_Adder FA_5164(s5164, c5164, in5164_1, in5164_2, pp11[47]);
    wire[0:0] s5165, in5165_1, in5165_2;
    wire c5165;
    assign in5165_1 = {pp15[43]};
    assign in5165_2 = {pp16[42]};
    Full_Adder FA_5165(s5165, c5165, in5165_1, in5165_2, pp14[44]);
    wire[0:0] s5166, in5166_1, in5166_2;
    wire c5166;
    assign in5166_1 = {pp18[40]};
    assign in5166_2 = {pp19[39]};
    Full_Adder FA_5166(s5166, c5166, in5166_1, in5166_2, pp17[41]);
    wire[0:0] s5167, in5167_1, in5167_2;
    wire c5167;
    assign in5167_1 = {pp21[37]};
    assign in5167_2 = {pp22[36]};
    Full_Adder FA_5167(s5167, c5167, in5167_1, in5167_2, pp20[38]);
    wire[0:0] s5168, in5168_1, in5168_2;
    wire c5168;
    assign in5168_1 = {pp24[34]};
    assign in5168_2 = {pp25[33]};
    Full_Adder FA_5168(s5168, c5168, in5168_1, in5168_2, pp23[35]);
    wire[0:0] s5169, in5169_1, in5169_2;
    wire c5169;
    assign in5169_1 = {pp27[31]};
    assign in5169_2 = {pp28[30]};
    Full_Adder FA_5169(s5169, c5169, in5169_1, in5169_2, pp26[32]);
    wire[0:0] s5170, in5170_1, in5170_2;
    wire c5170;
    assign in5170_1 = {pp30[28]};
    assign in5170_2 = {pp31[27]};
    Full_Adder FA_5170(s5170, c5170, in5170_1, in5170_2, pp29[29]);
    wire[0:0] s5171, in5171_1, in5171_2;
    wire c5171;
    assign in5171_1 = {pp33[25]};
    assign in5171_2 = {pp34[24]};
    Full_Adder FA_5171(s5171, c5171, in5171_1, in5171_2, pp32[26]);
    wire[0:0] s5172, in5172_1, in5172_2;
    wire c5172;
    assign in5172_1 = {pp36[22]};
    assign in5172_2 = {pp37[21]};
    Full_Adder FA_5172(s5172, c5172, in5172_1, in5172_2, pp35[23]);
    wire[0:0] s5173, in5173_1, in5173_2;
    wire c5173;
    assign in5173_1 = {pp39[19]};
    assign in5173_2 = {pp40[18]};
    Full_Adder FA_5173(s5173, c5173, in5173_1, in5173_2, pp38[20]);
    wire[0:0] s5174, in5174_1, in5174_2;
    wire c5174;
    assign in5174_1 = {pp42[16]};
    assign in5174_2 = {pp43[15]};
    Full_Adder FA_5174(s5174, c5174, in5174_1, in5174_2, pp41[17]);
    wire[0:0] s5175, in5175_1, in5175_2;
    wire c5175;
    assign in5175_1 = {pp45[13]};
    assign in5175_2 = {pp46[12]};
    Full_Adder FA_5175(s5175, c5175, in5175_1, in5175_2, pp44[14]);
    wire[0:0] s5176, in5176_1, in5176_2;
    wire c5176;
    assign in5176_1 = {pp48[10]};
    assign in5176_2 = {pp49[9]};
    Full_Adder FA_5176(s5176, c5176, in5176_1, in5176_2, pp47[11]);
    wire[0:0] s5177, in5177_1, in5177_2;
    wire c5177;
    assign in5177_1 = {pp51[7]};
    assign in5177_2 = {pp52[6]};
    Full_Adder FA_5177(s5177, c5177, in5177_1, in5177_2, pp50[8]);
    wire[0:0] s5178, in5178_1, in5178_2;
    wire c5178;
    assign in5178_1 = {pp54[4]};
    assign in5178_2 = {pp55[3]};
    Full_Adder FA_5178(s5178, c5178, in5178_1, in5178_2, pp53[5]);
    wire[0:0] s5179, in5179_1, in5179_2;
    wire c5179;
    assign in5179_1 = {pp57[1]};
    assign in5179_2 = {pp58[0]};
    Full_Adder FA_5179(s5179, c5179, in5179_1, in5179_2, pp56[2]);
    wire[0:0] s5180, in5180_1, in5180_2;
    wire c5180;
    assign in5180_1 = {pp6[53]};
    assign in5180_2 = {pp7[52]};
    Full_Adder FA_5180(s5180, c5180, in5180_1, in5180_2, pp5[54]);
    wire[0:0] s5181, in5181_1, in5181_2;
    wire c5181;
    assign in5181_1 = {pp9[50]};
    assign in5181_2 = {pp10[49]};
    Full_Adder FA_5181(s5181, c5181, in5181_1, in5181_2, pp8[51]);
    wire[0:0] s5182, in5182_1, in5182_2;
    wire c5182;
    assign in5182_1 = {pp12[47]};
    assign in5182_2 = {pp13[46]};
    Full_Adder FA_5182(s5182, c5182, in5182_1, in5182_2, pp11[48]);
    wire[0:0] s5183, in5183_1, in5183_2;
    wire c5183;
    assign in5183_1 = {pp15[44]};
    assign in5183_2 = {pp16[43]};
    Full_Adder FA_5183(s5183, c5183, in5183_1, in5183_2, pp14[45]);
    wire[0:0] s5184, in5184_1, in5184_2;
    wire c5184;
    assign in5184_1 = {pp18[41]};
    assign in5184_2 = {pp19[40]};
    Full_Adder FA_5184(s5184, c5184, in5184_1, in5184_2, pp17[42]);
    wire[0:0] s5185, in5185_1, in5185_2;
    wire c5185;
    assign in5185_1 = {pp21[38]};
    assign in5185_2 = {pp22[37]};
    Full_Adder FA_5185(s5185, c5185, in5185_1, in5185_2, pp20[39]);
    wire[0:0] s5186, in5186_1, in5186_2;
    wire c5186;
    assign in5186_1 = {pp24[35]};
    assign in5186_2 = {pp25[34]};
    Full_Adder FA_5186(s5186, c5186, in5186_1, in5186_2, pp23[36]);
    wire[0:0] s5187, in5187_1, in5187_2;
    wire c5187;
    assign in5187_1 = {pp27[32]};
    assign in5187_2 = {pp28[31]};
    Full_Adder FA_5187(s5187, c5187, in5187_1, in5187_2, pp26[33]);
    wire[0:0] s5188, in5188_1, in5188_2;
    wire c5188;
    assign in5188_1 = {pp30[29]};
    assign in5188_2 = {pp31[28]};
    Full_Adder FA_5188(s5188, c5188, in5188_1, in5188_2, pp29[30]);
    wire[0:0] s5189, in5189_1, in5189_2;
    wire c5189;
    assign in5189_1 = {pp33[26]};
    assign in5189_2 = {pp34[25]};
    Full_Adder FA_5189(s5189, c5189, in5189_1, in5189_2, pp32[27]);
    wire[0:0] s5190, in5190_1, in5190_2;
    wire c5190;
    assign in5190_1 = {pp36[23]};
    assign in5190_2 = {pp37[22]};
    Full_Adder FA_5190(s5190, c5190, in5190_1, in5190_2, pp35[24]);
    wire[0:0] s5191, in5191_1, in5191_2;
    wire c5191;
    assign in5191_1 = {pp39[20]};
    assign in5191_2 = {pp40[19]};
    Full_Adder FA_5191(s5191, c5191, in5191_1, in5191_2, pp38[21]);
    wire[0:0] s5192, in5192_1, in5192_2;
    wire c5192;
    assign in5192_1 = {pp42[17]};
    assign in5192_2 = {pp43[16]};
    Full_Adder FA_5192(s5192, c5192, in5192_1, in5192_2, pp41[18]);
    wire[0:0] s5193, in5193_1, in5193_2;
    wire c5193;
    assign in5193_1 = {pp45[14]};
    assign in5193_2 = {pp46[13]};
    Full_Adder FA_5193(s5193, c5193, in5193_1, in5193_2, pp44[15]);
    wire[0:0] s5194, in5194_1, in5194_2;
    wire c5194;
    assign in5194_1 = {pp48[11]};
    assign in5194_2 = {pp49[10]};
    Full_Adder FA_5194(s5194, c5194, in5194_1, in5194_2, pp47[12]);
    wire[0:0] s5195, in5195_1, in5195_2;
    wire c5195;
    assign in5195_1 = {pp51[8]};
    assign in5195_2 = {pp52[7]};
    Full_Adder FA_5195(s5195, c5195, in5195_1, in5195_2, pp50[9]);
    wire[0:0] s5196, in5196_1, in5196_2;
    wire c5196;
    assign in5196_1 = {pp54[5]};
    assign in5196_2 = {pp55[4]};
    Full_Adder FA_5196(s5196, c5196, in5196_1, in5196_2, pp53[6]);
    wire[0:0] s5197, in5197_1, in5197_2;
    wire c5197;
    assign in5197_1 = {pp57[2]};
    assign in5197_2 = {pp58[1]};
    Full_Adder FA_5197(s5197, c5197, in5197_1, in5197_2, pp56[3]);
    wire[0:0] s5198, in5198_1, in5198_2;
    wire c5198;
    assign in5198_1 = {c1807};
    assign in5198_2 = {s1808[0]};
    Full_Adder FA_5198(s5198, c5198, in5198_1, in5198_2, pp59[0]);
    wire[0:0] s5199, in5199_1, in5199_2;
    wire c5199;
    assign in5199_1 = {pp9[51]};
    assign in5199_2 = {pp10[50]};
    Full_Adder FA_5199(s5199, c5199, in5199_1, in5199_2, pp8[52]);
    wire[0:0] s5200, in5200_1, in5200_2;
    wire c5200;
    assign in5200_1 = {pp12[48]};
    assign in5200_2 = {pp13[47]};
    Full_Adder FA_5200(s5200, c5200, in5200_1, in5200_2, pp11[49]);
    wire[0:0] s5201, in5201_1, in5201_2;
    wire c5201;
    assign in5201_1 = {pp15[45]};
    assign in5201_2 = {pp16[44]};
    Full_Adder FA_5201(s5201, c5201, in5201_1, in5201_2, pp14[46]);
    wire[0:0] s5202, in5202_1, in5202_2;
    wire c5202;
    assign in5202_1 = {pp18[42]};
    assign in5202_2 = {pp19[41]};
    Full_Adder FA_5202(s5202, c5202, in5202_1, in5202_2, pp17[43]);
    wire[0:0] s5203, in5203_1, in5203_2;
    wire c5203;
    assign in5203_1 = {pp21[39]};
    assign in5203_2 = {pp22[38]};
    Full_Adder FA_5203(s5203, c5203, in5203_1, in5203_2, pp20[40]);
    wire[0:0] s5204, in5204_1, in5204_2;
    wire c5204;
    assign in5204_1 = {pp24[36]};
    assign in5204_2 = {pp25[35]};
    Full_Adder FA_5204(s5204, c5204, in5204_1, in5204_2, pp23[37]);
    wire[0:0] s5205, in5205_1, in5205_2;
    wire c5205;
    assign in5205_1 = {pp27[33]};
    assign in5205_2 = {pp28[32]};
    Full_Adder FA_5205(s5205, c5205, in5205_1, in5205_2, pp26[34]);
    wire[0:0] s5206, in5206_1, in5206_2;
    wire c5206;
    assign in5206_1 = {pp30[30]};
    assign in5206_2 = {pp31[29]};
    Full_Adder FA_5206(s5206, c5206, in5206_1, in5206_2, pp29[31]);
    wire[0:0] s5207, in5207_1, in5207_2;
    wire c5207;
    assign in5207_1 = {pp33[27]};
    assign in5207_2 = {pp34[26]};
    Full_Adder FA_5207(s5207, c5207, in5207_1, in5207_2, pp32[28]);
    wire[0:0] s5208, in5208_1, in5208_2;
    wire c5208;
    assign in5208_1 = {pp36[24]};
    assign in5208_2 = {pp37[23]};
    Full_Adder FA_5208(s5208, c5208, in5208_1, in5208_2, pp35[25]);
    wire[0:0] s5209, in5209_1, in5209_2;
    wire c5209;
    assign in5209_1 = {pp39[21]};
    assign in5209_2 = {pp40[20]};
    Full_Adder FA_5209(s5209, c5209, in5209_1, in5209_2, pp38[22]);
    wire[0:0] s5210, in5210_1, in5210_2;
    wire c5210;
    assign in5210_1 = {pp42[18]};
    assign in5210_2 = {pp43[17]};
    Full_Adder FA_5210(s5210, c5210, in5210_1, in5210_2, pp41[19]);
    wire[0:0] s5211, in5211_1, in5211_2;
    wire c5211;
    assign in5211_1 = {pp45[15]};
    assign in5211_2 = {pp46[14]};
    Full_Adder FA_5211(s5211, c5211, in5211_1, in5211_2, pp44[16]);
    wire[0:0] s5212, in5212_1, in5212_2;
    wire c5212;
    assign in5212_1 = {pp48[12]};
    assign in5212_2 = {pp49[11]};
    Full_Adder FA_5212(s5212, c5212, in5212_1, in5212_2, pp47[13]);
    wire[0:0] s5213, in5213_1, in5213_2;
    wire c5213;
    assign in5213_1 = {pp51[9]};
    assign in5213_2 = {pp52[8]};
    Full_Adder FA_5213(s5213, c5213, in5213_1, in5213_2, pp50[10]);
    wire[0:0] s5214, in5214_1, in5214_2;
    wire c5214;
    assign in5214_1 = {pp54[6]};
    assign in5214_2 = {pp55[5]};
    Full_Adder FA_5214(s5214, c5214, in5214_1, in5214_2, pp53[7]);
    wire[0:0] s5215, in5215_1, in5215_2;
    wire c5215;
    assign in5215_1 = {pp57[3]};
    assign in5215_2 = {pp58[2]};
    Full_Adder FA_5215(s5215, c5215, in5215_1, in5215_2, pp56[4]);
    wire[0:0] s5216, in5216_1, in5216_2;
    wire c5216;
    assign in5216_1 = {pp60[0]};
    assign in5216_2 = {c1808};
    Full_Adder FA_5216(s5216, c5216, in5216_1, in5216_2, pp59[1]);
    wire[0:0] s5217, in5217_1, in5217_2;
    wire c5217;
    assign in5217_1 = {s1810[0]};
    assign in5217_2 = {s1811[0]};
    Full_Adder FA_5217(s5217, c5217, in5217_1, in5217_2, c1809);
    wire[0:0] s5218, in5218_1, in5218_2;
    wire c5218;
    assign in5218_1 = {pp12[49]};
    assign in5218_2 = {pp13[48]};
    Full_Adder FA_5218(s5218, c5218, in5218_1, in5218_2, pp11[50]);
    wire[0:0] s5219, in5219_1, in5219_2;
    wire c5219;
    assign in5219_1 = {pp15[46]};
    assign in5219_2 = {pp16[45]};
    Full_Adder FA_5219(s5219, c5219, in5219_1, in5219_2, pp14[47]);
    wire[0:0] s5220, in5220_1, in5220_2;
    wire c5220;
    assign in5220_1 = {pp18[43]};
    assign in5220_2 = {pp19[42]};
    Full_Adder FA_5220(s5220, c5220, in5220_1, in5220_2, pp17[44]);
    wire[0:0] s5221, in5221_1, in5221_2;
    wire c5221;
    assign in5221_1 = {pp21[40]};
    assign in5221_2 = {pp22[39]};
    Full_Adder FA_5221(s5221, c5221, in5221_1, in5221_2, pp20[41]);
    wire[0:0] s5222, in5222_1, in5222_2;
    wire c5222;
    assign in5222_1 = {pp24[37]};
    assign in5222_2 = {pp25[36]};
    Full_Adder FA_5222(s5222, c5222, in5222_1, in5222_2, pp23[38]);
    wire[0:0] s5223, in5223_1, in5223_2;
    wire c5223;
    assign in5223_1 = {pp27[34]};
    assign in5223_2 = {pp28[33]};
    Full_Adder FA_5223(s5223, c5223, in5223_1, in5223_2, pp26[35]);
    wire[0:0] s5224, in5224_1, in5224_2;
    wire c5224;
    assign in5224_1 = {pp30[31]};
    assign in5224_2 = {pp31[30]};
    Full_Adder FA_5224(s5224, c5224, in5224_1, in5224_2, pp29[32]);
    wire[0:0] s5225, in5225_1, in5225_2;
    wire c5225;
    assign in5225_1 = {pp33[28]};
    assign in5225_2 = {pp34[27]};
    Full_Adder FA_5225(s5225, c5225, in5225_1, in5225_2, pp32[29]);
    wire[0:0] s5226, in5226_1, in5226_2;
    wire c5226;
    assign in5226_1 = {pp36[25]};
    assign in5226_2 = {pp37[24]};
    Full_Adder FA_5226(s5226, c5226, in5226_1, in5226_2, pp35[26]);
    wire[0:0] s5227, in5227_1, in5227_2;
    wire c5227;
    assign in5227_1 = {pp39[22]};
    assign in5227_2 = {pp40[21]};
    Full_Adder FA_5227(s5227, c5227, in5227_1, in5227_2, pp38[23]);
    wire[0:0] s5228, in5228_1, in5228_2;
    wire c5228;
    assign in5228_1 = {pp42[19]};
    assign in5228_2 = {pp43[18]};
    Full_Adder FA_5228(s5228, c5228, in5228_1, in5228_2, pp41[20]);
    wire[0:0] s5229, in5229_1, in5229_2;
    wire c5229;
    assign in5229_1 = {pp45[16]};
    assign in5229_2 = {pp46[15]};
    Full_Adder FA_5229(s5229, c5229, in5229_1, in5229_2, pp44[17]);
    wire[0:0] s5230, in5230_1, in5230_2;
    wire c5230;
    assign in5230_1 = {pp48[13]};
    assign in5230_2 = {pp49[12]};
    Full_Adder FA_5230(s5230, c5230, in5230_1, in5230_2, pp47[14]);
    wire[0:0] s5231, in5231_1, in5231_2;
    wire c5231;
    assign in5231_1 = {pp51[10]};
    assign in5231_2 = {pp52[9]};
    Full_Adder FA_5231(s5231, c5231, in5231_1, in5231_2, pp50[11]);
    wire[0:0] s5232, in5232_1, in5232_2;
    wire c5232;
    assign in5232_1 = {pp54[7]};
    assign in5232_2 = {pp55[6]};
    Full_Adder FA_5232(s5232, c5232, in5232_1, in5232_2, pp53[8]);
    wire[0:0] s5233, in5233_1, in5233_2;
    wire c5233;
    assign in5233_1 = {pp57[4]};
    assign in5233_2 = {pp58[3]};
    Full_Adder FA_5233(s5233, c5233, in5233_1, in5233_2, pp56[5]);
    wire[0:0] s5234, in5234_1, in5234_2;
    wire c5234;
    assign in5234_1 = {pp60[1]};
    assign in5234_2 = {pp61[0]};
    Full_Adder FA_5234(s5234, c5234, in5234_1, in5234_2, pp59[2]);
    wire[0:0] s5235, in5235_1, in5235_2;
    wire c5235;
    assign in5235_1 = {c1811};
    assign in5235_2 = {c1812};
    Full_Adder FA_5235(s5235, c5235, in5235_1, in5235_2, c1810);
    wire[0:0] s5236, in5236_1, in5236_2;
    wire c5236;
    assign in5236_1 = {s1814[0]};
    assign in5236_2 = {s1815[0]};
    Full_Adder FA_5236(s5236, c5236, in5236_1, in5236_2, s1813[0]);
    wire[0:0] s5237, in5237_1, in5237_2;
    wire c5237;
    assign in5237_1 = {pp15[47]};
    assign in5237_2 = {pp16[46]};
    Full_Adder FA_5237(s5237, c5237, in5237_1, in5237_2, pp14[48]);
    wire[0:0] s5238, in5238_1, in5238_2;
    wire c5238;
    assign in5238_1 = {pp18[44]};
    assign in5238_2 = {pp19[43]};
    Full_Adder FA_5238(s5238, c5238, in5238_1, in5238_2, pp17[45]);
    wire[0:0] s5239, in5239_1, in5239_2;
    wire c5239;
    assign in5239_1 = {pp21[41]};
    assign in5239_2 = {pp22[40]};
    Full_Adder FA_5239(s5239, c5239, in5239_1, in5239_2, pp20[42]);
    wire[0:0] s5240, in5240_1, in5240_2;
    wire c5240;
    assign in5240_1 = {pp24[38]};
    assign in5240_2 = {pp25[37]};
    Full_Adder FA_5240(s5240, c5240, in5240_1, in5240_2, pp23[39]);
    wire[0:0] s5241, in5241_1, in5241_2;
    wire c5241;
    assign in5241_1 = {pp27[35]};
    assign in5241_2 = {pp28[34]};
    Full_Adder FA_5241(s5241, c5241, in5241_1, in5241_2, pp26[36]);
    wire[0:0] s5242, in5242_1, in5242_2;
    wire c5242;
    assign in5242_1 = {pp30[32]};
    assign in5242_2 = {pp31[31]};
    Full_Adder FA_5242(s5242, c5242, in5242_1, in5242_2, pp29[33]);
    wire[0:0] s5243, in5243_1, in5243_2;
    wire c5243;
    assign in5243_1 = {pp33[29]};
    assign in5243_2 = {pp34[28]};
    Full_Adder FA_5243(s5243, c5243, in5243_1, in5243_2, pp32[30]);
    wire[0:0] s5244, in5244_1, in5244_2;
    wire c5244;
    assign in5244_1 = {pp36[26]};
    assign in5244_2 = {pp37[25]};
    Full_Adder FA_5244(s5244, c5244, in5244_1, in5244_2, pp35[27]);
    wire[0:0] s5245, in5245_1, in5245_2;
    wire c5245;
    assign in5245_1 = {pp39[23]};
    assign in5245_2 = {pp40[22]};
    Full_Adder FA_5245(s5245, c5245, in5245_1, in5245_2, pp38[24]);
    wire[0:0] s5246, in5246_1, in5246_2;
    wire c5246;
    assign in5246_1 = {pp42[20]};
    assign in5246_2 = {pp43[19]};
    Full_Adder FA_5246(s5246, c5246, in5246_1, in5246_2, pp41[21]);
    wire[0:0] s5247, in5247_1, in5247_2;
    wire c5247;
    assign in5247_1 = {pp45[17]};
    assign in5247_2 = {pp46[16]};
    Full_Adder FA_5247(s5247, c5247, in5247_1, in5247_2, pp44[18]);
    wire[0:0] s5248, in5248_1, in5248_2;
    wire c5248;
    assign in5248_1 = {pp48[14]};
    assign in5248_2 = {pp49[13]};
    Full_Adder FA_5248(s5248, c5248, in5248_1, in5248_2, pp47[15]);
    wire[0:0] s5249, in5249_1, in5249_2;
    wire c5249;
    assign in5249_1 = {pp51[11]};
    assign in5249_2 = {pp52[10]};
    Full_Adder FA_5249(s5249, c5249, in5249_1, in5249_2, pp50[12]);
    wire[0:0] s5250, in5250_1, in5250_2;
    wire c5250;
    assign in5250_1 = {pp54[8]};
    assign in5250_2 = {pp55[7]};
    Full_Adder FA_5250(s5250, c5250, in5250_1, in5250_2, pp53[9]);
    wire[0:0] s5251, in5251_1, in5251_2;
    wire c5251;
    assign in5251_1 = {pp57[5]};
    assign in5251_2 = {pp58[4]};
    Full_Adder FA_5251(s5251, c5251, in5251_1, in5251_2, pp56[6]);
    wire[0:0] s5252, in5252_1, in5252_2;
    wire c5252;
    assign in5252_1 = {pp60[2]};
    assign in5252_2 = {pp61[1]};
    Full_Adder FA_5252(s5252, c5252, in5252_1, in5252_2, pp59[3]);
    wire[0:0] s5253, in5253_1, in5253_2;
    wire c5253;
    assign in5253_1 = {c1813};
    assign in5253_2 = {c1814};
    Full_Adder FA_5253(s5253, c5253, in5253_1, in5253_2, pp62[0]);
    wire[0:0] s5254, in5254_1, in5254_2;
    wire c5254;
    assign in5254_1 = {c1816};
    assign in5254_2 = {s1817[0]};
    Full_Adder FA_5254(s5254, c5254, in5254_1, in5254_2, c1815);
    wire[0:0] s5255, in5255_1, in5255_2;
    wire c5255;
    assign in5255_1 = {s1819[0]};
    assign in5255_2 = {s1820[0]};
    Full_Adder FA_5255(s5255, c5255, in5255_1, in5255_2, s1818[0]);
    wire[0:0] s5256, in5256_1, in5256_2;
    wire c5256;
    assign in5256_1 = {pp18[45]};
    assign in5256_2 = {pp19[44]};
    Full_Adder FA_5256(s5256, c5256, in5256_1, in5256_2, pp17[46]);
    wire[0:0] s5257, in5257_1, in5257_2;
    wire c5257;
    assign in5257_1 = {pp21[42]};
    assign in5257_2 = {pp22[41]};
    Full_Adder FA_5257(s5257, c5257, in5257_1, in5257_2, pp20[43]);
    wire[0:0] s5258, in5258_1, in5258_2;
    wire c5258;
    assign in5258_1 = {pp24[39]};
    assign in5258_2 = {pp25[38]};
    Full_Adder FA_5258(s5258, c5258, in5258_1, in5258_2, pp23[40]);
    wire[0:0] s5259, in5259_1, in5259_2;
    wire c5259;
    assign in5259_1 = {pp27[36]};
    assign in5259_2 = {pp28[35]};
    Full_Adder FA_5259(s5259, c5259, in5259_1, in5259_2, pp26[37]);
    wire[0:0] s5260, in5260_1, in5260_2;
    wire c5260;
    assign in5260_1 = {pp30[33]};
    assign in5260_2 = {pp31[32]};
    Full_Adder FA_5260(s5260, c5260, in5260_1, in5260_2, pp29[34]);
    wire[0:0] s5261, in5261_1, in5261_2;
    wire c5261;
    assign in5261_1 = {pp33[30]};
    assign in5261_2 = {pp34[29]};
    Full_Adder FA_5261(s5261, c5261, in5261_1, in5261_2, pp32[31]);
    wire[0:0] s5262, in5262_1, in5262_2;
    wire c5262;
    assign in5262_1 = {pp36[27]};
    assign in5262_2 = {pp37[26]};
    Full_Adder FA_5262(s5262, c5262, in5262_1, in5262_2, pp35[28]);
    wire[0:0] s5263, in5263_1, in5263_2;
    wire c5263;
    assign in5263_1 = {pp39[24]};
    assign in5263_2 = {pp40[23]};
    Full_Adder FA_5263(s5263, c5263, in5263_1, in5263_2, pp38[25]);
    wire[0:0] s5264, in5264_1, in5264_2;
    wire c5264;
    assign in5264_1 = {pp42[21]};
    assign in5264_2 = {pp43[20]};
    Full_Adder FA_5264(s5264, c5264, in5264_1, in5264_2, pp41[22]);
    wire[0:0] s5265, in5265_1, in5265_2;
    wire c5265;
    assign in5265_1 = {pp45[18]};
    assign in5265_2 = {pp46[17]};
    Full_Adder FA_5265(s5265, c5265, in5265_1, in5265_2, pp44[19]);
    wire[0:0] s5266, in5266_1, in5266_2;
    wire c5266;
    assign in5266_1 = {pp48[15]};
    assign in5266_2 = {pp49[14]};
    Full_Adder FA_5266(s5266, c5266, in5266_1, in5266_2, pp47[16]);
    wire[0:0] s5267, in5267_1, in5267_2;
    wire c5267;
    assign in5267_1 = {pp51[12]};
    assign in5267_2 = {pp52[11]};
    Full_Adder FA_5267(s5267, c5267, in5267_1, in5267_2, pp50[13]);
    wire[0:0] s5268, in5268_1, in5268_2;
    wire c5268;
    assign in5268_1 = {pp54[9]};
    assign in5268_2 = {pp55[8]};
    Full_Adder FA_5268(s5268, c5268, in5268_1, in5268_2, pp53[10]);
    wire[0:0] s5269, in5269_1, in5269_2;
    wire c5269;
    assign in5269_1 = {pp57[6]};
    assign in5269_2 = {pp58[5]};
    Full_Adder FA_5269(s5269, c5269, in5269_1, in5269_2, pp56[7]);
    wire[0:0] s5270, in5270_1, in5270_2;
    wire c5270;
    assign in5270_1 = {pp60[3]};
    assign in5270_2 = {pp61[2]};
    Full_Adder FA_5270(s5270, c5270, in5270_1, in5270_2, pp59[4]);
    wire[0:0] s5271, in5271_1, in5271_2;
    wire c5271;
    assign in5271_1 = {pp63[0]};
    assign in5271_2 = {c1817};
    Full_Adder FA_5271(s5271, c5271, in5271_1, in5271_2, pp62[1]);
    wire[0:0] s5272, in5272_1, in5272_2;
    wire c5272;
    assign in5272_1 = {c1819};
    assign in5272_2 = {c1820};
    Full_Adder FA_5272(s5272, c5272, in5272_1, in5272_2, c1818);
    wire[0:0] s5273, in5273_1, in5273_2;
    wire c5273;
    assign in5273_1 = {s1822[0]};
    assign in5273_2 = {s1823[0]};
    Full_Adder FA_5273(s5273, c5273, in5273_1, in5273_2, c1821);
    wire[0:0] s5274, in5274_1, in5274_2;
    wire c5274;
    assign in5274_1 = {s1825[0]};
    assign in5274_2 = {s1826[0]};
    Full_Adder FA_5274(s5274, c5274, in5274_1, in5274_2, s1824[0]);
    wire[0:0] s5275, in5275_1, in5275_2;
    wire c5275;
    assign in5275_1 = {pp21[43]};
    assign in5275_2 = {pp22[42]};
    Full_Adder FA_5275(s5275, c5275, in5275_1, in5275_2, pp20[44]);
    wire[0:0] s5276, in5276_1, in5276_2;
    wire c5276;
    assign in5276_1 = {pp24[40]};
    assign in5276_2 = {pp25[39]};
    Full_Adder FA_5276(s5276, c5276, in5276_1, in5276_2, pp23[41]);
    wire[0:0] s5277, in5277_1, in5277_2;
    wire c5277;
    assign in5277_1 = {pp27[37]};
    assign in5277_2 = {pp28[36]};
    Full_Adder FA_5277(s5277, c5277, in5277_1, in5277_2, pp26[38]);
    wire[0:0] s5278, in5278_1, in5278_2;
    wire c5278;
    assign in5278_1 = {pp30[34]};
    assign in5278_2 = {pp31[33]};
    Full_Adder FA_5278(s5278, c5278, in5278_1, in5278_2, pp29[35]);
    wire[0:0] s5279, in5279_1, in5279_2;
    wire c5279;
    assign in5279_1 = {pp33[31]};
    assign in5279_2 = {pp34[30]};
    Full_Adder FA_5279(s5279, c5279, in5279_1, in5279_2, pp32[32]);
    wire[0:0] s5280, in5280_1, in5280_2;
    wire c5280;
    assign in5280_1 = {pp36[28]};
    assign in5280_2 = {pp37[27]};
    Full_Adder FA_5280(s5280, c5280, in5280_1, in5280_2, pp35[29]);
    wire[0:0] s5281, in5281_1, in5281_2;
    wire c5281;
    assign in5281_1 = {pp39[25]};
    assign in5281_2 = {pp40[24]};
    Full_Adder FA_5281(s5281, c5281, in5281_1, in5281_2, pp38[26]);
    wire[0:0] s5282, in5282_1, in5282_2;
    wire c5282;
    assign in5282_1 = {pp42[22]};
    assign in5282_2 = {pp43[21]};
    Full_Adder FA_5282(s5282, c5282, in5282_1, in5282_2, pp41[23]);
    wire[0:0] s5283, in5283_1, in5283_2;
    wire c5283;
    assign in5283_1 = {pp45[19]};
    assign in5283_2 = {pp46[18]};
    Full_Adder FA_5283(s5283, c5283, in5283_1, in5283_2, pp44[20]);
    wire[0:0] s5284, in5284_1, in5284_2;
    wire c5284;
    assign in5284_1 = {pp48[16]};
    assign in5284_2 = {pp49[15]};
    Full_Adder FA_5284(s5284, c5284, in5284_1, in5284_2, pp47[17]);
    wire[0:0] s5285, in5285_1, in5285_2;
    wire c5285;
    assign in5285_1 = {pp51[13]};
    assign in5285_2 = {pp52[12]};
    Full_Adder FA_5285(s5285, c5285, in5285_1, in5285_2, pp50[14]);
    wire[0:0] s5286, in5286_1, in5286_2;
    wire c5286;
    assign in5286_1 = {pp54[10]};
    assign in5286_2 = {pp55[9]};
    Full_Adder FA_5286(s5286, c5286, in5286_1, in5286_2, pp53[11]);
    wire[0:0] s5287, in5287_1, in5287_2;
    wire c5287;
    assign in5287_1 = {pp57[7]};
    assign in5287_2 = {pp58[6]};
    Full_Adder FA_5287(s5287, c5287, in5287_1, in5287_2, pp56[8]);
    wire[0:0] s5288, in5288_1, in5288_2;
    wire c5288;
    assign in5288_1 = {pp60[4]};
    assign in5288_2 = {pp61[3]};
    Full_Adder FA_5288(s5288, c5288, in5288_1, in5288_2, pp59[5]);
    wire[0:0] s5289, in5289_1, in5289_2;
    wire c5289;
    assign in5289_1 = {pp63[1]};
    assign in5289_2 = {pp64[0]};
    Full_Adder FA_5289(s5289, c5289, in5289_1, in5289_2, pp62[2]);
    wire[0:0] s5290, in5290_1, in5290_2;
    wire c5290;
    assign in5290_1 = {c1823};
    assign in5290_2 = {c1824};
    Full_Adder FA_5290(s5290, c5290, in5290_1, in5290_2, c1822);
    wire[0:0] s5291, in5291_1, in5291_2;
    wire c5291;
    assign in5291_1 = {c1826};
    assign in5291_2 = {c1827};
    Full_Adder FA_5291(s5291, c5291, in5291_1, in5291_2, c1825);
    wire[0:0] s5292, in5292_1, in5292_2;
    wire c5292;
    assign in5292_1 = {s1829[0]};
    assign in5292_2 = {s1830[0]};
    Full_Adder FA_5292(s5292, c5292, in5292_1, in5292_2, s1828[0]);
    wire[0:0] s5293, in5293_1, in5293_2;
    wire c5293;
    assign in5293_1 = {s1832[0]};
    assign in5293_2 = {s1833[0]};
    Full_Adder FA_5293(s5293, c5293, in5293_1, in5293_2, s1831[0]);
    wire[0:0] s5294, in5294_1, in5294_2;
    wire c5294;
    assign in5294_1 = {pp24[41]};
    assign in5294_2 = {pp25[40]};
    Full_Adder FA_5294(s5294, c5294, in5294_1, in5294_2, pp23[42]);
    wire[0:0] s5295, in5295_1, in5295_2;
    wire c5295;
    assign in5295_1 = {pp27[38]};
    assign in5295_2 = {pp28[37]};
    Full_Adder FA_5295(s5295, c5295, in5295_1, in5295_2, pp26[39]);
    wire[0:0] s5296, in5296_1, in5296_2;
    wire c5296;
    assign in5296_1 = {pp30[35]};
    assign in5296_2 = {pp31[34]};
    Full_Adder FA_5296(s5296, c5296, in5296_1, in5296_2, pp29[36]);
    wire[0:0] s5297, in5297_1, in5297_2;
    wire c5297;
    assign in5297_1 = {pp33[32]};
    assign in5297_2 = {pp34[31]};
    Full_Adder FA_5297(s5297, c5297, in5297_1, in5297_2, pp32[33]);
    wire[0:0] s5298, in5298_1, in5298_2;
    wire c5298;
    assign in5298_1 = {pp36[29]};
    assign in5298_2 = {pp37[28]};
    Full_Adder FA_5298(s5298, c5298, in5298_1, in5298_2, pp35[30]);
    wire[0:0] s5299, in5299_1, in5299_2;
    wire c5299;
    assign in5299_1 = {pp39[26]};
    assign in5299_2 = {pp40[25]};
    Full_Adder FA_5299(s5299, c5299, in5299_1, in5299_2, pp38[27]);
    wire[0:0] s5300, in5300_1, in5300_2;
    wire c5300;
    assign in5300_1 = {pp42[23]};
    assign in5300_2 = {pp43[22]};
    Full_Adder FA_5300(s5300, c5300, in5300_1, in5300_2, pp41[24]);
    wire[0:0] s5301, in5301_1, in5301_2;
    wire c5301;
    assign in5301_1 = {pp45[20]};
    assign in5301_2 = {pp46[19]};
    Full_Adder FA_5301(s5301, c5301, in5301_1, in5301_2, pp44[21]);
    wire[0:0] s5302, in5302_1, in5302_2;
    wire c5302;
    assign in5302_1 = {pp48[17]};
    assign in5302_2 = {pp49[16]};
    Full_Adder FA_5302(s5302, c5302, in5302_1, in5302_2, pp47[18]);
    wire[0:0] s5303, in5303_1, in5303_2;
    wire c5303;
    assign in5303_1 = {pp51[14]};
    assign in5303_2 = {pp52[13]};
    Full_Adder FA_5303(s5303, c5303, in5303_1, in5303_2, pp50[15]);
    wire[0:0] s5304, in5304_1, in5304_2;
    wire c5304;
    assign in5304_1 = {pp54[11]};
    assign in5304_2 = {pp55[10]};
    Full_Adder FA_5304(s5304, c5304, in5304_1, in5304_2, pp53[12]);
    wire[0:0] s5305, in5305_1, in5305_2;
    wire c5305;
    assign in5305_1 = {pp57[8]};
    assign in5305_2 = {pp58[7]};
    Full_Adder FA_5305(s5305, c5305, in5305_1, in5305_2, pp56[9]);
    wire[0:0] s5306, in5306_1, in5306_2;
    wire c5306;
    assign in5306_1 = {pp60[5]};
    assign in5306_2 = {pp61[4]};
    Full_Adder FA_5306(s5306, c5306, in5306_1, in5306_2, pp59[6]);
    wire[0:0] s5307, in5307_1, in5307_2;
    wire c5307;
    assign in5307_1 = {pp63[2]};
    assign in5307_2 = {pp64[1]};
    Full_Adder FA_5307(s5307, c5307, in5307_1, in5307_2, pp62[3]);
    wire[0:0] s5308, in5308_1, in5308_2;
    wire c5308;
    assign in5308_1 = {c1828};
    assign in5308_2 = {c1829};
    Full_Adder FA_5308(s5308, c5308, in5308_1, in5308_2, pp65[0]);
    wire[0:0] s5309, in5309_1, in5309_2;
    wire c5309;
    assign in5309_1 = {c1831};
    assign in5309_2 = {c1832};
    Full_Adder FA_5309(s5309, c5309, in5309_1, in5309_2, c1830);
    wire[0:0] s5310, in5310_1, in5310_2;
    wire c5310;
    assign in5310_1 = {c1834};
    assign in5310_2 = {s1835[0]};
    Full_Adder FA_5310(s5310, c5310, in5310_1, in5310_2, c1833);
    wire[0:0] s5311, in5311_1, in5311_2;
    wire c5311;
    assign in5311_1 = {s1837[0]};
    assign in5311_2 = {s1838[0]};
    Full_Adder FA_5311(s5311, c5311, in5311_1, in5311_2, s1836[0]);
    wire[0:0] s5312, in5312_1, in5312_2;
    wire c5312;
    assign in5312_1 = {s1840[0]};
    assign in5312_2 = {s1841[0]};
    Full_Adder FA_5312(s5312, c5312, in5312_1, in5312_2, s1839[0]);
    wire[0:0] s5313, in5313_1, in5313_2;
    wire c5313;
    assign in5313_1 = {pp27[39]};
    assign in5313_2 = {pp28[38]};
    Full_Adder FA_5313(s5313, c5313, in5313_1, in5313_2, pp26[40]);
    wire[0:0] s5314, in5314_1, in5314_2;
    wire c5314;
    assign in5314_1 = {pp30[36]};
    assign in5314_2 = {pp31[35]};
    Full_Adder FA_5314(s5314, c5314, in5314_1, in5314_2, pp29[37]);
    wire[0:0] s5315, in5315_1, in5315_2;
    wire c5315;
    assign in5315_1 = {pp33[33]};
    assign in5315_2 = {pp34[32]};
    Full_Adder FA_5315(s5315, c5315, in5315_1, in5315_2, pp32[34]);
    wire[0:0] s5316, in5316_1, in5316_2;
    wire c5316;
    assign in5316_1 = {pp36[30]};
    assign in5316_2 = {pp37[29]};
    Full_Adder FA_5316(s5316, c5316, in5316_1, in5316_2, pp35[31]);
    wire[0:0] s5317, in5317_1, in5317_2;
    wire c5317;
    assign in5317_1 = {pp39[27]};
    assign in5317_2 = {pp40[26]};
    Full_Adder FA_5317(s5317, c5317, in5317_1, in5317_2, pp38[28]);
    wire[0:0] s5318, in5318_1, in5318_2;
    wire c5318;
    assign in5318_1 = {pp42[24]};
    assign in5318_2 = {pp43[23]};
    Full_Adder FA_5318(s5318, c5318, in5318_1, in5318_2, pp41[25]);
    wire[0:0] s5319, in5319_1, in5319_2;
    wire c5319;
    assign in5319_1 = {pp45[21]};
    assign in5319_2 = {pp46[20]};
    Full_Adder FA_5319(s5319, c5319, in5319_1, in5319_2, pp44[22]);
    wire[0:0] s5320, in5320_1, in5320_2;
    wire c5320;
    assign in5320_1 = {pp48[18]};
    assign in5320_2 = {pp49[17]};
    Full_Adder FA_5320(s5320, c5320, in5320_1, in5320_2, pp47[19]);
    wire[0:0] s5321, in5321_1, in5321_2;
    wire c5321;
    assign in5321_1 = {pp51[15]};
    assign in5321_2 = {pp52[14]};
    Full_Adder FA_5321(s5321, c5321, in5321_1, in5321_2, pp50[16]);
    wire[0:0] s5322, in5322_1, in5322_2;
    wire c5322;
    assign in5322_1 = {pp54[12]};
    assign in5322_2 = {pp55[11]};
    Full_Adder FA_5322(s5322, c5322, in5322_1, in5322_2, pp53[13]);
    wire[0:0] s5323, in5323_1, in5323_2;
    wire c5323;
    assign in5323_1 = {pp57[9]};
    assign in5323_2 = {pp58[8]};
    Full_Adder FA_5323(s5323, c5323, in5323_1, in5323_2, pp56[10]);
    wire[0:0] s5324, in5324_1, in5324_2;
    wire c5324;
    assign in5324_1 = {pp60[6]};
    assign in5324_2 = {pp61[5]};
    Full_Adder FA_5324(s5324, c5324, in5324_1, in5324_2, pp59[7]);
    wire[0:0] s5325, in5325_1, in5325_2;
    wire c5325;
    assign in5325_1 = {pp63[3]};
    assign in5325_2 = {pp64[2]};
    Full_Adder FA_5325(s5325, c5325, in5325_1, in5325_2, pp62[4]);
    wire[0:0] s5326, in5326_1, in5326_2;
    wire c5326;
    assign in5326_1 = {pp66[0]};
    assign in5326_2 = {c1835};
    Full_Adder FA_5326(s5326, c5326, in5326_1, in5326_2, pp65[1]);
    wire[0:0] s5327, in5327_1, in5327_2;
    wire c5327;
    assign in5327_1 = {c1837};
    assign in5327_2 = {c1838};
    Full_Adder FA_5327(s5327, c5327, in5327_1, in5327_2, c1836);
    wire[0:0] s5328, in5328_1, in5328_2;
    wire c5328;
    assign in5328_1 = {c1840};
    assign in5328_2 = {c1841};
    Full_Adder FA_5328(s5328, c5328, in5328_1, in5328_2, c1839);
    wire[0:0] s5329, in5329_1, in5329_2;
    wire c5329;
    assign in5329_1 = {s1843[0]};
    assign in5329_2 = {s1844[0]};
    Full_Adder FA_5329(s5329, c5329, in5329_1, in5329_2, c1842);
    wire[0:0] s5330, in5330_1, in5330_2;
    wire c5330;
    assign in5330_1 = {s1846[0]};
    assign in5330_2 = {s1847[0]};
    Full_Adder FA_5330(s5330, c5330, in5330_1, in5330_2, s1845[0]);
    wire[0:0] s5331, in5331_1, in5331_2;
    wire c5331;
    assign in5331_1 = {s1849[0]};
    assign in5331_2 = {s1850[0]};
    Full_Adder FA_5331(s5331, c5331, in5331_1, in5331_2, s1848[0]);
    wire[0:0] s5332, in5332_1, in5332_2;
    wire c5332;
    assign in5332_1 = {pp30[37]};
    assign in5332_2 = {pp31[36]};
    Full_Adder FA_5332(s5332, c5332, in5332_1, in5332_2, pp29[38]);
    wire[0:0] s5333, in5333_1, in5333_2;
    wire c5333;
    assign in5333_1 = {pp33[34]};
    assign in5333_2 = {pp34[33]};
    Full_Adder FA_5333(s5333, c5333, in5333_1, in5333_2, pp32[35]);
    wire[0:0] s5334, in5334_1, in5334_2;
    wire c5334;
    assign in5334_1 = {pp36[31]};
    assign in5334_2 = {pp37[30]};
    Full_Adder FA_5334(s5334, c5334, in5334_1, in5334_2, pp35[32]);
    wire[0:0] s5335, in5335_1, in5335_2;
    wire c5335;
    assign in5335_1 = {pp39[28]};
    assign in5335_2 = {pp40[27]};
    Full_Adder FA_5335(s5335, c5335, in5335_1, in5335_2, pp38[29]);
    wire[0:0] s5336, in5336_1, in5336_2;
    wire c5336;
    assign in5336_1 = {pp42[25]};
    assign in5336_2 = {pp43[24]};
    Full_Adder FA_5336(s5336, c5336, in5336_1, in5336_2, pp41[26]);
    wire[0:0] s5337, in5337_1, in5337_2;
    wire c5337;
    assign in5337_1 = {pp45[22]};
    assign in5337_2 = {pp46[21]};
    Full_Adder FA_5337(s5337, c5337, in5337_1, in5337_2, pp44[23]);
    wire[0:0] s5338, in5338_1, in5338_2;
    wire c5338;
    assign in5338_1 = {pp48[19]};
    assign in5338_2 = {pp49[18]};
    Full_Adder FA_5338(s5338, c5338, in5338_1, in5338_2, pp47[20]);
    wire[0:0] s5339, in5339_1, in5339_2;
    wire c5339;
    assign in5339_1 = {pp51[16]};
    assign in5339_2 = {pp52[15]};
    Full_Adder FA_5339(s5339, c5339, in5339_1, in5339_2, pp50[17]);
    wire[0:0] s5340, in5340_1, in5340_2;
    wire c5340;
    assign in5340_1 = {pp54[13]};
    assign in5340_2 = {pp55[12]};
    Full_Adder FA_5340(s5340, c5340, in5340_1, in5340_2, pp53[14]);
    wire[0:0] s5341, in5341_1, in5341_2;
    wire c5341;
    assign in5341_1 = {pp57[10]};
    assign in5341_2 = {pp58[9]};
    Full_Adder FA_5341(s5341, c5341, in5341_1, in5341_2, pp56[11]);
    wire[0:0] s5342, in5342_1, in5342_2;
    wire c5342;
    assign in5342_1 = {pp60[7]};
    assign in5342_2 = {pp61[6]};
    Full_Adder FA_5342(s5342, c5342, in5342_1, in5342_2, pp59[8]);
    wire[0:0] s5343, in5343_1, in5343_2;
    wire c5343;
    assign in5343_1 = {pp63[4]};
    assign in5343_2 = {pp64[3]};
    Full_Adder FA_5343(s5343, c5343, in5343_1, in5343_2, pp62[5]);
    wire[0:0] s5344, in5344_1, in5344_2;
    wire c5344;
    assign in5344_1 = {pp66[1]};
    assign in5344_2 = {pp67[0]};
    Full_Adder FA_5344(s5344, c5344, in5344_1, in5344_2, pp65[2]);
    wire[0:0] s5345, in5345_1, in5345_2;
    wire c5345;
    assign in5345_1 = {c1844};
    assign in5345_2 = {c1845};
    Full_Adder FA_5345(s5345, c5345, in5345_1, in5345_2, c1843);
    wire[0:0] s5346, in5346_1, in5346_2;
    wire c5346;
    assign in5346_1 = {c1847};
    assign in5346_2 = {c1848};
    Full_Adder FA_5346(s5346, c5346, in5346_1, in5346_2, c1846);
    wire[0:0] s5347, in5347_1, in5347_2;
    wire c5347;
    assign in5347_1 = {c1850};
    assign in5347_2 = {c1851};
    Full_Adder FA_5347(s5347, c5347, in5347_1, in5347_2, c1849);
    wire[0:0] s5348, in5348_1, in5348_2;
    wire c5348;
    assign in5348_1 = {s1853[0]};
    assign in5348_2 = {s1854[0]};
    Full_Adder FA_5348(s5348, c5348, in5348_1, in5348_2, s1852[0]);
    wire[0:0] s5349, in5349_1, in5349_2;
    wire c5349;
    assign in5349_1 = {s1856[0]};
    assign in5349_2 = {s1857[0]};
    Full_Adder FA_5349(s5349, c5349, in5349_1, in5349_2, s1855[0]);
    wire[0:0] s5350, in5350_1, in5350_2;
    wire c5350;
    assign in5350_1 = {s1859[0]};
    assign in5350_2 = {s1860[0]};
    Full_Adder FA_5350(s5350, c5350, in5350_1, in5350_2, s1858[0]);
    wire[0:0] s5351, in5351_1, in5351_2;
    wire c5351;
    assign in5351_1 = {pp33[35]};
    assign in5351_2 = {pp34[34]};
    Full_Adder FA_5351(s5351, c5351, in5351_1, in5351_2, pp32[36]);
    wire[0:0] s5352, in5352_1, in5352_2;
    wire c5352;
    assign in5352_1 = {pp36[32]};
    assign in5352_2 = {pp37[31]};
    Full_Adder FA_5352(s5352, c5352, in5352_1, in5352_2, pp35[33]);
    wire[0:0] s5353, in5353_1, in5353_2;
    wire c5353;
    assign in5353_1 = {pp39[29]};
    assign in5353_2 = {pp40[28]};
    Full_Adder FA_5353(s5353, c5353, in5353_1, in5353_2, pp38[30]);
    wire[0:0] s5354, in5354_1, in5354_2;
    wire c5354;
    assign in5354_1 = {pp42[26]};
    assign in5354_2 = {pp43[25]};
    Full_Adder FA_5354(s5354, c5354, in5354_1, in5354_2, pp41[27]);
    wire[0:0] s5355, in5355_1, in5355_2;
    wire c5355;
    assign in5355_1 = {pp45[23]};
    assign in5355_2 = {pp46[22]};
    Full_Adder FA_5355(s5355, c5355, in5355_1, in5355_2, pp44[24]);
    wire[0:0] s5356, in5356_1, in5356_2;
    wire c5356;
    assign in5356_1 = {pp48[20]};
    assign in5356_2 = {pp49[19]};
    Full_Adder FA_5356(s5356, c5356, in5356_1, in5356_2, pp47[21]);
    wire[0:0] s5357, in5357_1, in5357_2;
    wire c5357;
    assign in5357_1 = {pp51[17]};
    assign in5357_2 = {pp52[16]};
    Full_Adder FA_5357(s5357, c5357, in5357_1, in5357_2, pp50[18]);
    wire[0:0] s5358, in5358_1, in5358_2;
    wire c5358;
    assign in5358_1 = {pp54[14]};
    assign in5358_2 = {pp55[13]};
    Full_Adder FA_5358(s5358, c5358, in5358_1, in5358_2, pp53[15]);
    wire[0:0] s5359, in5359_1, in5359_2;
    wire c5359;
    assign in5359_1 = {pp57[11]};
    assign in5359_2 = {pp58[10]};
    Full_Adder FA_5359(s5359, c5359, in5359_1, in5359_2, pp56[12]);
    wire[0:0] s5360, in5360_1, in5360_2;
    wire c5360;
    assign in5360_1 = {pp60[8]};
    assign in5360_2 = {pp61[7]};
    Full_Adder FA_5360(s5360, c5360, in5360_1, in5360_2, pp59[9]);
    wire[0:0] s5361, in5361_1, in5361_2;
    wire c5361;
    assign in5361_1 = {pp63[5]};
    assign in5361_2 = {pp64[4]};
    Full_Adder FA_5361(s5361, c5361, in5361_1, in5361_2, pp62[6]);
    wire[0:0] s5362, in5362_1, in5362_2;
    wire c5362;
    assign in5362_1 = {pp66[2]};
    assign in5362_2 = {pp67[1]};
    Full_Adder FA_5362(s5362, c5362, in5362_1, in5362_2, pp65[3]);
    wire[0:0] s5363, in5363_1, in5363_2;
    wire c5363;
    assign in5363_1 = {c1852};
    assign in5363_2 = {c1853};
    Full_Adder FA_5363(s5363, c5363, in5363_1, in5363_2, pp68[0]);
    wire[0:0] s5364, in5364_1, in5364_2;
    wire c5364;
    assign in5364_1 = {c1855};
    assign in5364_2 = {c1856};
    Full_Adder FA_5364(s5364, c5364, in5364_1, in5364_2, c1854);
    wire[0:0] s5365, in5365_1, in5365_2;
    wire c5365;
    assign in5365_1 = {c1858};
    assign in5365_2 = {c1859};
    Full_Adder FA_5365(s5365, c5365, in5365_1, in5365_2, c1857);
    wire[0:0] s5366, in5366_1, in5366_2;
    wire c5366;
    assign in5366_1 = {c1861};
    assign in5366_2 = {s1862[0]};
    Full_Adder FA_5366(s5366, c5366, in5366_1, in5366_2, c1860);
    wire[0:0] s5367, in5367_1, in5367_2;
    wire c5367;
    assign in5367_1 = {s1864[0]};
    assign in5367_2 = {s1865[0]};
    Full_Adder FA_5367(s5367, c5367, in5367_1, in5367_2, s1863[0]);
    wire[0:0] s5368, in5368_1, in5368_2;
    wire c5368;
    assign in5368_1 = {s1867[0]};
    assign in5368_2 = {s1868[0]};
    Full_Adder FA_5368(s5368, c5368, in5368_1, in5368_2, s1866[0]);
    wire[0:0] s5369, in5369_1, in5369_2;
    wire c5369;
    assign in5369_1 = {s1870[0]};
    assign in5369_2 = {s1871[0]};
    Full_Adder FA_5369(s5369, c5369, in5369_1, in5369_2, s1869[0]);
    wire[0:0] s5370, in5370_1, in5370_2;
    wire c5370;
    assign in5370_1 = {pp36[33]};
    assign in5370_2 = {pp37[32]};
    Full_Adder FA_5370(s5370, c5370, in5370_1, in5370_2, pp35[34]);
    wire[0:0] s5371, in5371_1, in5371_2;
    wire c5371;
    assign in5371_1 = {pp39[30]};
    assign in5371_2 = {pp40[29]};
    Full_Adder FA_5371(s5371, c5371, in5371_1, in5371_2, pp38[31]);
    wire[0:0] s5372, in5372_1, in5372_2;
    wire c5372;
    assign in5372_1 = {pp42[27]};
    assign in5372_2 = {pp43[26]};
    Full_Adder FA_5372(s5372, c5372, in5372_1, in5372_2, pp41[28]);
    wire[0:0] s5373, in5373_1, in5373_2;
    wire c5373;
    assign in5373_1 = {pp45[24]};
    assign in5373_2 = {pp46[23]};
    Full_Adder FA_5373(s5373, c5373, in5373_1, in5373_2, pp44[25]);
    wire[0:0] s5374, in5374_1, in5374_2;
    wire c5374;
    assign in5374_1 = {pp48[21]};
    assign in5374_2 = {pp49[20]};
    Full_Adder FA_5374(s5374, c5374, in5374_1, in5374_2, pp47[22]);
    wire[0:0] s5375, in5375_1, in5375_2;
    wire c5375;
    assign in5375_1 = {pp51[18]};
    assign in5375_2 = {pp52[17]};
    Full_Adder FA_5375(s5375, c5375, in5375_1, in5375_2, pp50[19]);
    wire[0:0] s5376, in5376_1, in5376_2;
    wire c5376;
    assign in5376_1 = {pp54[15]};
    assign in5376_2 = {pp55[14]};
    Full_Adder FA_5376(s5376, c5376, in5376_1, in5376_2, pp53[16]);
    wire[0:0] s5377, in5377_1, in5377_2;
    wire c5377;
    assign in5377_1 = {pp57[12]};
    assign in5377_2 = {pp58[11]};
    Full_Adder FA_5377(s5377, c5377, in5377_1, in5377_2, pp56[13]);
    wire[0:0] s5378, in5378_1, in5378_2;
    wire c5378;
    assign in5378_1 = {pp60[9]};
    assign in5378_2 = {pp61[8]};
    Full_Adder FA_5378(s5378, c5378, in5378_1, in5378_2, pp59[10]);
    wire[0:0] s5379, in5379_1, in5379_2;
    wire c5379;
    assign in5379_1 = {pp63[6]};
    assign in5379_2 = {pp64[5]};
    Full_Adder FA_5379(s5379, c5379, in5379_1, in5379_2, pp62[7]);
    wire[0:0] s5380, in5380_1, in5380_2;
    wire c5380;
    assign in5380_1 = {pp66[3]};
    assign in5380_2 = {pp67[2]};
    Full_Adder FA_5380(s5380, c5380, in5380_1, in5380_2, pp65[4]);
    wire[0:0] s5381, in5381_1, in5381_2;
    wire c5381;
    assign in5381_1 = {pp69[0]};
    assign in5381_2 = {c1862};
    Full_Adder FA_5381(s5381, c5381, in5381_1, in5381_2, pp68[1]);
    wire[0:0] s5382, in5382_1, in5382_2;
    wire c5382;
    assign in5382_1 = {c1864};
    assign in5382_2 = {c1865};
    Full_Adder FA_5382(s5382, c5382, in5382_1, in5382_2, c1863);
    wire[0:0] s5383, in5383_1, in5383_2;
    wire c5383;
    assign in5383_1 = {c1867};
    assign in5383_2 = {c1868};
    Full_Adder FA_5383(s5383, c5383, in5383_1, in5383_2, c1866);
    wire[0:0] s5384, in5384_1, in5384_2;
    wire c5384;
    assign in5384_1 = {c1870};
    assign in5384_2 = {c1871};
    Full_Adder FA_5384(s5384, c5384, in5384_1, in5384_2, c1869);
    wire[0:0] s5385, in5385_1, in5385_2;
    wire c5385;
    assign in5385_1 = {s1873[0]};
    assign in5385_2 = {s1874[0]};
    Full_Adder FA_5385(s5385, c5385, in5385_1, in5385_2, c1872);
    wire[0:0] s5386, in5386_1, in5386_2;
    wire c5386;
    assign in5386_1 = {s1876[0]};
    assign in5386_2 = {s1877[0]};
    Full_Adder FA_5386(s5386, c5386, in5386_1, in5386_2, s1875[0]);
    wire[0:0] s5387, in5387_1, in5387_2;
    wire c5387;
    assign in5387_1 = {s1879[0]};
    assign in5387_2 = {s1880[0]};
    Full_Adder FA_5387(s5387, c5387, in5387_1, in5387_2, s1878[0]);
    wire[0:0] s5388, in5388_1, in5388_2;
    wire c5388;
    assign in5388_1 = {s1882[0]};
    assign in5388_2 = {s1883[0]};
    Full_Adder FA_5388(s5388, c5388, in5388_1, in5388_2, s1881[0]);
    wire[0:0] s5389, in5389_1, in5389_2;
    wire c5389;
    assign in5389_1 = {pp39[31]};
    assign in5389_2 = {pp40[30]};
    Full_Adder FA_5389(s5389, c5389, in5389_1, in5389_2, pp38[32]);
    wire[0:0] s5390, in5390_1, in5390_2;
    wire c5390;
    assign in5390_1 = {pp42[28]};
    assign in5390_2 = {pp43[27]};
    Full_Adder FA_5390(s5390, c5390, in5390_1, in5390_2, pp41[29]);
    wire[0:0] s5391, in5391_1, in5391_2;
    wire c5391;
    assign in5391_1 = {pp45[25]};
    assign in5391_2 = {pp46[24]};
    Full_Adder FA_5391(s5391, c5391, in5391_1, in5391_2, pp44[26]);
    wire[0:0] s5392, in5392_1, in5392_2;
    wire c5392;
    assign in5392_1 = {pp48[22]};
    assign in5392_2 = {pp49[21]};
    Full_Adder FA_5392(s5392, c5392, in5392_1, in5392_2, pp47[23]);
    wire[0:0] s5393, in5393_1, in5393_2;
    wire c5393;
    assign in5393_1 = {pp51[19]};
    assign in5393_2 = {pp52[18]};
    Full_Adder FA_5393(s5393, c5393, in5393_1, in5393_2, pp50[20]);
    wire[0:0] s5394, in5394_1, in5394_2;
    wire c5394;
    assign in5394_1 = {pp54[16]};
    assign in5394_2 = {pp55[15]};
    Full_Adder FA_5394(s5394, c5394, in5394_1, in5394_2, pp53[17]);
    wire[0:0] s5395, in5395_1, in5395_2;
    wire c5395;
    assign in5395_1 = {pp57[13]};
    assign in5395_2 = {pp58[12]};
    Full_Adder FA_5395(s5395, c5395, in5395_1, in5395_2, pp56[14]);
    wire[0:0] s5396, in5396_1, in5396_2;
    wire c5396;
    assign in5396_1 = {pp60[10]};
    assign in5396_2 = {pp61[9]};
    Full_Adder FA_5396(s5396, c5396, in5396_1, in5396_2, pp59[11]);
    wire[0:0] s5397, in5397_1, in5397_2;
    wire c5397;
    assign in5397_1 = {pp63[7]};
    assign in5397_2 = {pp64[6]};
    Full_Adder FA_5397(s5397, c5397, in5397_1, in5397_2, pp62[8]);
    wire[0:0] s5398, in5398_1, in5398_2;
    wire c5398;
    assign in5398_1 = {pp66[4]};
    assign in5398_2 = {pp67[3]};
    Full_Adder FA_5398(s5398, c5398, in5398_1, in5398_2, pp65[5]);
    wire[0:0] s5399, in5399_1, in5399_2;
    wire c5399;
    assign in5399_1 = {pp69[1]};
    assign in5399_2 = {pp70[0]};
    Full_Adder FA_5399(s5399, c5399, in5399_1, in5399_2, pp68[2]);
    wire[0:0] s5400, in5400_1, in5400_2;
    wire c5400;
    assign in5400_1 = {c1874};
    assign in5400_2 = {c1875};
    Full_Adder FA_5400(s5400, c5400, in5400_1, in5400_2, c1873);
    wire[0:0] s5401, in5401_1, in5401_2;
    wire c5401;
    assign in5401_1 = {c1877};
    assign in5401_2 = {c1878};
    Full_Adder FA_5401(s5401, c5401, in5401_1, in5401_2, c1876);
    wire[0:0] s5402, in5402_1, in5402_2;
    wire c5402;
    assign in5402_1 = {c1880};
    assign in5402_2 = {c1881};
    Full_Adder FA_5402(s5402, c5402, in5402_1, in5402_2, c1879);
    wire[0:0] s5403, in5403_1, in5403_2;
    wire c5403;
    assign in5403_1 = {c1883};
    assign in5403_2 = {c1884};
    Full_Adder FA_5403(s5403, c5403, in5403_1, in5403_2, c1882);
    wire[0:0] s5404, in5404_1, in5404_2;
    wire c5404;
    assign in5404_1 = {s1886[0]};
    assign in5404_2 = {s1887[0]};
    Full_Adder FA_5404(s5404, c5404, in5404_1, in5404_2, s1885[0]);
    wire[0:0] s5405, in5405_1, in5405_2;
    wire c5405;
    assign in5405_1 = {s1889[0]};
    assign in5405_2 = {s1890[0]};
    Full_Adder FA_5405(s5405, c5405, in5405_1, in5405_2, s1888[0]);
    wire[0:0] s5406, in5406_1, in5406_2;
    wire c5406;
    assign in5406_1 = {s1892[0]};
    assign in5406_2 = {s1893[0]};
    Full_Adder FA_5406(s5406, c5406, in5406_1, in5406_2, s1891[0]);
    wire[0:0] s5407, in5407_1, in5407_2;
    wire c5407;
    assign in5407_1 = {s1895[0]};
    assign in5407_2 = {s1896[0]};
    Full_Adder FA_5407(s5407, c5407, in5407_1, in5407_2, s1894[0]);
    wire[0:0] s5408, in5408_1, in5408_2;
    wire c5408;
    assign in5408_1 = {pp42[29]};
    assign in5408_2 = {pp43[28]};
    Full_Adder FA_5408(s5408, c5408, in5408_1, in5408_2, pp41[30]);
    wire[0:0] s5409, in5409_1, in5409_2;
    wire c5409;
    assign in5409_1 = {pp45[26]};
    assign in5409_2 = {pp46[25]};
    Full_Adder FA_5409(s5409, c5409, in5409_1, in5409_2, pp44[27]);
    wire[0:0] s5410, in5410_1, in5410_2;
    wire c5410;
    assign in5410_1 = {pp48[23]};
    assign in5410_2 = {pp49[22]};
    Full_Adder FA_5410(s5410, c5410, in5410_1, in5410_2, pp47[24]);
    wire[0:0] s5411, in5411_1, in5411_2;
    wire c5411;
    assign in5411_1 = {pp51[20]};
    assign in5411_2 = {pp52[19]};
    Full_Adder FA_5411(s5411, c5411, in5411_1, in5411_2, pp50[21]);
    wire[0:0] s5412, in5412_1, in5412_2;
    wire c5412;
    assign in5412_1 = {pp54[17]};
    assign in5412_2 = {pp55[16]};
    Full_Adder FA_5412(s5412, c5412, in5412_1, in5412_2, pp53[18]);
    wire[0:0] s5413, in5413_1, in5413_2;
    wire c5413;
    assign in5413_1 = {pp57[14]};
    assign in5413_2 = {pp58[13]};
    Full_Adder FA_5413(s5413, c5413, in5413_1, in5413_2, pp56[15]);
    wire[0:0] s5414, in5414_1, in5414_2;
    wire c5414;
    assign in5414_1 = {pp60[11]};
    assign in5414_2 = {pp61[10]};
    Full_Adder FA_5414(s5414, c5414, in5414_1, in5414_2, pp59[12]);
    wire[0:0] s5415, in5415_1, in5415_2;
    wire c5415;
    assign in5415_1 = {pp63[8]};
    assign in5415_2 = {pp64[7]};
    Full_Adder FA_5415(s5415, c5415, in5415_1, in5415_2, pp62[9]);
    wire[0:0] s5416, in5416_1, in5416_2;
    wire c5416;
    assign in5416_1 = {pp66[5]};
    assign in5416_2 = {pp67[4]};
    Full_Adder FA_5416(s5416, c5416, in5416_1, in5416_2, pp65[6]);
    wire[0:0] s5417, in5417_1, in5417_2;
    wire c5417;
    assign in5417_1 = {pp69[2]};
    assign in5417_2 = {pp70[1]};
    Full_Adder FA_5417(s5417, c5417, in5417_1, in5417_2, pp68[3]);
    wire[0:0] s5418, in5418_1, in5418_2;
    wire c5418;
    assign in5418_1 = {c1885};
    assign in5418_2 = {c1886};
    Full_Adder FA_5418(s5418, c5418, in5418_1, in5418_2, pp71[0]);
    wire[0:0] s5419, in5419_1, in5419_2;
    wire c5419;
    assign in5419_1 = {c1888};
    assign in5419_2 = {c1889};
    Full_Adder FA_5419(s5419, c5419, in5419_1, in5419_2, c1887);
    wire[0:0] s5420, in5420_1, in5420_2;
    wire c5420;
    assign in5420_1 = {c1891};
    assign in5420_2 = {c1892};
    Full_Adder FA_5420(s5420, c5420, in5420_1, in5420_2, c1890);
    wire[0:0] s5421, in5421_1, in5421_2;
    wire c5421;
    assign in5421_1 = {c1894};
    assign in5421_2 = {c1895};
    Full_Adder FA_5421(s5421, c5421, in5421_1, in5421_2, c1893);
    wire[0:0] s5422, in5422_1, in5422_2;
    wire c5422;
    assign in5422_1 = {c1897};
    assign in5422_2 = {s1898[0]};
    Full_Adder FA_5422(s5422, c5422, in5422_1, in5422_2, c1896);
    wire[0:0] s5423, in5423_1, in5423_2;
    wire c5423;
    assign in5423_1 = {s1900[0]};
    assign in5423_2 = {s1901[0]};
    Full_Adder FA_5423(s5423, c5423, in5423_1, in5423_2, s1899[0]);
    wire[0:0] s5424, in5424_1, in5424_2;
    wire c5424;
    assign in5424_1 = {s1903[0]};
    assign in5424_2 = {s1904[0]};
    Full_Adder FA_5424(s5424, c5424, in5424_1, in5424_2, s1902[0]);
    wire[0:0] s5425, in5425_1, in5425_2;
    wire c5425;
    assign in5425_1 = {s1906[0]};
    assign in5425_2 = {s1907[0]};
    Full_Adder FA_5425(s5425, c5425, in5425_1, in5425_2, s1905[0]);
    wire[0:0] s5426, in5426_1, in5426_2;
    wire c5426;
    assign in5426_1 = {s1909[0]};
    assign in5426_2 = {s1910[0]};
    Full_Adder FA_5426(s5426, c5426, in5426_1, in5426_2, s1908[0]);
    wire[0:0] s5427, in5427_1, in5427_2;
    wire c5427;
    assign in5427_1 = {pp45[27]};
    assign in5427_2 = {pp46[26]};
    Full_Adder FA_5427(s5427, c5427, in5427_1, in5427_2, pp44[28]);
    wire[0:0] s5428, in5428_1, in5428_2;
    wire c5428;
    assign in5428_1 = {pp48[24]};
    assign in5428_2 = {pp49[23]};
    Full_Adder FA_5428(s5428, c5428, in5428_1, in5428_2, pp47[25]);
    wire[0:0] s5429, in5429_1, in5429_2;
    wire c5429;
    assign in5429_1 = {pp51[21]};
    assign in5429_2 = {pp52[20]};
    Full_Adder FA_5429(s5429, c5429, in5429_1, in5429_2, pp50[22]);
    wire[0:0] s5430, in5430_1, in5430_2;
    wire c5430;
    assign in5430_1 = {pp54[18]};
    assign in5430_2 = {pp55[17]};
    Full_Adder FA_5430(s5430, c5430, in5430_1, in5430_2, pp53[19]);
    wire[0:0] s5431, in5431_1, in5431_2;
    wire c5431;
    assign in5431_1 = {pp57[15]};
    assign in5431_2 = {pp58[14]};
    Full_Adder FA_5431(s5431, c5431, in5431_1, in5431_2, pp56[16]);
    wire[0:0] s5432, in5432_1, in5432_2;
    wire c5432;
    assign in5432_1 = {pp60[12]};
    assign in5432_2 = {pp61[11]};
    Full_Adder FA_5432(s5432, c5432, in5432_1, in5432_2, pp59[13]);
    wire[0:0] s5433, in5433_1, in5433_2;
    wire c5433;
    assign in5433_1 = {pp63[9]};
    assign in5433_2 = {pp64[8]};
    Full_Adder FA_5433(s5433, c5433, in5433_1, in5433_2, pp62[10]);
    wire[0:0] s5434, in5434_1, in5434_2;
    wire c5434;
    assign in5434_1 = {pp66[6]};
    assign in5434_2 = {pp67[5]};
    Full_Adder FA_5434(s5434, c5434, in5434_1, in5434_2, pp65[7]);
    wire[0:0] s5435, in5435_1, in5435_2;
    wire c5435;
    assign in5435_1 = {pp69[3]};
    assign in5435_2 = {pp70[2]};
    Full_Adder FA_5435(s5435, c5435, in5435_1, in5435_2, pp68[4]);
    wire[0:0] s5436, in5436_1, in5436_2;
    wire c5436;
    assign in5436_1 = {pp72[0]};
    assign in5436_2 = {c1898};
    Full_Adder FA_5436(s5436, c5436, in5436_1, in5436_2, pp71[1]);
    wire[0:0] s5437, in5437_1, in5437_2;
    wire c5437;
    assign in5437_1 = {c1900};
    assign in5437_2 = {c1901};
    Full_Adder FA_5437(s5437, c5437, in5437_1, in5437_2, c1899);
    wire[0:0] s5438, in5438_1, in5438_2;
    wire c5438;
    assign in5438_1 = {c1903};
    assign in5438_2 = {c1904};
    Full_Adder FA_5438(s5438, c5438, in5438_1, in5438_2, c1902);
    wire[0:0] s5439, in5439_1, in5439_2;
    wire c5439;
    assign in5439_1 = {c1906};
    assign in5439_2 = {c1907};
    Full_Adder FA_5439(s5439, c5439, in5439_1, in5439_2, c1905);
    wire[0:0] s5440, in5440_1, in5440_2;
    wire c5440;
    assign in5440_1 = {c1909};
    assign in5440_2 = {c1910};
    Full_Adder FA_5440(s5440, c5440, in5440_1, in5440_2, c1908);
    wire[0:0] s5441, in5441_1, in5441_2;
    wire c5441;
    assign in5441_1 = {s1912[0]};
    assign in5441_2 = {s1913[0]};
    Full_Adder FA_5441(s5441, c5441, in5441_1, in5441_2, c1911);
    wire[0:0] s5442, in5442_1, in5442_2;
    wire c5442;
    assign in5442_1 = {s1915[0]};
    assign in5442_2 = {s1916[0]};
    Full_Adder FA_5442(s5442, c5442, in5442_1, in5442_2, s1914[0]);
    wire[0:0] s5443, in5443_1, in5443_2;
    wire c5443;
    assign in5443_1 = {s1918[0]};
    assign in5443_2 = {s1919[0]};
    Full_Adder FA_5443(s5443, c5443, in5443_1, in5443_2, s1917[0]);
    wire[0:0] s5444, in5444_1, in5444_2;
    wire c5444;
    assign in5444_1 = {s1921[0]};
    assign in5444_2 = {s1922[0]};
    Full_Adder FA_5444(s5444, c5444, in5444_1, in5444_2, s1920[0]);
    wire[0:0] s5445, in5445_1, in5445_2;
    wire c5445;
    assign in5445_1 = {s1924[0]};
    assign in5445_2 = {s1925[0]};
    Full_Adder FA_5445(s5445, c5445, in5445_1, in5445_2, s1923[0]);
    wire[0:0] s5446, in5446_1, in5446_2;
    wire c5446;
    assign in5446_1 = {pp48[25]};
    assign in5446_2 = {pp49[24]};
    Full_Adder FA_5446(s5446, c5446, in5446_1, in5446_2, pp47[26]);
    wire[0:0] s5447, in5447_1, in5447_2;
    wire c5447;
    assign in5447_1 = {pp51[22]};
    assign in5447_2 = {pp52[21]};
    Full_Adder FA_5447(s5447, c5447, in5447_1, in5447_2, pp50[23]);
    wire[0:0] s5448, in5448_1, in5448_2;
    wire c5448;
    assign in5448_1 = {pp54[19]};
    assign in5448_2 = {pp55[18]};
    Full_Adder FA_5448(s5448, c5448, in5448_1, in5448_2, pp53[20]);
    wire[0:0] s5449, in5449_1, in5449_2;
    wire c5449;
    assign in5449_1 = {pp57[16]};
    assign in5449_2 = {pp58[15]};
    Full_Adder FA_5449(s5449, c5449, in5449_1, in5449_2, pp56[17]);
    wire[0:0] s5450, in5450_1, in5450_2;
    wire c5450;
    assign in5450_1 = {pp60[13]};
    assign in5450_2 = {pp61[12]};
    Full_Adder FA_5450(s5450, c5450, in5450_1, in5450_2, pp59[14]);
    wire[0:0] s5451, in5451_1, in5451_2;
    wire c5451;
    assign in5451_1 = {pp63[10]};
    assign in5451_2 = {pp64[9]};
    Full_Adder FA_5451(s5451, c5451, in5451_1, in5451_2, pp62[11]);
    wire[0:0] s5452, in5452_1, in5452_2;
    wire c5452;
    assign in5452_1 = {pp66[7]};
    assign in5452_2 = {pp67[6]};
    Full_Adder FA_5452(s5452, c5452, in5452_1, in5452_2, pp65[8]);
    wire[0:0] s5453, in5453_1, in5453_2;
    wire c5453;
    assign in5453_1 = {pp69[4]};
    assign in5453_2 = {pp70[3]};
    Full_Adder FA_5453(s5453, c5453, in5453_1, in5453_2, pp68[5]);
    wire[0:0] s5454, in5454_1, in5454_2;
    wire c5454;
    assign in5454_1 = {pp72[1]};
    assign in5454_2 = {pp73[0]};
    Full_Adder FA_5454(s5454, c5454, in5454_1, in5454_2, pp71[2]);
    wire[0:0] s5455, in5455_1, in5455_2;
    wire c5455;
    assign in5455_1 = {c1913};
    assign in5455_2 = {c1914};
    Full_Adder FA_5455(s5455, c5455, in5455_1, in5455_2, c1912);
    wire[0:0] s5456, in5456_1, in5456_2;
    wire c5456;
    assign in5456_1 = {c1916};
    assign in5456_2 = {c1917};
    Full_Adder FA_5456(s5456, c5456, in5456_1, in5456_2, c1915);
    wire[0:0] s5457, in5457_1, in5457_2;
    wire c5457;
    assign in5457_1 = {c1919};
    assign in5457_2 = {c1920};
    Full_Adder FA_5457(s5457, c5457, in5457_1, in5457_2, c1918);
    wire[0:0] s5458, in5458_1, in5458_2;
    wire c5458;
    assign in5458_1 = {c1922};
    assign in5458_2 = {c1923};
    Full_Adder FA_5458(s5458, c5458, in5458_1, in5458_2, c1921);
    wire[0:0] s5459, in5459_1, in5459_2;
    wire c5459;
    assign in5459_1 = {c1925};
    assign in5459_2 = {c1926};
    Full_Adder FA_5459(s5459, c5459, in5459_1, in5459_2, c1924);
    wire[0:0] s5460, in5460_1, in5460_2;
    wire c5460;
    assign in5460_1 = {s1928[0]};
    assign in5460_2 = {s1929[0]};
    Full_Adder FA_5460(s5460, c5460, in5460_1, in5460_2, s1927[0]);
    wire[0:0] s5461, in5461_1, in5461_2;
    wire c5461;
    assign in5461_1 = {s1931[0]};
    assign in5461_2 = {s1932[0]};
    Full_Adder FA_5461(s5461, c5461, in5461_1, in5461_2, s1930[0]);
    wire[0:0] s5462, in5462_1, in5462_2;
    wire c5462;
    assign in5462_1 = {s1934[0]};
    assign in5462_2 = {s1935[0]};
    Full_Adder FA_5462(s5462, c5462, in5462_1, in5462_2, s1933[0]);
    wire[0:0] s5463, in5463_1, in5463_2;
    wire c5463;
    assign in5463_1 = {s1937[0]};
    assign in5463_2 = {s1938[0]};
    Full_Adder FA_5463(s5463, c5463, in5463_1, in5463_2, s1936[0]);
    wire[0:0] s5464, in5464_1, in5464_2;
    wire c5464;
    assign in5464_1 = {s1940[0]};
    assign in5464_2 = {s1941[0]};
    Full_Adder FA_5464(s5464, c5464, in5464_1, in5464_2, s1939[0]);
    wire[0:0] s5465, in5465_1, in5465_2;
    wire c5465;
    assign in5465_1 = {pp51[23]};
    assign in5465_2 = {pp52[22]};
    Full_Adder FA_5465(s5465, c5465, in5465_1, in5465_2, pp50[24]);
    wire[0:0] s5466, in5466_1, in5466_2;
    wire c5466;
    assign in5466_1 = {pp54[20]};
    assign in5466_2 = {pp55[19]};
    Full_Adder FA_5466(s5466, c5466, in5466_1, in5466_2, pp53[21]);
    wire[0:0] s5467, in5467_1, in5467_2;
    wire c5467;
    assign in5467_1 = {pp57[17]};
    assign in5467_2 = {pp58[16]};
    Full_Adder FA_5467(s5467, c5467, in5467_1, in5467_2, pp56[18]);
    wire[0:0] s5468, in5468_1, in5468_2;
    wire c5468;
    assign in5468_1 = {pp60[14]};
    assign in5468_2 = {pp61[13]};
    Full_Adder FA_5468(s5468, c5468, in5468_1, in5468_2, pp59[15]);
    wire[0:0] s5469, in5469_1, in5469_2;
    wire c5469;
    assign in5469_1 = {pp63[11]};
    assign in5469_2 = {pp64[10]};
    Full_Adder FA_5469(s5469, c5469, in5469_1, in5469_2, pp62[12]);
    wire[0:0] s5470, in5470_1, in5470_2;
    wire c5470;
    assign in5470_1 = {pp66[8]};
    assign in5470_2 = {pp67[7]};
    Full_Adder FA_5470(s5470, c5470, in5470_1, in5470_2, pp65[9]);
    wire[0:0] s5471, in5471_1, in5471_2;
    wire c5471;
    assign in5471_1 = {pp69[5]};
    assign in5471_2 = {pp70[4]};
    Full_Adder FA_5471(s5471, c5471, in5471_1, in5471_2, pp68[6]);
    wire[0:0] s5472, in5472_1, in5472_2;
    wire c5472;
    assign in5472_1 = {pp72[2]};
    assign in5472_2 = {pp73[1]};
    Full_Adder FA_5472(s5472, c5472, in5472_1, in5472_2, pp71[3]);
    wire[0:0] s5473, in5473_1, in5473_2;
    wire c5473;
    assign in5473_1 = {c1927};
    assign in5473_2 = {c1928};
    Full_Adder FA_5473(s5473, c5473, in5473_1, in5473_2, pp74[0]);
    wire[0:0] s5474, in5474_1, in5474_2;
    wire c5474;
    assign in5474_1 = {c1930};
    assign in5474_2 = {c1931};
    Full_Adder FA_5474(s5474, c5474, in5474_1, in5474_2, c1929);
    wire[0:0] s5475, in5475_1, in5475_2;
    wire c5475;
    assign in5475_1 = {c1933};
    assign in5475_2 = {c1934};
    Full_Adder FA_5475(s5475, c5475, in5475_1, in5475_2, c1932);
    wire[0:0] s5476, in5476_1, in5476_2;
    wire c5476;
    assign in5476_1 = {c1936};
    assign in5476_2 = {c1937};
    Full_Adder FA_5476(s5476, c5476, in5476_1, in5476_2, c1935);
    wire[0:0] s5477, in5477_1, in5477_2;
    wire c5477;
    assign in5477_1 = {c1939};
    assign in5477_2 = {c1940};
    Full_Adder FA_5477(s5477, c5477, in5477_1, in5477_2, c1938);
    wire[0:0] s5478, in5478_1, in5478_2;
    wire c5478;
    assign in5478_1 = {c1942};
    assign in5478_2 = {s1943[0]};
    Full_Adder FA_5478(s5478, c5478, in5478_1, in5478_2, c1941);
    wire[0:0] s5479, in5479_1, in5479_2;
    wire c5479;
    assign in5479_1 = {s1945[0]};
    assign in5479_2 = {s1946[0]};
    Full_Adder FA_5479(s5479, c5479, in5479_1, in5479_2, s1944[0]);
    wire[0:0] s5480, in5480_1, in5480_2;
    wire c5480;
    assign in5480_1 = {s1948[0]};
    assign in5480_2 = {s1949[0]};
    Full_Adder FA_5480(s5480, c5480, in5480_1, in5480_2, s1947[0]);
    wire[0:0] s5481, in5481_1, in5481_2;
    wire c5481;
    assign in5481_1 = {s1951[0]};
    assign in5481_2 = {s1952[0]};
    Full_Adder FA_5481(s5481, c5481, in5481_1, in5481_2, s1950[0]);
    wire[0:0] s5482, in5482_1, in5482_2;
    wire c5482;
    assign in5482_1 = {s1954[0]};
    assign in5482_2 = {s1955[0]};
    Full_Adder FA_5482(s5482, c5482, in5482_1, in5482_2, s1953[0]);
    wire[0:0] s5483, in5483_1, in5483_2;
    wire c5483;
    assign in5483_1 = {s1957[0]};
    assign in5483_2 = {s1958[0]};
    Full_Adder FA_5483(s5483, c5483, in5483_1, in5483_2, s1956[0]);
    wire[0:0] s5484, in5484_1, in5484_2;
    wire c5484;
    assign in5484_1 = {pp54[21]};
    assign in5484_2 = {pp55[20]};
    Full_Adder FA_5484(s5484, c5484, in5484_1, in5484_2, pp53[22]);
    wire[0:0] s5485, in5485_1, in5485_2;
    wire c5485;
    assign in5485_1 = {pp57[18]};
    assign in5485_2 = {pp58[17]};
    Full_Adder FA_5485(s5485, c5485, in5485_1, in5485_2, pp56[19]);
    wire[0:0] s5486, in5486_1, in5486_2;
    wire c5486;
    assign in5486_1 = {pp60[15]};
    assign in5486_2 = {pp61[14]};
    Full_Adder FA_5486(s5486, c5486, in5486_1, in5486_2, pp59[16]);
    wire[0:0] s5487, in5487_1, in5487_2;
    wire c5487;
    assign in5487_1 = {pp63[12]};
    assign in5487_2 = {pp64[11]};
    Full_Adder FA_5487(s5487, c5487, in5487_1, in5487_2, pp62[13]);
    wire[0:0] s5488, in5488_1, in5488_2;
    wire c5488;
    assign in5488_1 = {pp66[9]};
    assign in5488_2 = {pp67[8]};
    Full_Adder FA_5488(s5488, c5488, in5488_1, in5488_2, pp65[10]);
    wire[0:0] s5489, in5489_1, in5489_2;
    wire c5489;
    assign in5489_1 = {pp69[6]};
    assign in5489_2 = {pp70[5]};
    Full_Adder FA_5489(s5489, c5489, in5489_1, in5489_2, pp68[7]);
    wire[0:0] s5490, in5490_1, in5490_2;
    wire c5490;
    assign in5490_1 = {pp72[3]};
    assign in5490_2 = {pp73[2]};
    Full_Adder FA_5490(s5490, c5490, in5490_1, in5490_2, pp71[4]);
    wire[0:0] s5491, in5491_1, in5491_2;
    wire c5491;
    assign in5491_1 = {pp75[0]};
    assign in5491_2 = {c1943};
    Full_Adder FA_5491(s5491, c5491, in5491_1, in5491_2, pp74[1]);
    wire[0:0] s5492, in5492_1, in5492_2;
    wire c5492;
    assign in5492_1 = {c1945};
    assign in5492_2 = {c1946};
    Full_Adder FA_5492(s5492, c5492, in5492_1, in5492_2, c1944);
    wire[0:0] s5493, in5493_1, in5493_2;
    wire c5493;
    assign in5493_1 = {c1948};
    assign in5493_2 = {c1949};
    Full_Adder FA_5493(s5493, c5493, in5493_1, in5493_2, c1947);
    wire[0:0] s5494, in5494_1, in5494_2;
    wire c5494;
    assign in5494_1 = {c1951};
    assign in5494_2 = {c1952};
    Full_Adder FA_5494(s5494, c5494, in5494_1, in5494_2, c1950);
    wire[0:0] s5495, in5495_1, in5495_2;
    wire c5495;
    assign in5495_1 = {c1954};
    assign in5495_2 = {c1955};
    Full_Adder FA_5495(s5495, c5495, in5495_1, in5495_2, c1953);
    wire[0:0] s5496, in5496_1, in5496_2;
    wire c5496;
    assign in5496_1 = {c1957};
    assign in5496_2 = {c1958};
    Full_Adder FA_5496(s5496, c5496, in5496_1, in5496_2, c1956);
    wire[0:0] s5497, in5497_1, in5497_2;
    wire c5497;
    assign in5497_1 = {s1960[0]};
    assign in5497_2 = {s1961[0]};
    Full_Adder FA_5497(s5497, c5497, in5497_1, in5497_2, c1959);
    wire[0:0] s5498, in5498_1, in5498_2;
    wire c5498;
    assign in5498_1 = {s1963[0]};
    assign in5498_2 = {s1964[0]};
    Full_Adder FA_5498(s5498, c5498, in5498_1, in5498_2, s1962[0]);
    wire[0:0] s5499, in5499_1, in5499_2;
    wire c5499;
    assign in5499_1 = {s1966[0]};
    assign in5499_2 = {s1967[0]};
    Full_Adder FA_5499(s5499, c5499, in5499_1, in5499_2, s1965[0]);
    wire[0:0] s5500, in5500_1, in5500_2;
    wire c5500;
    assign in5500_1 = {s1969[0]};
    assign in5500_2 = {s1970[0]};
    Full_Adder FA_5500(s5500, c5500, in5500_1, in5500_2, s1968[0]);
    wire[0:0] s5501, in5501_1, in5501_2;
    wire c5501;
    assign in5501_1 = {s1972[0]};
    assign in5501_2 = {s1973[0]};
    Full_Adder FA_5501(s5501, c5501, in5501_1, in5501_2, s1971[0]);
    wire[0:0] s5502, in5502_1, in5502_2;
    wire c5502;
    assign in5502_1 = {s1975[0]};
    assign in5502_2 = {s1976[0]};
    Full_Adder FA_5502(s5502, c5502, in5502_1, in5502_2, s1974[0]);
    wire[0:0] s5503, in5503_1, in5503_2;
    wire c5503;
    assign in5503_1 = {pp57[19]};
    assign in5503_2 = {pp58[18]};
    Full_Adder FA_5503(s5503, c5503, in5503_1, in5503_2, pp56[20]);
    wire[0:0] s5504, in5504_1, in5504_2;
    wire c5504;
    assign in5504_1 = {pp60[16]};
    assign in5504_2 = {pp61[15]};
    Full_Adder FA_5504(s5504, c5504, in5504_1, in5504_2, pp59[17]);
    wire[0:0] s5505, in5505_1, in5505_2;
    wire c5505;
    assign in5505_1 = {pp63[13]};
    assign in5505_2 = {pp64[12]};
    Full_Adder FA_5505(s5505, c5505, in5505_1, in5505_2, pp62[14]);
    wire[0:0] s5506, in5506_1, in5506_2;
    wire c5506;
    assign in5506_1 = {pp66[10]};
    assign in5506_2 = {pp67[9]};
    Full_Adder FA_5506(s5506, c5506, in5506_1, in5506_2, pp65[11]);
    wire[0:0] s5507, in5507_1, in5507_2;
    wire c5507;
    assign in5507_1 = {pp69[7]};
    assign in5507_2 = {pp70[6]};
    Full_Adder FA_5507(s5507, c5507, in5507_1, in5507_2, pp68[8]);
    wire[0:0] s5508, in5508_1, in5508_2;
    wire c5508;
    assign in5508_1 = {pp72[4]};
    assign in5508_2 = {pp73[3]};
    Full_Adder FA_5508(s5508, c5508, in5508_1, in5508_2, pp71[5]);
    wire[0:0] s5509, in5509_1, in5509_2;
    wire c5509;
    assign in5509_1 = {pp75[1]};
    assign in5509_2 = {pp76[0]};
    Full_Adder FA_5509(s5509, c5509, in5509_1, in5509_2, pp74[2]);
    wire[0:0] s5510, in5510_1, in5510_2;
    wire c5510;
    assign in5510_1 = {c1961};
    assign in5510_2 = {c1962};
    Full_Adder FA_5510(s5510, c5510, in5510_1, in5510_2, c1960);
    wire[0:0] s5511, in5511_1, in5511_2;
    wire c5511;
    assign in5511_1 = {c1964};
    assign in5511_2 = {c1965};
    Full_Adder FA_5511(s5511, c5511, in5511_1, in5511_2, c1963);
    wire[0:0] s5512, in5512_1, in5512_2;
    wire c5512;
    assign in5512_1 = {c1967};
    assign in5512_2 = {c1968};
    Full_Adder FA_5512(s5512, c5512, in5512_1, in5512_2, c1966);
    wire[0:0] s5513, in5513_1, in5513_2;
    wire c5513;
    assign in5513_1 = {c1970};
    assign in5513_2 = {c1971};
    Full_Adder FA_5513(s5513, c5513, in5513_1, in5513_2, c1969);
    wire[0:0] s5514, in5514_1, in5514_2;
    wire c5514;
    assign in5514_1 = {c1973};
    assign in5514_2 = {c1974};
    Full_Adder FA_5514(s5514, c5514, in5514_1, in5514_2, c1972);
    wire[0:0] s5515, in5515_1, in5515_2;
    wire c5515;
    assign in5515_1 = {c1976};
    assign in5515_2 = {c1977};
    Full_Adder FA_5515(s5515, c5515, in5515_1, in5515_2, c1975);
    wire[0:0] s5516, in5516_1, in5516_2;
    wire c5516;
    assign in5516_1 = {s1979[0]};
    assign in5516_2 = {s1980[0]};
    Full_Adder FA_5516(s5516, c5516, in5516_1, in5516_2, s1978[0]);
    wire[0:0] s5517, in5517_1, in5517_2;
    wire c5517;
    assign in5517_1 = {s1982[0]};
    assign in5517_2 = {s1983[0]};
    Full_Adder FA_5517(s5517, c5517, in5517_1, in5517_2, s1981[0]);
    wire[0:0] s5518, in5518_1, in5518_2;
    wire c5518;
    assign in5518_1 = {s1985[0]};
    assign in5518_2 = {s1986[0]};
    Full_Adder FA_5518(s5518, c5518, in5518_1, in5518_2, s1984[0]);
    wire[0:0] s5519, in5519_1, in5519_2;
    wire c5519;
    assign in5519_1 = {s1988[0]};
    assign in5519_2 = {s1989[0]};
    Full_Adder FA_5519(s5519, c5519, in5519_1, in5519_2, s1987[0]);
    wire[0:0] s5520, in5520_1, in5520_2;
    wire c5520;
    assign in5520_1 = {s1991[0]};
    assign in5520_2 = {s1992[0]};
    Full_Adder FA_5520(s5520, c5520, in5520_1, in5520_2, s1990[0]);
    wire[0:0] s5521, in5521_1, in5521_2;
    wire c5521;
    assign in5521_1 = {s1994[0]};
    assign in5521_2 = {s1995[0]};
    Full_Adder FA_5521(s5521, c5521, in5521_1, in5521_2, s1993[0]);
    wire[0:0] s5522, in5522_1, in5522_2;
    wire c5522;
    assign in5522_1 = {pp60[17]};
    assign in5522_2 = {pp61[16]};
    Full_Adder FA_5522(s5522, c5522, in5522_1, in5522_2, pp59[18]);
    wire[0:0] s5523, in5523_1, in5523_2;
    wire c5523;
    assign in5523_1 = {pp63[14]};
    assign in5523_2 = {pp64[13]};
    Full_Adder FA_5523(s5523, c5523, in5523_1, in5523_2, pp62[15]);
    wire[0:0] s5524, in5524_1, in5524_2;
    wire c5524;
    assign in5524_1 = {pp66[11]};
    assign in5524_2 = {pp67[10]};
    Full_Adder FA_5524(s5524, c5524, in5524_1, in5524_2, pp65[12]);
    wire[0:0] s5525, in5525_1, in5525_2;
    wire c5525;
    assign in5525_1 = {pp69[8]};
    assign in5525_2 = {pp70[7]};
    Full_Adder FA_5525(s5525, c5525, in5525_1, in5525_2, pp68[9]);
    wire[0:0] s5526, in5526_1, in5526_2;
    wire c5526;
    assign in5526_1 = {pp72[5]};
    assign in5526_2 = {pp73[4]};
    Full_Adder FA_5526(s5526, c5526, in5526_1, in5526_2, pp71[6]);
    wire[0:0] s5527, in5527_1, in5527_2;
    wire c5527;
    assign in5527_1 = {pp75[2]};
    assign in5527_2 = {pp76[1]};
    Full_Adder FA_5527(s5527, c5527, in5527_1, in5527_2, pp74[3]);
    wire[0:0] s5528, in5528_1, in5528_2;
    wire c5528;
    assign in5528_1 = {c1978};
    assign in5528_2 = {c1979};
    Full_Adder FA_5528(s5528, c5528, in5528_1, in5528_2, pp77[0]);
    wire[0:0] s5529, in5529_1, in5529_2;
    wire c5529;
    assign in5529_1 = {c1981};
    assign in5529_2 = {c1982};
    Full_Adder FA_5529(s5529, c5529, in5529_1, in5529_2, c1980);
    wire[0:0] s5530, in5530_1, in5530_2;
    wire c5530;
    assign in5530_1 = {c1984};
    assign in5530_2 = {c1985};
    Full_Adder FA_5530(s5530, c5530, in5530_1, in5530_2, c1983);
    wire[0:0] s5531, in5531_1, in5531_2;
    wire c5531;
    assign in5531_1 = {c1987};
    assign in5531_2 = {c1988};
    Full_Adder FA_5531(s5531, c5531, in5531_1, in5531_2, c1986);
    wire[0:0] s5532, in5532_1, in5532_2;
    wire c5532;
    assign in5532_1 = {c1990};
    assign in5532_2 = {c1991};
    Full_Adder FA_5532(s5532, c5532, in5532_1, in5532_2, c1989);
    wire[0:0] s5533, in5533_1, in5533_2;
    wire c5533;
    assign in5533_1 = {c1993};
    assign in5533_2 = {c1994};
    Full_Adder FA_5533(s5533, c5533, in5533_1, in5533_2, c1992);
    wire[0:0] s5534, in5534_1, in5534_2;
    wire c5534;
    assign in5534_1 = {c1996};
    assign in5534_2 = {s1997[0]};
    Full_Adder FA_5534(s5534, c5534, in5534_1, in5534_2, c1995);
    wire[0:0] s5535, in5535_1, in5535_2;
    wire c5535;
    assign in5535_1 = {s1999[0]};
    assign in5535_2 = {s2000[0]};
    Full_Adder FA_5535(s5535, c5535, in5535_1, in5535_2, s1998[0]);
    wire[0:0] s5536, in5536_1, in5536_2;
    wire c5536;
    assign in5536_1 = {s2002[0]};
    assign in5536_2 = {s2003[0]};
    Full_Adder FA_5536(s5536, c5536, in5536_1, in5536_2, s2001[0]);
    wire[0:0] s5537, in5537_1, in5537_2;
    wire c5537;
    assign in5537_1 = {s2005[0]};
    assign in5537_2 = {s2006[0]};
    Full_Adder FA_5537(s5537, c5537, in5537_1, in5537_2, s2004[0]);
    wire[0:0] s5538, in5538_1, in5538_2;
    wire c5538;
    assign in5538_1 = {s2008[0]};
    assign in5538_2 = {s2009[0]};
    Full_Adder FA_5538(s5538, c5538, in5538_1, in5538_2, s2007[0]);
    wire[0:0] s5539, in5539_1, in5539_2;
    wire c5539;
    assign in5539_1 = {s2011[0]};
    assign in5539_2 = {s2012[0]};
    Full_Adder FA_5539(s5539, c5539, in5539_1, in5539_2, s2010[0]);
    wire[0:0] s5540, in5540_1, in5540_2;
    wire c5540;
    assign in5540_1 = {s2014[0]};
    assign in5540_2 = {s2015[0]};
    Full_Adder FA_5540(s5540, c5540, in5540_1, in5540_2, s2013[0]);
    wire[0:0] s5541, in5541_1, in5541_2;
    wire c5541;
    assign in5541_1 = {pp63[15]};
    assign in5541_2 = {pp64[14]};
    Full_Adder FA_5541(s5541, c5541, in5541_1, in5541_2, pp62[16]);
    wire[0:0] s5542, in5542_1, in5542_2;
    wire c5542;
    assign in5542_1 = {pp66[12]};
    assign in5542_2 = {pp67[11]};
    Full_Adder FA_5542(s5542, c5542, in5542_1, in5542_2, pp65[13]);
    wire[0:0] s5543, in5543_1, in5543_2;
    wire c5543;
    assign in5543_1 = {pp69[9]};
    assign in5543_2 = {pp70[8]};
    Full_Adder FA_5543(s5543, c5543, in5543_1, in5543_2, pp68[10]);
    wire[0:0] s5544, in5544_1, in5544_2;
    wire c5544;
    assign in5544_1 = {pp72[6]};
    assign in5544_2 = {pp73[5]};
    Full_Adder FA_5544(s5544, c5544, in5544_1, in5544_2, pp71[7]);
    wire[0:0] s5545, in5545_1, in5545_2;
    wire c5545;
    assign in5545_1 = {pp75[3]};
    assign in5545_2 = {pp76[2]};
    Full_Adder FA_5545(s5545, c5545, in5545_1, in5545_2, pp74[4]);
    wire[0:0] s5546, in5546_1, in5546_2;
    wire c5546;
    assign in5546_1 = {pp78[0]};
    assign in5546_2 = {c1997};
    Full_Adder FA_5546(s5546, c5546, in5546_1, in5546_2, pp77[1]);
    wire[0:0] s5547, in5547_1, in5547_2;
    wire c5547;
    assign in5547_1 = {c1999};
    assign in5547_2 = {c2000};
    Full_Adder FA_5547(s5547, c5547, in5547_1, in5547_2, c1998);
    wire[0:0] s5548, in5548_1, in5548_2;
    wire c5548;
    assign in5548_1 = {c2002};
    assign in5548_2 = {c2003};
    Full_Adder FA_5548(s5548, c5548, in5548_1, in5548_2, c2001);
    wire[0:0] s5549, in5549_1, in5549_2;
    wire c5549;
    assign in5549_1 = {c2005};
    assign in5549_2 = {c2006};
    Full_Adder FA_5549(s5549, c5549, in5549_1, in5549_2, c2004);
    wire[0:0] s5550, in5550_1, in5550_2;
    wire c5550;
    assign in5550_1 = {c2008};
    assign in5550_2 = {c2009};
    Full_Adder FA_5550(s5550, c5550, in5550_1, in5550_2, c2007);
    wire[0:0] s5551, in5551_1, in5551_2;
    wire c5551;
    assign in5551_1 = {c2011};
    assign in5551_2 = {c2012};
    Full_Adder FA_5551(s5551, c5551, in5551_1, in5551_2, c2010);
    wire[0:0] s5552, in5552_1, in5552_2;
    wire c5552;
    assign in5552_1 = {c2014};
    assign in5552_2 = {c2015};
    Full_Adder FA_5552(s5552, c5552, in5552_1, in5552_2, c2013);
    wire[0:0] s5553, in5553_1, in5553_2;
    wire c5553;
    assign in5553_1 = {s2017[0]};
    assign in5553_2 = {s2018[0]};
    Full_Adder FA_5553(s5553, c5553, in5553_1, in5553_2, c2016);
    wire[0:0] s5554, in5554_1, in5554_2;
    wire c5554;
    assign in5554_1 = {s2020[0]};
    assign in5554_2 = {s2021[0]};
    Full_Adder FA_5554(s5554, c5554, in5554_1, in5554_2, s2019[0]);
    wire[0:0] s5555, in5555_1, in5555_2;
    wire c5555;
    assign in5555_1 = {s2023[0]};
    assign in5555_2 = {s2024[0]};
    Full_Adder FA_5555(s5555, c5555, in5555_1, in5555_2, s2022[0]);
    wire[0:0] s5556, in5556_1, in5556_2;
    wire c5556;
    assign in5556_1 = {s2026[0]};
    assign in5556_2 = {s2027[0]};
    Full_Adder FA_5556(s5556, c5556, in5556_1, in5556_2, s2025[0]);
    wire[0:0] s5557, in5557_1, in5557_2;
    wire c5557;
    assign in5557_1 = {s2029[0]};
    assign in5557_2 = {s2030[0]};
    Full_Adder FA_5557(s5557, c5557, in5557_1, in5557_2, s2028[0]);
    wire[0:0] s5558, in5558_1, in5558_2;
    wire c5558;
    assign in5558_1 = {s2032[0]};
    assign in5558_2 = {s2033[0]};
    Full_Adder FA_5558(s5558, c5558, in5558_1, in5558_2, s2031[0]);
    wire[0:0] s5559, in5559_1, in5559_2;
    wire c5559;
    assign in5559_1 = {s2035[0]};
    assign in5559_2 = {s2036[0]};
    Full_Adder FA_5559(s5559, c5559, in5559_1, in5559_2, s2034[0]);
    wire[0:0] s5560, in5560_1, in5560_2;
    wire c5560;
    assign in5560_1 = {pp66[13]};
    assign in5560_2 = {pp67[12]};
    Full_Adder FA_5560(s5560, c5560, in5560_1, in5560_2, pp65[14]);
    wire[0:0] s5561, in5561_1, in5561_2;
    wire c5561;
    assign in5561_1 = {pp69[10]};
    assign in5561_2 = {pp70[9]};
    Full_Adder FA_5561(s5561, c5561, in5561_1, in5561_2, pp68[11]);
    wire[0:0] s5562, in5562_1, in5562_2;
    wire c5562;
    assign in5562_1 = {pp72[7]};
    assign in5562_2 = {pp73[6]};
    Full_Adder FA_5562(s5562, c5562, in5562_1, in5562_2, pp71[8]);
    wire[0:0] s5563, in5563_1, in5563_2;
    wire c5563;
    assign in5563_1 = {pp75[4]};
    assign in5563_2 = {pp76[3]};
    Full_Adder FA_5563(s5563, c5563, in5563_1, in5563_2, pp74[5]);
    wire[0:0] s5564, in5564_1, in5564_2;
    wire c5564;
    assign in5564_1 = {pp78[1]};
    assign in5564_2 = {pp79[0]};
    Full_Adder FA_5564(s5564, c5564, in5564_1, in5564_2, pp77[2]);
    wire[0:0] s5565, in5565_1, in5565_2;
    wire c5565;
    assign in5565_1 = {c2018};
    assign in5565_2 = {c2019};
    Full_Adder FA_5565(s5565, c5565, in5565_1, in5565_2, c2017);
    wire[0:0] s5566, in5566_1, in5566_2;
    wire c5566;
    assign in5566_1 = {c2021};
    assign in5566_2 = {c2022};
    Full_Adder FA_5566(s5566, c5566, in5566_1, in5566_2, c2020);
    wire[0:0] s5567, in5567_1, in5567_2;
    wire c5567;
    assign in5567_1 = {c2024};
    assign in5567_2 = {c2025};
    Full_Adder FA_5567(s5567, c5567, in5567_1, in5567_2, c2023);
    wire[0:0] s5568, in5568_1, in5568_2;
    wire c5568;
    assign in5568_1 = {c2027};
    assign in5568_2 = {c2028};
    Full_Adder FA_5568(s5568, c5568, in5568_1, in5568_2, c2026);
    wire[0:0] s5569, in5569_1, in5569_2;
    wire c5569;
    assign in5569_1 = {c2030};
    assign in5569_2 = {c2031};
    Full_Adder FA_5569(s5569, c5569, in5569_1, in5569_2, c2029);
    wire[0:0] s5570, in5570_1, in5570_2;
    wire c5570;
    assign in5570_1 = {c2033};
    assign in5570_2 = {c2034};
    Full_Adder FA_5570(s5570, c5570, in5570_1, in5570_2, c2032);
    wire[0:0] s5571, in5571_1, in5571_2;
    wire c5571;
    assign in5571_1 = {c2036};
    assign in5571_2 = {c2037};
    Full_Adder FA_5571(s5571, c5571, in5571_1, in5571_2, c2035);
    wire[0:0] s5572, in5572_1, in5572_2;
    wire c5572;
    assign in5572_1 = {s2039[0]};
    assign in5572_2 = {s2040[0]};
    Full_Adder FA_5572(s5572, c5572, in5572_1, in5572_2, s2038[0]);
    wire[0:0] s5573, in5573_1, in5573_2;
    wire c5573;
    assign in5573_1 = {s2042[0]};
    assign in5573_2 = {s2043[0]};
    Full_Adder FA_5573(s5573, c5573, in5573_1, in5573_2, s2041[0]);
    wire[0:0] s5574, in5574_1, in5574_2;
    wire c5574;
    assign in5574_1 = {s2045[0]};
    assign in5574_2 = {s2046[0]};
    Full_Adder FA_5574(s5574, c5574, in5574_1, in5574_2, s2044[0]);
    wire[0:0] s5575, in5575_1, in5575_2;
    wire c5575;
    assign in5575_1 = {s2048[0]};
    assign in5575_2 = {s2049[0]};
    Full_Adder FA_5575(s5575, c5575, in5575_1, in5575_2, s2047[0]);
    wire[0:0] s5576, in5576_1, in5576_2;
    wire c5576;
    assign in5576_1 = {s2051[0]};
    assign in5576_2 = {s2052[0]};
    Full_Adder FA_5576(s5576, c5576, in5576_1, in5576_2, s2050[0]);
    wire[0:0] s5577, in5577_1, in5577_2;
    wire c5577;
    assign in5577_1 = {s2054[0]};
    assign in5577_2 = {s2055[0]};
    Full_Adder FA_5577(s5577, c5577, in5577_1, in5577_2, s2053[0]);
    wire[0:0] s5578, in5578_1, in5578_2;
    wire c5578;
    assign in5578_1 = {s2057[0]};
    assign in5578_2 = {s2058[0]};
    Full_Adder FA_5578(s5578, c5578, in5578_1, in5578_2, s2056[0]);
    wire[0:0] s5579, in5579_1, in5579_2;
    wire c5579;
    assign in5579_1 = {pp69[11]};
    assign in5579_2 = {pp70[10]};
    Full_Adder FA_5579(s5579, c5579, in5579_1, in5579_2, pp68[12]);
    wire[0:0] s5580, in5580_1, in5580_2;
    wire c5580;
    assign in5580_1 = {pp72[8]};
    assign in5580_2 = {pp73[7]};
    Full_Adder FA_5580(s5580, c5580, in5580_1, in5580_2, pp71[9]);
    wire[0:0] s5581, in5581_1, in5581_2;
    wire c5581;
    assign in5581_1 = {pp75[5]};
    assign in5581_2 = {pp76[4]};
    Full_Adder FA_5581(s5581, c5581, in5581_1, in5581_2, pp74[6]);
    wire[0:0] s5582, in5582_1, in5582_2;
    wire c5582;
    assign in5582_1 = {pp78[2]};
    assign in5582_2 = {pp79[1]};
    Full_Adder FA_5582(s5582, c5582, in5582_1, in5582_2, pp77[3]);
    wire[0:0] s5583, in5583_1, in5583_2;
    wire c5583;
    assign in5583_1 = {c2038};
    assign in5583_2 = {c2039};
    Full_Adder FA_5583(s5583, c5583, in5583_1, in5583_2, pp80[0]);
    wire[0:0] s5584, in5584_1, in5584_2;
    wire c5584;
    assign in5584_1 = {c2041};
    assign in5584_2 = {c2042};
    Full_Adder FA_5584(s5584, c5584, in5584_1, in5584_2, c2040);
    wire[0:0] s5585, in5585_1, in5585_2;
    wire c5585;
    assign in5585_1 = {c2044};
    assign in5585_2 = {c2045};
    Full_Adder FA_5585(s5585, c5585, in5585_1, in5585_2, c2043);
    wire[0:0] s5586, in5586_1, in5586_2;
    wire c5586;
    assign in5586_1 = {c2047};
    assign in5586_2 = {c2048};
    Full_Adder FA_5586(s5586, c5586, in5586_1, in5586_2, c2046);
    wire[0:0] s5587, in5587_1, in5587_2;
    wire c5587;
    assign in5587_1 = {c2050};
    assign in5587_2 = {c2051};
    Full_Adder FA_5587(s5587, c5587, in5587_1, in5587_2, c2049);
    wire[0:0] s5588, in5588_1, in5588_2;
    wire c5588;
    assign in5588_1 = {c2053};
    assign in5588_2 = {c2054};
    Full_Adder FA_5588(s5588, c5588, in5588_1, in5588_2, c2052);
    wire[0:0] s5589, in5589_1, in5589_2;
    wire c5589;
    assign in5589_1 = {c2056};
    assign in5589_2 = {c2057};
    Full_Adder FA_5589(s5589, c5589, in5589_1, in5589_2, c2055);
    wire[0:0] s5590, in5590_1, in5590_2;
    wire c5590;
    assign in5590_1 = {c2059};
    assign in5590_2 = {s2060[0]};
    Full_Adder FA_5590(s5590, c5590, in5590_1, in5590_2, c2058);
    wire[0:0] s5591, in5591_1, in5591_2;
    wire c5591;
    assign in5591_1 = {s2062[0]};
    assign in5591_2 = {s2063[0]};
    Full_Adder FA_5591(s5591, c5591, in5591_1, in5591_2, s2061[0]);
    wire[0:0] s5592, in5592_1, in5592_2;
    wire c5592;
    assign in5592_1 = {s2065[0]};
    assign in5592_2 = {s2066[0]};
    Full_Adder FA_5592(s5592, c5592, in5592_1, in5592_2, s2064[0]);
    wire[0:0] s5593, in5593_1, in5593_2;
    wire c5593;
    assign in5593_1 = {s2068[0]};
    assign in5593_2 = {s2069[0]};
    Full_Adder FA_5593(s5593, c5593, in5593_1, in5593_2, s2067[0]);
    wire[0:0] s5594, in5594_1, in5594_2;
    wire c5594;
    assign in5594_1 = {s2071[0]};
    assign in5594_2 = {s2072[0]};
    Full_Adder FA_5594(s5594, c5594, in5594_1, in5594_2, s2070[0]);
    wire[0:0] s5595, in5595_1, in5595_2;
    wire c5595;
    assign in5595_1 = {s2074[0]};
    assign in5595_2 = {s2075[0]};
    Full_Adder FA_5595(s5595, c5595, in5595_1, in5595_2, s2073[0]);
    wire[0:0] s5596, in5596_1, in5596_2;
    wire c5596;
    assign in5596_1 = {s2077[0]};
    assign in5596_2 = {s2078[0]};
    Full_Adder FA_5596(s5596, c5596, in5596_1, in5596_2, s2076[0]);
    wire[0:0] s5597, in5597_1, in5597_2;
    wire c5597;
    assign in5597_1 = {s2080[0]};
    assign in5597_2 = {s2081[0]};
    Full_Adder FA_5597(s5597, c5597, in5597_1, in5597_2, s2079[0]);
    wire[0:0] s5598, in5598_1, in5598_2;
    wire c5598;
    assign in5598_1 = {pp72[9]};
    assign in5598_2 = {pp73[8]};
    Full_Adder FA_5598(s5598, c5598, in5598_1, in5598_2, pp71[10]);
    wire[0:0] s5599, in5599_1, in5599_2;
    wire c5599;
    assign in5599_1 = {pp75[6]};
    assign in5599_2 = {pp76[5]};
    Full_Adder FA_5599(s5599, c5599, in5599_1, in5599_2, pp74[7]);
    wire[0:0] s5600, in5600_1, in5600_2;
    wire c5600;
    assign in5600_1 = {pp78[3]};
    assign in5600_2 = {pp79[2]};
    Full_Adder FA_5600(s5600, c5600, in5600_1, in5600_2, pp77[4]);
    wire[0:0] s5601, in5601_1, in5601_2;
    wire c5601;
    assign in5601_1 = {pp81[0]};
    assign in5601_2 = {c2060};
    Full_Adder FA_5601(s5601, c5601, in5601_1, in5601_2, pp80[1]);
    wire[0:0] s5602, in5602_1, in5602_2;
    wire c5602;
    assign in5602_1 = {c2062};
    assign in5602_2 = {c2063};
    Full_Adder FA_5602(s5602, c5602, in5602_1, in5602_2, c2061);
    wire[0:0] s5603, in5603_1, in5603_2;
    wire c5603;
    assign in5603_1 = {c2065};
    assign in5603_2 = {c2066};
    Full_Adder FA_5603(s5603, c5603, in5603_1, in5603_2, c2064);
    wire[0:0] s5604, in5604_1, in5604_2;
    wire c5604;
    assign in5604_1 = {c2068};
    assign in5604_2 = {c2069};
    Full_Adder FA_5604(s5604, c5604, in5604_1, in5604_2, c2067);
    wire[0:0] s5605, in5605_1, in5605_2;
    wire c5605;
    assign in5605_1 = {c2071};
    assign in5605_2 = {c2072};
    Full_Adder FA_5605(s5605, c5605, in5605_1, in5605_2, c2070);
    wire[0:0] s5606, in5606_1, in5606_2;
    wire c5606;
    assign in5606_1 = {c2074};
    assign in5606_2 = {c2075};
    Full_Adder FA_5606(s5606, c5606, in5606_1, in5606_2, c2073);
    wire[0:0] s5607, in5607_1, in5607_2;
    wire c5607;
    assign in5607_1 = {c2077};
    assign in5607_2 = {c2078};
    Full_Adder FA_5607(s5607, c5607, in5607_1, in5607_2, c2076);
    wire[0:0] s5608, in5608_1, in5608_2;
    wire c5608;
    assign in5608_1 = {c2080};
    assign in5608_2 = {c2081};
    Full_Adder FA_5608(s5608, c5608, in5608_1, in5608_2, c2079);
    wire[0:0] s5609, in5609_1, in5609_2;
    wire c5609;
    assign in5609_1 = {s2083[0]};
    assign in5609_2 = {s2084[0]};
    Full_Adder FA_5609(s5609, c5609, in5609_1, in5609_2, c2082);
    wire[0:0] s5610, in5610_1, in5610_2;
    wire c5610;
    assign in5610_1 = {s2086[0]};
    assign in5610_2 = {s2087[0]};
    Full_Adder FA_5610(s5610, c5610, in5610_1, in5610_2, s2085[0]);
    wire[0:0] s5611, in5611_1, in5611_2;
    wire c5611;
    assign in5611_1 = {s2089[0]};
    assign in5611_2 = {s2090[0]};
    Full_Adder FA_5611(s5611, c5611, in5611_1, in5611_2, s2088[0]);
    wire[0:0] s5612, in5612_1, in5612_2;
    wire c5612;
    assign in5612_1 = {s2092[0]};
    assign in5612_2 = {s2093[0]};
    Full_Adder FA_5612(s5612, c5612, in5612_1, in5612_2, s2091[0]);
    wire[0:0] s5613, in5613_1, in5613_2;
    wire c5613;
    assign in5613_1 = {s2095[0]};
    assign in5613_2 = {s2096[0]};
    Full_Adder FA_5613(s5613, c5613, in5613_1, in5613_2, s2094[0]);
    wire[0:0] s5614, in5614_1, in5614_2;
    wire c5614;
    assign in5614_1 = {s2098[0]};
    assign in5614_2 = {s2099[0]};
    Full_Adder FA_5614(s5614, c5614, in5614_1, in5614_2, s2097[0]);
    wire[0:0] s5615, in5615_1, in5615_2;
    wire c5615;
    assign in5615_1 = {s2101[0]};
    assign in5615_2 = {s2102[0]};
    Full_Adder FA_5615(s5615, c5615, in5615_1, in5615_2, s2100[0]);
    wire[0:0] s5616, in5616_1, in5616_2;
    wire c5616;
    assign in5616_1 = {s2104[0]};
    assign in5616_2 = {s2105[0]};
    Full_Adder FA_5616(s5616, c5616, in5616_1, in5616_2, s2103[0]);
    wire[0:0] s5617, in5617_1, in5617_2;
    wire c5617;
    assign in5617_1 = {pp75[7]};
    assign in5617_2 = {pp76[6]};
    Full_Adder FA_5617(s5617, c5617, in5617_1, in5617_2, pp74[8]);
    wire[0:0] s5618, in5618_1, in5618_2;
    wire c5618;
    assign in5618_1 = {pp78[4]};
    assign in5618_2 = {pp79[3]};
    Full_Adder FA_5618(s5618, c5618, in5618_1, in5618_2, pp77[5]);
    wire[0:0] s5619, in5619_1, in5619_2;
    wire c5619;
    assign in5619_1 = {pp81[1]};
    assign in5619_2 = {pp82[0]};
    Full_Adder FA_5619(s5619, c5619, in5619_1, in5619_2, pp80[2]);
    wire[0:0] s5620, in5620_1, in5620_2;
    wire c5620;
    assign in5620_1 = {c2084};
    assign in5620_2 = {c2085};
    Full_Adder FA_5620(s5620, c5620, in5620_1, in5620_2, c2083);
    wire[0:0] s5621, in5621_1, in5621_2;
    wire c5621;
    assign in5621_1 = {c2087};
    assign in5621_2 = {c2088};
    Full_Adder FA_5621(s5621, c5621, in5621_1, in5621_2, c2086);
    wire[0:0] s5622, in5622_1, in5622_2;
    wire c5622;
    assign in5622_1 = {c2090};
    assign in5622_2 = {c2091};
    Full_Adder FA_5622(s5622, c5622, in5622_1, in5622_2, c2089);
    wire[0:0] s5623, in5623_1, in5623_2;
    wire c5623;
    assign in5623_1 = {c2093};
    assign in5623_2 = {c2094};
    Full_Adder FA_5623(s5623, c5623, in5623_1, in5623_2, c2092);
    wire[0:0] s5624, in5624_1, in5624_2;
    wire c5624;
    assign in5624_1 = {c2096};
    assign in5624_2 = {c2097};
    Full_Adder FA_5624(s5624, c5624, in5624_1, in5624_2, c2095);
    wire[0:0] s5625, in5625_1, in5625_2;
    wire c5625;
    assign in5625_1 = {c2099};
    assign in5625_2 = {c2100};
    Full_Adder FA_5625(s5625, c5625, in5625_1, in5625_2, c2098);
    wire[0:0] s5626, in5626_1, in5626_2;
    wire c5626;
    assign in5626_1 = {c2102};
    assign in5626_2 = {c2103};
    Full_Adder FA_5626(s5626, c5626, in5626_1, in5626_2, c2101);
    wire[0:0] s5627, in5627_1, in5627_2;
    wire c5627;
    assign in5627_1 = {c2105};
    assign in5627_2 = {c2106};
    Full_Adder FA_5627(s5627, c5627, in5627_1, in5627_2, c2104);
    wire[0:0] s5628, in5628_1, in5628_2;
    wire c5628;
    assign in5628_1 = {s2108[0]};
    assign in5628_2 = {s2109[0]};
    Full_Adder FA_5628(s5628, c5628, in5628_1, in5628_2, s2107[0]);
    wire[0:0] s5629, in5629_1, in5629_2;
    wire c5629;
    assign in5629_1 = {s2111[0]};
    assign in5629_2 = {s2112[0]};
    Full_Adder FA_5629(s5629, c5629, in5629_1, in5629_2, s2110[0]);
    wire[0:0] s5630, in5630_1, in5630_2;
    wire c5630;
    assign in5630_1 = {s2114[0]};
    assign in5630_2 = {s2115[0]};
    Full_Adder FA_5630(s5630, c5630, in5630_1, in5630_2, s2113[0]);
    wire[0:0] s5631, in5631_1, in5631_2;
    wire c5631;
    assign in5631_1 = {s2117[0]};
    assign in5631_2 = {s2118[0]};
    Full_Adder FA_5631(s5631, c5631, in5631_1, in5631_2, s2116[0]);
    wire[0:0] s5632, in5632_1, in5632_2;
    wire c5632;
    assign in5632_1 = {s2120[0]};
    assign in5632_2 = {s2121[0]};
    Full_Adder FA_5632(s5632, c5632, in5632_1, in5632_2, s2119[0]);
    wire[0:0] s5633, in5633_1, in5633_2;
    wire c5633;
    assign in5633_1 = {s2123[0]};
    assign in5633_2 = {s2124[0]};
    Full_Adder FA_5633(s5633, c5633, in5633_1, in5633_2, s2122[0]);
    wire[0:0] s5634, in5634_1, in5634_2;
    wire c5634;
    assign in5634_1 = {s2126[0]};
    assign in5634_2 = {s2127[0]};
    Full_Adder FA_5634(s5634, c5634, in5634_1, in5634_2, s2125[0]);
    wire[0:0] s5635, in5635_1, in5635_2;
    wire c5635;
    assign in5635_1 = {s2129[0]};
    assign in5635_2 = {s2130[0]};
    Full_Adder FA_5635(s5635, c5635, in5635_1, in5635_2, s2128[0]);
    wire[0:0] s5636, in5636_1, in5636_2;
    wire c5636;
    assign in5636_1 = {pp78[5]};
    assign in5636_2 = {pp79[4]};
    Full_Adder FA_5636(s5636, c5636, in5636_1, in5636_2, pp77[6]);
    wire[0:0] s5637, in5637_1, in5637_2;
    wire c5637;
    assign in5637_1 = {pp81[2]};
    assign in5637_2 = {pp82[1]};
    Full_Adder FA_5637(s5637, c5637, in5637_1, in5637_2, pp80[3]);
    wire[0:0] s5638, in5638_1, in5638_2;
    wire c5638;
    assign in5638_1 = {c2107};
    assign in5638_2 = {c2108};
    Full_Adder FA_5638(s5638, c5638, in5638_1, in5638_2, pp83[0]);
    wire[0:0] s5639, in5639_1, in5639_2;
    wire c5639;
    assign in5639_1 = {c2110};
    assign in5639_2 = {c2111};
    Full_Adder FA_5639(s5639, c5639, in5639_1, in5639_2, c2109);
    wire[0:0] s5640, in5640_1, in5640_2;
    wire c5640;
    assign in5640_1 = {c2113};
    assign in5640_2 = {c2114};
    Full_Adder FA_5640(s5640, c5640, in5640_1, in5640_2, c2112);
    wire[0:0] s5641, in5641_1, in5641_2;
    wire c5641;
    assign in5641_1 = {c2116};
    assign in5641_2 = {c2117};
    Full_Adder FA_5641(s5641, c5641, in5641_1, in5641_2, c2115);
    wire[0:0] s5642, in5642_1, in5642_2;
    wire c5642;
    assign in5642_1 = {c2119};
    assign in5642_2 = {c2120};
    Full_Adder FA_5642(s5642, c5642, in5642_1, in5642_2, c2118);
    wire[0:0] s5643, in5643_1, in5643_2;
    wire c5643;
    assign in5643_1 = {c2122};
    assign in5643_2 = {c2123};
    Full_Adder FA_5643(s5643, c5643, in5643_1, in5643_2, c2121);
    wire[0:0] s5644, in5644_1, in5644_2;
    wire c5644;
    assign in5644_1 = {c2125};
    assign in5644_2 = {c2126};
    Full_Adder FA_5644(s5644, c5644, in5644_1, in5644_2, c2124);
    wire[0:0] s5645, in5645_1, in5645_2;
    wire c5645;
    assign in5645_1 = {c2128};
    assign in5645_2 = {c2129};
    Full_Adder FA_5645(s5645, c5645, in5645_1, in5645_2, c2127);
    wire[0:0] s5646, in5646_1, in5646_2;
    wire c5646;
    assign in5646_1 = {c2131};
    assign in5646_2 = {s2132[0]};
    Full_Adder FA_5646(s5646, c5646, in5646_1, in5646_2, c2130);
    wire[0:0] s5647, in5647_1, in5647_2;
    wire c5647;
    assign in5647_1 = {s2134[0]};
    assign in5647_2 = {s2135[0]};
    Full_Adder FA_5647(s5647, c5647, in5647_1, in5647_2, s2133[0]);
    wire[0:0] s5648, in5648_1, in5648_2;
    wire c5648;
    assign in5648_1 = {s2137[0]};
    assign in5648_2 = {s2138[0]};
    Full_Adder FA_5648(s5648, c5648, in5648_1, in5648_2, s2136[0]);
    wire[0:0] s5649, in5649_1, in5649_2;
    wire c5649;
    assign in5649_1 = {s2140[0]};
    assign in5649_2 = {s2141[0]};
    Full_Adder FA_5649(s5649, c5649, in5649_1, in5649_2, s2139[0]);
    wire[0:0] s5650, in5650_1, in5650_2;
    wire c5650;
    assign in5650_1 = {s2143[0]};
    assign in5650_2 = {s2144[0]};
    Full_Adder FA_5650(s5650, c5650, in5650_1, in5650_2, s2142[0]);
    wire[0:0] s5651, in5651_1, in5651_2;
    wire c5651;
    assign in5651_1 = {s2146[0]};
    assign in5651_2 = {s2147[0]};
    Full_Adder FA_5651(s5651, c5651, in5651_1, in5651_2, s2145[0]);
    wire[0:0] s5652, in5652_1, in5652_2;
    wire c5652;
    assign in5652_1 = {s2149[0]};
    assign in5652_2 = {s2150[0]};
    Full_Adder FA_5652(s5652, c5652, in5652_1, in5652_2, s2148[0]);
    wire[0:0] s5653, in5653_1, in5653_2;
    wire c5653;
    assign in5653_1 = {s2152[0]};
    assign in5653_2 = {s2153[0]};
    Full_Adder FA_5653(s5653, c5653, in5653_1, in5653_2, s2151[0]);
    wire[0:0] s5654, in5654_1, in5654_2;
    wire c5654;
    assign in5654_1 = {s2155[0]};
    assign in5654_2 = {s2156[0]};
    Full_Adder FA_5654(s5654, c5654, in5654_1, in5654_2, s2154[0]);
    wire[0:0] s5655, in5655_1, in5655_2;
    wire c5655;
    assign in5655_1 = {pp81[3]};
    assign in5655_2 = {pp82[2]};
    Full_Adder FA_5655(s5655, c5655, in5655_1, in5655_2, pp80[4]);
    wire[0:0] s5656, in5656_1, in5656_2;
    wire c5656;
    assign in5656_1 = {pp84[0]};
    assign in5656_2 = {c2132};
    Full_Adder FA_5656(s5656, c5656, in5656_1, in5656_2, pp83[1]);
    wire[0:0] s5657, in5657_1, in5657_2;
    wire c5657;
    assign in5657_1 = {c2134};
    assign in5657_2 = {c2135};
    Full_Adder FA_5657(s5657, c5657, in5657_1, in5657_2, c2133);
    wire[0:0] s5658, in5658_1, in5658_2;
    wire c5658;
    assign in5658_1 = {c2137};
    assign in5658_2 = {c2138};
    Full_Adder FA_5658(s5658, c5658, in5658_1, in5658_2, c2136);
    wire[0:0] s5659, in5659_1, in5659_2;
    wire c5659;
    assign in5659_1 = {c2140};
    assign in5659_2 = {c2141};
    Full_Adder FA_5659(s5659, c5659, in5659_1, in5659_2, c2139);
    wire[0:0] s5660, in5660_1, in5660_2;
    wire c5660;
    assign in5660_1 = {c2143};
    assign in5660_2 = {c2144};
    Full_Adder FA_5660(s5660, c5660, in5660_1, in5660_2, c2142);
    wire[0:0] s5661, in5661_1, in5661_2;
    wire c5661;
    assign in5661_1 = {c2146};
    assign in5661_2 = {c2147};
    Full_Adder FA_5661(s5661, c5661, in5661_1, in5661_2, c2145);
    wire[0:0] s5662, in5662_1, in5662_2;
    wire c5662;
    assign in5662_1 = {c2149};
    assign in5662_2 = {c2150};
    Full_Adder FA_5662(s5662, c5662, in5662_1, in5662_2, c2148);
    wire[0:0] s5663, in5663_1, in5663_2;
    wire c5663;
    assign in5663_1 = {c2152};
    assign in5663_2 = {c2153};
    Full_Adder FA_5663(s5663, c5663, in5663_1, in5663_2, c2151);
    wire[0:0] s5664, in5664_1, in5664_2;
    wire c5664;
    assign in5664_1 = {c2155};
    assign in5664_2 = {c2156};
    Full_Adder FA_5664(s5664, c5664, in5664_1, in5664_2, c2154);
    wire[0:0] s5665, in5665_1, in5665_2;
    wire c5665;
    assign in5665_1 = {s2158[0]};
    assign in5665_2 = {s2159[0]};
    Full_Adder FA_5665(s5665, c5665, in5665_1, in5665_2, c2157);
    wire[0:0] s5666, in5666_1, in5666_2;
    wire c5666;
    assign in5666_1 = {s2161[0]};
    assign in5666_2 = {s2162[0]};
    Full_Adder FA_5666(s5666, c5666, in5666_1, in5666_2, s2160[0]);
    wire[0:0] s5667, in5667_1, in5667_2;
    wire c5667;
    assign in5667_1 = {s2164[0]};
    assign in5667_2 = {s2165[0]};
    Full_Adder FA_5667(s5667, c5667, in5667_1, in5667_2, s2163[0]);
    wire[0:0] s5668, in5668_1, in5668_2;
    wire c5668;
    assign in5668_1 = {s2167[0]};
    assign in5668_2 = {s2168[0]};
    Full_Adder FA_5668(s5668, c5668, in5668_1, in5668_2, s2166[0]);
    wire[0:0] s5669, in5669_1, in5669_2;
    wire c5669;
    assign in5669_1 = {s2170[0]};
    assign in5669_2 = {s2171[0]};
    Full_Adder FA_5669(s5669, c5669, in5669_1, in5669_2, s2169[0]);
    wire[0:0] s5670, in5670_1, in5670_2;
    wire c5670;
    assign in5670_1 = {s2173[0]};
    assign in5670_2 = {s2174[0]};
    Full_Adder FA_5670(s5670, c5670, in5670_1, in5670_2, s2172[0]);
    wire[0:0] s5671, in5671_1, in5671_2;
    wire c5671;
    assign in5671_1 = {s2176[0]};
    assign in5671_2 = {s2177[0]};
    Full_Adder FA_5671(s5671, c5671, in5671_1, in5671_2, s2175[0]);
    wire[0:0] s5672, in5672_1, in5672_2;
    wire c5672;
    assign in5672_1 = {s2179[0]};
    assign in5672_2 = {s2180[0]};
    Full_Adder FA_5672(s5672, c5672, in5672_1, in5672_2, s2178[0]);
    wire[0:0] s5673, in5673_1, in5673_2;
    wire c5673;
    assign in5673_1 = {s2182[0]};
    assign in5673_2 = {s2183[0]};
    Full_Adder FA_5673(s5673, c5673, in5673_1, in5673_2, s2181[0]);
    wire[0:0] s5674, in5674_1, in5674_2;
    wire c5674;
    assign in5674_1 = {pp84[1]};
    assign in5674_2 = {pp85[0]};
    Full_Adder FA_5674(s5674, c5674, in5674_1, in5674_2, pp83[2]);
    wire[0:0] s5675, in5675_1, in5675_2;
    wire c5675;
    assign in5675_1 = {c2159};
    assign in5675_2 = {c2160};
    Full_Adder FA_5675(s5675, c5675, in5675_1, in5675_2, c2158);
    wire[0:0] s5676, in5676_1, in5676_2;
    wire c5676;
    assign in5676_1 = {c2162};
    assign in5676_2 = {c2163};
    Full_Adder FA_5676(s5676, c5676, in5676_1, in5676_2, c2161);
    wire[0:0] s5677, in5677_1, in5677_2;
    wire c5677;
    assign in5677_1 = {c2165};
    assign in5677_2 = {c2166};
    Full_Adder FA_5677(s5677, c5677, in5677_1, in5677_2, c2164);
    wire[0:0] s5678, in5678_1, in5678_2;
    wire c5678;
    assign in5678_1 = {c2168};
    assign in5678_2 = {c2169};
    Full_Adder FA_5678(s5678, c5678, in5678_1, in5678_2, c2167);
    wire[0:0] s5679, in5679_1, in5679_2;
    wire c5679;
    assign in5679_1 = {c2171};
    assign in5679_2 = {c2172};
    Full_Adder FA_5679(s5679, c5679, in5679_1, in5679_2, c2170);
    wire[0:0] s5680, in5680_1, in5680_2;
    wire c5680;
    assign in5680_1 = {c2174};
    assign in5680_2 = {c2175};
    Full_Adder FA_5680(s5680, c5680, in5680_1, in5680_2, c2173);
    wire[0:0] s5681, in5681_1, in5681_2;
    wire c5681;
    assign in5681_1 = {c2177};
    assign in5681_2 = {c2178};
    Full_Adder FA_5681(s5681, c5681, in5681_1, in5681_2, c2176);
    wire[0:0] s5682, in5682_1, in5682_2;
    wire c5682;
    assign in5682_1 = {c2180};
    assign in5682_2 = {c2181};
    Full_Adder FA_5682(s5682, c5682, in5682_1, in5682_2, c2179);
    wire[0:0] s5683, in5683_1, in5683_2;
    wire c5683;
    assign in5683_1 = {c2183};
    assign in5683_2 = {c2184};
    Full_Adder FA_5683(s5683, c5683, in5683_1, in5683_2, c2182);
    wire[0:0] s5684, in5684_1, in5684_2;
    wire c5684;
    assign in5684_1 = {s2186[0]};
    assign in5684_2 = {s2187[0]};
    Full_Adder FA_5684(s5684, c5684, in5684_1, in5684_2, s2185[0]);
    wire[0:0] s5685, in5685_1, in5685_2;
    wire c5685;
    assign in5685_1 = {s2189[0]};
    assign in5685_2 = {s2190[0]};
    Full_Adder FA_5685(s5685, c5685, in5685_1, in5685_2, s2188[0]);
    wire[0:0] s5686, in5686_1, in5686_2;
    wire c5686;
    assign in5686_1 = {s2192[0]};
    assign in5686_2 = {s2193[0]};
    Full_Adder FA_5686(s5686, c5686, in5686_1, in5686_2, s2191[0]);
    wire[0:0] s5687, in5687_1, in5687_2;
    wire c5687;
    assign in5687_1 = {s2195[0]};
    assign in5687_2 = {s2196[0]};
    Full_Adder FA_5687(s5687, c5687, in5687_1, in5687_2, s2194[0]);
    wire[0:0] s5688, in5688_1, in5688_2;
    wire c5688;
    assign in5688_1 = {s2198[0]};
    assign in5688_2 = {s2199[0]};
    Full_Adder FA_5688(s5688, c5688, in5688_1, in5688_2, s2197[0]);
    wire[0:0] s5689, in5689_1, in5689_2;
    wire c5689;
    assign in5689_1 = {s2201[0]};
    assign in5689_2 = {s2202[0]};
    Full_Adder FA_5689(s5689, c5689, in5689_1, in5689_2, s2200[0]);
    wire[0:0] s5690, in5690_1, in5690_2;
    wire c5690;
    assign in5690_1 = {s2204[0]};
    assign in5690_2 = {s2205[0]};
    Full_Adder FA_5690(s5690, c5690, in5690_1, in5690_2, s2203[0]);
    wire[0:0] s5691, in5691_1, in5691_2;
    wire c5691;
    assign in5691_1 = {s2207[0]};
    assign in5691_2 = {s2208[0]};
    Full_Adder FA_5691(s5691, c5691, in5691_1, in5691_2, s2206[0]);
    wire[0:0] s5692, in5692_1, in5692_2;
    wire c5692;
    assign in5692_1 = {s2210[0]};
    assign in5692_2 = {s2211[0]};
    Full_Adder FA_5692(s5692, c5692, in5692_1, in5692_2, s2209[0]);
    wire[0:0] s5693, in5693_1, in5693_2;
    wire c5693;
    assign in5693_1 = {s1[0]};
    assign in5693_2 = {c2185};
    Full_Adder FA_5693(s5693, c5693, in5693_1, in5693_2, pp86[0]);
    wire[0:0] s5694, in5694_1, in5694_2;
    wire c5694;
    assign in5694_1 = {c2187};
    assign in5694_2 = {c2188};
    Full_Adder FA_5694(s5694, c5694, in5694_1, in5694_2, c2186);
    wire[0:0] s5695, in5695_1, in5695_2;
    wire c5695;
    assign in5695_1 = {c2190};
    assign in5695_2 = {c2191};
    Full_Adder FA_5695(s5695, c5695, in5695_1, in5695_2, c2189);
    wire[0:0] s5696, in5696_1, in5696_2;
    wire c5696;
    assign in5696_1 = {c2193};
    assign in5696_2 = {c2194};
    Full_Adder FA_5696(s5696, c5696, in5696_1, in5696_2, c2192);
    wire[0:0] s5697, in5697_1, in5697_2;
    wire c5697;
    assign in5697_1 = {c2196};
    assign in5697_2 = {c2197};
    Full_Adder FA_5697(s5697, c5697, in5697_1, in5697_2, c2195);
    wire[0:0] s5698, in5698_1, in5698_2;
    wire c5698;
    assign in5698_1 = {c2199};
    assign in5698_2 = {c2200};
    Full_Adder FA_5698(s5698, c5698, in5698_1, in5698_2, c2198);
    wire[0:0] s5699, in5699_1, in5699_2;
    wire c5699;
    assign in5699_1 = {c2202};
    assign in5699_2 = {c2203};
    Full_Adder FA_5699(s5699, c5699, in5699_1, in5699_2, c2201);
    wire[0:0] s5700, in5700_1, in5700_2;
    wire c5700;
    assign in5700_1 = {c2205};
    assign in5700_2 = {c2206};
    Full_Adder FA_5700(s5700, c5700, in5700_1, in5700_2, c2204);
    wire[0:0] s5701, in5701_1, in5701_2;
    wire c5701;
    assign in5701_1 = {c2208};
    assign in5701_2 = {c2209};
    Full_Adder FA_5701(s5701, c5701, in5701_1, in5701_2, c2207);
    wire[0:0] s5702, in5702_1, in5702_2;
    wire c5702;
    assign in5702_1 = {c2211};
    assign in5702_2 = {c2212};
    Full_Adder FA_5702(s5702, c5702, in5702_1, in5702_2, c2210);
    wire[0:0] s5703, in5703_1, in5703_2;
    wire c5703;
    assign in5703_1 = {s2214[0]};
    assign in5703_2 = {s2215[0]};
    Full_Adder FA_5703(s5703, c5703, in5703_1, in5703_2, s2213[0]);
    wire[0:0] s5704, in5704_1, in5704_2;
    wire c5704;
    assign in5704_1 = {s2217[0]};
    assign in5704_2 = {s2218[0]};
    Full_Adder FA_5704(s5704, c5704, in5704_1, in5704_2, s2216[0]);
    wire[0:0] s5705, in5705_1, in5705_2;
    wire c5705;
    assign in5705_1 = {s2220[0]};
    assign in5705_2 = {s2221[0]};
    Full_Adder FA_5705(s5705, c5705, in5705_1, in5705_2, s2219[0]);
    wire[0:0] s5706, in5706_1, in5706_2;
    wire c5706;
    assign in5706_1 = {s2223[0]};
    assign in5706_2 = {s2224[0]};
    Full_Adder FA_5706(s5706, c5706, in5706_1, in5706_2, s2222[0]);
    wire[0:0] s5707, in5707_1, in5707_2;
    wire c5707;
    assign in5707_1 = {s2226[0]};
    assign in5707_2 = {s2227[0]};
    Full_Adder FA_5707(s5707, c5707, in5707_1, in5707_2, s2225[0]);
    wire[0:0] s5708, in5708_1, in5708_2;
    wire c5708;
    assign in5708_1 = {s2229[0]};
    assign in5708_2 = {s2230[0]};
    Full_Adder FA_5708(s5708, c5708, in5708_1, in5708_2, s2228[0]);
    wire[0:0] s5709, in5709_1, in5709_2;
    wire c5709;
    assign in5709_1 = {s2232[0]};
    assign in5709_2 = {s2233[0]};
    Full_Adder FA_5709(s5709, c5709, in5709_1, in5709_2, s2231[0]);
    wire[0:0] s5710, in5710_1, in5710_2;
    wire c5710;
    assign in5710_1 = {s2235[0]};
    assign in5710_2 = {s2236[0]};
    Full_Adder FA_5710(s5710, c5710, in5710_1, in5710_2, s2234[0]);
    wire[0:0] s5711, in5711_1, in5711_2;
    wire c5711;
    assign in5711_1 = {s2238[0]};
    assign in5711_2 = {s2239[0]};
    Full_Adder FA_5711(s5711, c5711, in5711_1, in5711_2, s2237[0]);
    wire[0:0] s5712, in5712_1, in5712_2;
    wire c5712;
    assign in5712_1 = {s3[0]};
    assign in5712_2 = {c2213};
    Full_Adder FA_5712(s5712, c5712, in5712_1, in5712_2, s2[0]);
    wire[0:0] s5713, in5713_1, in5713_2;
    wire c5713;
    assign in5713_1 = {c2215};
    assign in5713_2 = {c2216};
    Full_Adder FA_5713(s5713, c5713, in5713_1, in5713_2, c2214);
    wire[0:0] s5714, in5714_1, in5714_2;
    wire c5714;
    assign in5714_1 = {c2218};
    assign in5714_2 = {c2219};
    Full_Adder FA_5714(s5714, c5714, in5714_1, in5714_2, c2217);
    wire[0:0] s5715, in5715_1, in5715_2;
    wire c5715;
    assign in5715_1 = {c2221};
    assign in5715_2 = {c2222};
    Full_Adder FA_5715(s5715, c5715, in5715_1, in5715_2, c2220);
    wire[0:0] s5716, in5716_1, in5716_2;
    wire c5716;
    assign in5716_1 = {c2224};
    assign in5716_2 = {c2225};
    Full_Adder FA_5716(s5716, c5716, in5716_1, in5716_2, c2223);
    wire[0:0] s5717, in5717_1, in5717_2;
    wire c5717;
    assign in5717_1 = {c2227};
    assign in5717_2 = {c2228};
    Full_Adder FA_5717(s5717, c5717, in5717_1, in5717_2, c2226);
    wire[0:0] s5718, in5718_1, in5718_2;
    wire c5718;
    assign in5718_1 = {c2230};
    assign in5718_2 = {c2231};
    Full_Adder FA_5718(s5718, c5718, in5718_1, in5718_2, c2229);
    wire[0:0] s5719, in5719_1, in5719_2;
    wire c5719;
    assign in5719_1 = {c2233};
    assign in5719_2 = {c2234};
    Full_Adder FA_5719(s5719, c5719, in5719_1, in5719_2, c2232);
    wire[0:0] s5720, in5720_1, in5720_2;
    wire c5720;
    assign in5720_1 = {c2236};
    assign in5720_2 = {c2237};
    Full_Adder FA_5720(s5720, c5720, in5720_1, in5720_2, c2235);
    wire[0:0] s5721, in5721_1, in5721_2;
    wire c5721;
    assign in5721_1 = {c2239};
    assign in5721_2 = {c2240};
    Full_Adder FA_5721(s5721, c5721, in5721_1, in5721_2, c2238);
    wire[0:0] s5722, in5722_1, in5722_2;
    wire c5722;
    assign in5722_1 = {s2242[0]};
    assign in5722_2 = {s2243[0]};
    Full_Adder FA_5722(s5722, c5722, in5722_1, in5722_2, s2241[0]);
    wire[0:0] s5723, in5723_1, in5723_2;
    wire c5723;
    assign in5723_1 = {s2245[0]};
    assign in5723_2 = {s2246[0]};
    Full_Adder FA_5723(s5723, c5723, in5723_1, in5723_2, s2244[0]);
    wire[0:0] s5724, in5724_1, in5724_2;
    wire c5724;
    assign in5724_1 = {s2248[0]};
    assign in5724_2 = {s2249[0]};
    Full_Adder FA_5724(s5724, c5724, in5724_1, in5724_2, s2247[0]);
    wire[0:0] s5725, in5725_1, in5725_2;
    wire c5725;
    assign in5725_1 = {s2251[0]};
    assign in5725_2 = {s2252[0]};
    Full_Adder FA_5725(s5725, c5725, in5725_1, in5725_2, s2250[0]);
    wire[0:0] s5726, in5726_1, in5726_2;
    wire c5726;
    assign in5726_1 = {s2254[0]};
    assign in5726_2 = {s2255[0]};
    Full_Adder FA_5726(s5726, c5726, in5726_1, in5726_2, s2253[0]);
    wire[0:0] s5727, in5727_1, in5727_2;
    wire c5727;
    assign in5727_1 = {s2257[0]};
    assign in5727_2 = {s2258[0]};
    Full_Adder FA_5727(s5727, c5727, in5727_1, in5727_2, s2256[0]);
    wire[0:0] s5728, in5728_1, in5728_2;
    wire c5728;
    assign in5728_1 = {s2260[0]};
    assign in5728_2 = {s2261[0]};
    Full_Adder FA_5728(s5728, c5728, in5728_1, in5728_2, s2259[0]);
    wire[0:0] s5729, in5729_1, in5729_2;
    wire c5729;
    assign in5729_1 = {s2263[0]};
    assign in5729_2 = {s2264[0]};
    Full_Adder FA_5729(s5729, c5729, in5729_1, in5729_2, s2262[0]);
    wire[0:0] s5730, in5730_1, in5730_2;
    wire c5730;
    assign in5730_1 = {s2266[0]};
    assign in5730_2 = {s2267[0]};
    Full_Adder FA_5730(s5730, c5730, in5730_1, in5730_2, s2265[0]);
    wire[0:0] s5731, in5731_1, in5731_2;
    wire c5731;
    assign in5731_1 = {s6[0]};
    assign in5731_2 = {c2241};
    Full_Adder FA_5731(s5731, c5731, in5731_1, in5731_2, s5[0]);
    wire[0:0] s5732, in5732_1, in5732_2;
    wire c5732;
    assign in5732_1 = {c2243};
    assign in5732_2 = {c2244};
    Full_Adder FA_5732(s5732, c5732, in5732_1, in5732_2, c2242);
    wire[0:0] s5733, in5733_1, in5733_2;
    wire c5733;
    assign in5733_1 = {c2246};
    assign in5733_2 = {c2247};
    Full_Adder FA_5733(s5733, c5733, in5733_1, in5733_2, c2245);
    wire[0:0] s5734, in5734_1, in5734_2;
    wire c5734;
    assign in5734_1 = {c2249};
    assign in5734_2 = {c2250};
    Full_Adder FA_5734(s5734, c5734, in5734_1, in5734_2, c2248);
    wire[0:0] s5735, in5735_1, in5735_2;
    wire c5735;
    assign in5735_1 = {c2252};
    assign in5735_2 = {c2253};
    Full_Adder FA_5735(s5735, c5735, in5735_1, in5735_2, c2251);
    wire[0:0] s5736, in5736_1, in5736_2;
    wire c5736;
    assign in5736_1 = {c2255};
    assign in5736_2 = {c2256};
    Full_Adder FA_5736(s5736, c5736, in5736_1, in5736_2, c2254);
    wire[0:0] s5737, in5737_1, in5737_2;
    wire c5737;
    assign in5737_1 = {c2258};
    assign in5737_2 = {c2259};
    Full_Adder FA_5737(s5737, c5737, in5737_1, in5737_2, c2257);
    wire[0:0] s5738, in5738_1, in5738_2;
    wire c5738;
    assign in5738_1 = {c2261};
    assign in5738_2 = {c2262};
    Full_Adder FA_5738(s5738, c5738, in5738_1, in5738_2, c2260);
    wire[0:0] s5739, in5739_1, in5739_2;
    wire c5739;
    assign in5739_1 = {c2264};
    assign in5739_2 = {c2265};
    Full_Adder FA_5739(s5739, c5739, in5739_1, in5739_2, c2263);
    wire[0:0] s5740, in5740_1, in5740_2;
    wire c5740;
    assign in5740_1 = {c2267};
    assign in5740_2 = {c2268};
    Full_Adder FA_5740(s5740, c5740, in5740_1, in5740_2, c2266);
    wire[0:0] s5741, in5741_1, in5741_2;
    wire c5741;
    assign in5741_1 = {s2270[0]};
    assign in5741_2 = {s2271[0]};
    Full_Adder FA_5741(s5741, c5741, in5741_1, in5741_2, s2269[0]);
    wire[0:0] s5742, in5742_1, in5742_2;
    wire c5742;
    assign in5742_1 = {s2273[0]};
    assign in5742_2 = {s2274[0]};
    Full_Adder FA_5742(s5742, c5742, in5742_1, in5742_2, s2272[0]);
    wire[0:0] s5743, in5743_1, in5743_2;
    wire c5743;
    assign in5743_1 = {s2276[0]};
    assign in5743_2 = {s2277[0]};
    Full_Adder FA_5743(s5743, c5743, in5743_1, in5743_2, s2275[0]);
    wire[0:0] s5744, in5744_1, in5744_2;
    wire c5744;
    assign in5744_1 = {s2279[0]};
    assign in5744_2 = {s2280[0]};
    Full_Adder FA_5744(s5744, c5744, in5744_1, in5744_2, s2278[0]);
    wire[0:0] s5745, in5745_1, in5745_2;
    wire c5745;
    assign in5745_1 = {s2282[0]};
    assign in5745_2 = {s2283[0]};
    Full_Adder FA_5745(s5745, c5745, in5745_1, in5745_2, s2281[0]);
    wire[0:0] s5746, in5746_1, in5746_2;
    wire c5746;
    assign in5746_1 = {s2285[0]};
    assign in5746_2 = {s2286[0]};
    Full_Adder FA_5746(s5746, c5746, in5746_1, in5746_2, s2284[0]);
    wire[0:0] s5747, in5747_1, in5747_2;
    wire c5747;
    assign in5747_1 = {s2288[0]};
    assign in5747_2 = {s2289[0]};
    Full_Adder FA_5747(s5747, c5747, in5747_1, in5747_2, s2287[0]);
    wire[0:0] s5748, in5748_1, in5748_2;
    wire c5748;
    assign in5748_1 = {s2291[0]};
    assign in5748_2 = {s2292[0]};
    Full_Adder FA_5748(s5748, c5748, in5748_1, in5748_2, s2290[0]);
    wire[0:0] s5749, in5749_1, in5749_2;
    wire c5749;
    assign in5749_1 = {s2294[0]};
    assign in5749_2 = {s2295[0]};
    Full_Adder FA_5749(s5749, c5749, in5749_1, in5749_2, s2293[0]);
    wire[0:0] s5750, in5750_1, in5750_2;
    wire c5750;
    assign in5750_1 = {s10[0]};
    assign in5750_2 = {c2269};
    Full_Adder FA_5750(s5750, c5750, in5750_1, in5750_2, s9[0]);
    wire[0:0] s5751, in5751_1, in5751_2;
    wire c5751;
    assign in5751_1 = {c2271};
    assign in5751_2 = {c2272};
    Full_Adder FA_5751(s5751, c5751, in5751_1, in5751_2, c2270);
    wire[0:0] s5752, in5752_1, in5752_2;
    wire c5752;
    assign in5752_1 = {c2274};
    assign in5752_2 = {c2275};
    Full_Adder FA_5752(s5752, c5752, in5752_1, in5752_2, c2273);
    wire[0:0] s5753, in5753_1, in5753_2;
    wire c5753;
    assign in5753_1 = {c2277};
    assign in5753_2 = {c2278};
    Full_Adder FA_5753(s5753, c5753, in5753_1, in5753_2, c2276);
    wire[0:0] s5754, in5754_1, in5754_2;
    wire c5754;
    assign in5754_1 = {c2280};
    assign in5754_2 = {c2281};
    Full_Adder FA_5754(s5754, c5754, in5754_1, in5754_2, c2279);
    wire[0:0] s5755, in5755_1, in5755_2;
    wire c5755;
    assign in5755_1 = {c2283};
    assign in5755_2 = {c2284};
    Full_Adder FA_5755(s5755, c5755, in5755_1, in5755_2, c2282);
    wire[0:0] s5756, in5756_1, in5756_2;
    wire c5756;
    assign in5756_1 = {c2286};
    assign in5756_2 = {c2287};
    Full_Adder FA_5756(s5756, c5756, in5756_1, in5756_2, c2285);
    wire[0:0] s5757, in5757_1, in5757_2;
    wire c5757;
    assign in5757_1 = {c2289};
    assign in5757_2 = {c2290};
    Full_Adder FA_5757(s5757, c5757, in5757_1, in5757_2, c2288);
    wire[0:0] s5758, in5758_1, in5758_2;
    wire c5758;
    assign in5758_1 = {c2292};
    assign in5758_2 = {c2293};
    Full_Adder FA_5758(s5758, c5758, in5758_1, in5758_2, c2291);
    wire[0:0] s5759, in5759_1, in5759_2;
    wire c5759;
    assign in5759_1 = {c2295};
    assign in5759_2 = {c2296};
    Full_Adder FA_5759(s5759, c5759, in5759_1, in5759_2, c2294);
    wire[0:0] s5760, in5760_1, in5760_2;
    wire c5760;
    assign in5760_1 = {s2298[0]};
    assign in5760_2 = {s2299[0]};
    Full_Adder FA_5760(s5760, c5760, in5760_1, in5760_2, s2297[0]);
    wire[0:0] s5761, in5761_1, in5761_2;
    wire c5761;
    assign in5761_1 = {s2301[0]};
    assign in5761_2 = {s2302[0]};
    Full_Adder FA_5761(s5761, c5761, in5761_1, in5761_2, s2300[0]);
    wire[0:0] s5762, in5762_1, in5762_2;
    wire c5762;
    assign in5762_1 = {s2304[0]};
    assign in5762_2 = {s2305[0]};
    Full_Adder FA_5762(s5762, c5762, in5762_1, in5762_2, s2303[0]);
    wire[0:0] s5763, in5763_1, in5763_2;
    wire c5763;
    assign in5763_1 = {s2307[0]};
    assign in5763_2 = {s2308[0]};
    Full_Adder FA_5763(s5763, c5763, in5763_1, in5763_2, s2306[0]);
    wire[0:0] s5764, in5764_1, in5764_2;
    wire c5764;
    assign in5764_1 = {s2310[0]};
    assign in5764_2 = {s2311[0]};
    Full_Adder FA_5764(s5764, c5764, in5764_1, in5764_2, s2309[0]);
    wire[0:0] s5765, in5765_1, in5765_2;
    wire c5765;
    assign in5765_1 = {s2313[0]};
    assign in5765_2 = {s2314[0]};
    Full_Adder FA_5765(s5765, c5765, in5765_1, in5765_2, s2312[0]);
    wire[0:0] s5766, in5766_1, in5766_2;
    wire c5766;
    assign in5766_1 = {s2316[0]};
    assign in5766_2 = {s2317[0]};
    Full_Adder FA_5766(s5766, c5766, in5766_1, in5766_2, s2315[0]);
    wire[0:0] s5767, in5767_1, in5767_2;
    wire c5767;
    assign in5767_1 = {s2319[0]};
    assign in5767_2 = {s2320[0]};
    Full_Adder FA_5767(s5767, c5767, in5767_1, in5767_2, s2318[0]);
    wire[0:0] s5768, in5768_1, in5768_2;
    wire c5768;
    assign in5768_1 = {s2322[0]};
    assign in5768_2 = {s2323[0]};
    Full_Adder FA_5768(s5768, c5768, in5768_1, in5768_2, s2321[0]);
    wire[0:0] s5769, in5769_1, in5769_2;
    wire c5769;
    assign in5769_1 = {s15[0]};
    assign in5769_2 = {c2297};
    Full_Adder FA_5769(s5769, c5769, in5769_1, in5769_2, s14[0]);
    wire[0:0] s5770, in5770_1, in5770_2;
    wire c5770;
    assign in5770_1 = {c2299};
    assign in5770_2 = {c2300};
    Full_Adder FA_5770(s5770, c5770, in5770_1, in5770_2, c2298);
    wire[0:0] s5771, in5771_1, in5771_2;
    wire c5771;
    assign in5771_1 = {c2302};
    assign in5771_2 = {c2303};
    Full_Adder FA_5771(s5771, c5771, in5771_1, in5771_2, c2301);
    wire[0:0] s5772, in5772_1, in5772_2;
    wire c5772;
    assign in5772_1 = {c2305};
    assign in5772_2 = {c2306};
    Full_Adder FA_5772(s5772, c5772, in5772_1, in5772_2, c2304);
    wire[0:0] s5773, in5773_1, in5773_2;
    wire c5773;
    assign in5773_1 = {c2308};
    assign in5773_2 = {c2309};
    Full_Adder FA_5773(s5773, c5773, in5773_1, in5773_2, c2307);
    wire[0:0] s5774, in5774_1, in5774_2;
    wire c5774;
    assign in5774_1 = {c2311};
    assign in5774_2 = {c2312};
    Full_Adder FA_5774(s5774, c5774, in5774_1, in5774_2, c2310);
    wire[0:0] s5775, in5775_1, in5775_2;
    wire c5775;
    assign in5775_1 = {c2314};
    assign in5775_2 = {c2315};
    Full_Adder FA_5775(s5775, c5775, in5775_1, in5775_2, c2313);
    wire[0:0] s5776, in5776_1, in5776_2;
    wire c5776;
    assign in5776_1 = {c2317};
    assign in5776_2 = {c2318};
    Full_Adder FA_5776(s5776, c5776, in5776_1, in5776_2, c2316);
    wire[0:0] s5777, in5777_1, in5777_2;
    wire c5777;
    assign in5777_1 = {c2320};
    assign in5777_2 = {c2321};
    Full_Adder FA_5777(s5777, c5777, in5777_1, in5777_2, c2319);
    wire[0:0] s5778, in5778_1, in5778_2;
    wire c5778;
    assign in5778_1 = {c2323};
    assign in5778_2 = {c2324};
    Full_Adder FA_5778(s5778, c5778, in5778_1, in5778_2, c2322);
    wire[0:0] s5779, in5779_1, in5779_2;
    wire c5779;
    assign in5779_1 = {s2326[0]};
    assign in5779_2 = {s2327[0]};
    Full_Adder FA_5779(s5779, c5779, in5779_1, in5779_2, s2325[0]);
    wire[0:0] s5780, in5780_1, in5780_2;
    wire c5780;
    assign in5780_1 = {s2329[0]};
    assign in5780_2 = {s2330[0]};
    Full_Adder FA_5780(s5780, c5780, in5780_1, in5780_2, s2328[0]);
    wire[0:0] s5781, in5781_1, in5781_2;
    wire c5781;
    assign in5781_1 = {s2332[0]};
    assign in5781_2 = {s2333[0]};
    Full_Adder FA_5781(s5781, c5781, in5781_1, in5781_2, s2331[0]);
    wire[0:0] s5782, in5782_1, in5782_2;
    wire c5782;
    assign in5782_1 = {s2335[0]};
    assign in5782_2 = {s2336[0]};
    Full_Adder FA_5782(s5782, c5782, in5782_1, in5782_2, s2334[0]);
    wire[0:0] s5783, in5783_1, in5783_2;
    wire c5783;
    assign in5783_1 = {s2338[0]};
    assign in5783_2 = {s2339[0]};
    Full_Adder FA_5783(s5783, c5783, in5783_1, in5783_2, s2337[0]);
    wire[0:0] s5784, in5784_1, in5784_2;
    wire c5784;
    assign in5784_1 = {s2341[0]};
    assign in5784_2 = {s2342[0]};
    Full_Adder FA_5784(s5784, c5784, in5784_1, in5784_2, s2340[0]);
    wire[0:0] s5785, in5785_1, in5785_2;
    wire c5785;
    assign in5785_1 = {s2344[0]};
    assign in5785_2 = {s2345[0]};
    Full_Adder FA_5785(s5785, c5785, in5785_1, in5785_2, s2343[0]);
    wire[0:0] s5786, in5786_1, in5786_2;
    wire c5786;
    assign in5786_1 = {s2347[0]};
    assign in5786_2 = {s2348[0]};
    Full_Adder FA_5786(s5786, c5786, in5786_1, in5786_2, s2346[0]);
    wire[0:0] s5787, in5787_1, in5787_2;
    wire c5787;
    assign in5787_1 = {s2350[0]};
    assign in5787_2 = {s2351[0]};
    Full_Adder FA_5787(s5787, c5787, in5787_1, in5787_2, s2349[0]);
    wire[0:0] s5788, in5788_1, in5788_2;
    wire c5788;
    assign in5788_1 = {s21[0]};
    assign in5788_2 = {c2325};
    Full_Adder FA_5788(s5788, c5788, in5788_1, in5788_2, s20[0]);
    wire[0:0] s5789, in5789_1, in5789_2;
    wire c5789;
    assign in5789_1 = {c2327};
    assign in5789_2 = {c2328};
    Full_Adder FA_5789(s5789, c5789, in5789_1, in5789_2, c2326);
    wire[0:0] s5790, in5790_1, in5790_2;
    wire c5790;
    assign in5790_1 = {c2330};
    assign in5790_2 = {c2331};
    Full_Adder FA_5790(s5790, c5790, in5790_1, in5790_2, c2329);
    wire[0:0] s5791, in5791_1, in5791_2;
    wire c5791;
    assign in5791_1 = {c2333};
    assign in5791_2 = {c2334};
    Full_Adder FA_5791(s5791, c5791, in5791_1, in5791_2, c2332);
    wire[0:0] s5792, in5792_1, in5792_2;
    wire c5792;
    assign in5792_1 = {c2336};
    assign in5792_2 = {c2337};
    Full_Adder FA_5792(s5792, c5792, in5792_1, in5792_2, c2335);
    wire[0:0] s5793, in5793_1, in5793_2;
    wire c5793;
    assign in5793_1 = {c2339};
    assign in5793_2 = {c2340};
    Full_Adder FA_5793(s5793, c5793, in5793_1, in5793_2, c2338);
    wire[0:0] s5794, in5794_1, in5794_2;
    wire c5794;
    assign in5794_1 = {c2342};
    assign in5794_2 = {c2343};
    Full_Adder FA_5794(s5794, c5794, in5794_1, in5794_2, c2341);
    wire[0:0] s5795, in5795_1, in5795_2;
    wire c5795;
    assign in5795_1 = {c2345};
    assign in5795_2 = {c2346};
    Full_Adder FA_5795(s5795, c5795, in5795_1, in5795_2, c2344);
    wire[0:0] s5796, in5796_1, in5796_2;
    wire c5796;
    assign in5796_1 = {c2348};
    assign in5796_2 = {c2349};
    Full_Adder FA_5796(s5796, c5796, in5796_1, in5796_2, c2347);
    wire[0:0] s5797, in5797_1, in5797_2;
    wire c5797;
    assign in5797_1 = {c2351};
    assign in5797_2 = {c2352};
    Full_Adder FA_5797(s5797, c5797, in5797_1, in5797_2, c2350);
    wire[0:0] s5798, in5798_1, in5798_2;
    wire c5798;
    assign in5798_1 = {s2354[0]};
    assign in5798_2 = {s2355[0]};
    Full_Adder FA_5798(s5798, c5798, in5798_1, in5798_2, s2353[0]);
    wire[0:0] s5799, in5799_1, in5799_2;
    wire c5799;
    assign in5799_1 = {s2357[0]};
    assign in5799_2 = {s2358[0]};
    Full_Adder FA_5799(s5799, c5799, in5799_1, in5799_2, s2356[0]);
    wire[0:0] s5800, in5800_1, in5800_2;
    wire c5800;
    assign in5800_1 = {s2360[0]};
    assign in5800_2 = {s2361[0]};
    Full_Adder FA_5800(s5800, c5800, in5800_1, in5800_2, s2359[0]);
    wire[0:0] s5801, in5801_1, in5801_2;
    wire c5801;
    assign in5801_1 = {s2363[0]};
    assign in5801_2 = {s2364[0]};
    Full_Adder FA_5801(s5801, c5801, in5801_1, in5801_2, s2362[0]);
    wire[0:0] s5802, in5802_1, in5802_2;
    wire c5802;
    assign in5802_1 = {s2366[0]};
    assign in5802_2 = {s2367[0]};
    Full_Adder FA_5802(s5802, c5802, in5802_1, in5802_2, s2365[0]);
    wire[0:0] s5803, in5803_1, in5803_2;
    wire c5803;
    assign in5803_1 = {s2369[0]};
    assign in5803_2 = {s2370[0]};
    Full_Adder FA_5803(s5803, c5803, in5803_1, in5803_2, s2368[0]);
    wire[0:0] s5804, in5804_1, in5804_2;
    wire c5804;
    assign in5804_1 = {s2372[0]};
    assign in5804_2 = {s2373[0]};
    Full_Adder FA_5804(s5804, c5804, in5804_1, in5804_2, s2371[0]);
    wire[0:0] s5805, in5805_1, in5805_2;
    wire c5805;
    assign in5805_1 = {s2375[0]};
    assign in5805_2 = {s2376[0]};
    Full_Adder FA_5805(s5805, c5805, in5805_1, in5805_2, s2374[0]);
    wire[0:0] s5806, in5806_1, in5806_2;
    wire c5806;
    assign in5806_1 = {s2378[0]};
    assign in5806_2 = {s2379[0]};
    Full_Adder FA_5806(s5806, c5806, in5806_1, in5806_2, s2377[0]);
    wire[0:0] s5807, in5807_1, in5807_2;
    wire c5807;
    assign in5807_1 = {s28[0]};
    assign in5807_2 = {c2353};
    Full_Adder FA_5807(s5807, c5807, in5807_1, in5807_2, s27[0]);
    wire[0:0] s5808, in5808_1, in5808_2;
    wire c5808;
    assign in5808_1 = {c2355};
    assign in5808_2 = {c2356};
    Full_Adder FA_5808(s5808, c5808, in5808_1, in5808_2, c2354);
    wire[0:0] s5809, in5809_1, in5809_2;
    wire c5809;
    assign in5809_1 = {c2358};
    assign in5809_2 = {c2359};
    Full_Adder FA_5809(s5809, c5809, in5809_1, in5809_2, c2357);
    wire[0:0] s5810, in5810_1, in5810_2;
    wire c5810;
    assign in5810_1 = {c2361};
    assign in5810_2 = {c2362};
    Full_Adder FA_5810(s5810, c5810, in5810_1, in5810_2, c2360);
    wire[0:0] s5811, in5811_1, in5811_2;
    wire c5811;
    assign in5811_1 = {c2364};
    assign in5811_2 = {c2365};
    Full_Adder FA_5811(s5811, c5811, in5811_1, in5811_2, c2363);
    wire[0:0] s5812, in5812_1, in5812_2;
    wire c5812;
    assign in5812_1 = {c2367};
    assign in5812_2 = {c2368};
    Full_Adder FA_5812(s5812, c5812, in5812_1, in5812_2, c2366);
    wire[0:0] s5813, in5813_1, in5813_2;
    wire c5813;
    assign in5813_1 = {c2370};
    assign in5813_2 = {c2371};
    Full_Adder FA_5813(s5813, c5813, in5813_1, in5813_2, c2369);
    wire[0:0] s5814, in5814_1, in5814_2;
    wire c5814;
    assign in5814_1 = {c2373};
    assign in5814_2 = {c2374};
    Full_Adder FA_5814(s5814, c5814, in5814_1, in5814_2, c2372);
    wire[0:0] s5815, in5815_1, in5815_2;
    wire c5815;
    assign in5815_1 = {c2376};
    assign in5815_2 = {c2377};
    Full_Adder FA_5815(s5815, c5815, in5815_1, in5815_2, c2375);
    wire[0:0] s5816, in5816_1, in5816_2;
    wire c5816;
    assign in5816_1 = {c2379};
    assign in5816_2 = {c2380};
    Full_Adder FA_5816(s5816, c5816, in5816_1, in5816_2, c2378);
    wire[0:0] s5817, in5817_1, in5817_2;
    wire c5817;
    assign in5817_1 = {s2382[0]};
    assign in5817_2 = {s2383[0]};
    Full_Adder FA_5817(s5817, c5817, in5817_1, in5817_2, s2381[0]);
    wire[0:0] s5818, in5818_1, in5818_2;
    wire c5818;
    assign in5818_1 = {s2385[0]};
    assign in5818_2 = {s2386[0]};
    Full_Adder FA_5818(s5818, c5818, in5818_1, in5818_2, s2384[0]);
    wire[0:0] s5819, in5819_1, in5819_2;
    wire c5819;
    assign in5819_1 = {s2388[0]};
    assign in5819_2 = {s2389[0]};
    Full_Adder FA_5819(s5819, c5819, in5819_1, in5819_2, s2387[0]);
    wire[0:0] s5820, in5820_1, in5820_2;
    wire c5820;
    assign in5820_1 = {s2391[0]};
    assign in5820_2 = {s2392[0]};
    Full_Adder FA_5820(s5820, c5820, in5820_1, in5820_2, s2390[0]);
    wire[0:0] s5821, in5821_1, in5821_2;
    wire c5821;
    assign in5821_1 = {s2394[0]};
    assign in5821_2 = {s2395[0]};
    Full_Adder FA_5821(s5821, c5821, in5821_1, in5821_2, s2393[0]);
    wire[0:0] s5822, in5822_1, in5822_2;
    wire c5822;
    assign in5822_1 = {s2397[0]};
    assign in5822_2 = {s2398[0]};
    Full_Adder FA_5822(s5822, c5822, in5822_1, in5822_2, s2396[0]);
    wire[0:0] s5823, in5823_1, in5823_2;
    wire c5823;
    assign in5823_1 = {s2400[0]};
    assign in5823_2 = {s2401[0]};
    Full_Adder FA_5823(s5823, c5823, in5823_1, in5823_2, s2399[0]);
    wire[0:0] s5824, in5824_1, in5824_2;
    wire c5824;
    assign in5824_1 = {s2403[0]};
    assign in5824_2 = {s2404[0]};
    Full_Adder FA_5824(s5824, c5824, in5824_1, in5824_2, s2402[0]);
    wire[0:0] s5825, in5825_1, in5825_2;
    wire c5825;
    assign in5825_1 = {s2406[0]};
    assign in5825_2 = {s2407[0]};
    Full_Adder FA_5825(s5825, c5825, in5825_1, in5825_2, s2405[0]);
    wire[0:0] s5826, in5826_1, in5826_2;
    wire c5826;
    assign in5826_1 = {s36[0]};
    assign in5826_2 = {c2381};
    Full_Adder FA_5826(s5826, c5826, in5826_1, in5826_2, s35[0]);
    wire[0:0] s5827, in5827_1, in5827_2;
    wire c5827;
    assign in5827_1 = {c2383};
    assign in5827_2 = {c2384};
    Full_Adder FA_5827(s5827, c5827, in5827_1, in5827_2, c2382);
    wire[0:0] s5828, in5828_1, in5828_2;
    wire c5828;
    assign in5828_1 = {c2386};
    assign in5828_2 = {c2387};
    Full_Adder FA_5828(s5828, c5828, in5828_1, in5828_2, c2385);
    wire[0:0] s5829, in5829_1, in5829_2;
    wire c5829;
    assign in5829_1 = {c2389};
    assign in5829_2 = {c2390};
    Full_Adder FA_5829(s5829, c5829, in5829_1, in5829_2, c2388);
    wire[0:0] s5830, in5830_1, in5830_2;
    wire c5830;
    assign in5830_1 = {c2392};
    assign in5830_2 = {c2393};
    Full_Adder FA_5830(s5830, c5830, in5830_1, in5830_2, c2391);
    wire[0:0] s5831, in5831_1, in5831_2;
    wire c5831;
    assign in5831_1 = {c2395};
    assign in5831_2 = {c2396};
    Full_Adder FA_5831(s5831, c5831, in5831_1, in5831_2, c2394);
    wire[0:0] s5832, in5832_1, in5832_2;
    wire c5832;
    assign in5832_1 = {c2398};
    assign in5832_2 = {c2399};
    Full_Adder FA_5832(s5832, c5832, in5832_1, in5832_2, c2397);
    wire[0:0] s5833, in5833_1, in5833_2;
    wire c5833;
    assign in5833_1 = {c2401};
    assign in5833_2 = {c2402};
    Full_Adder FA_5833(s5833, c5833, in5833_1, in5833_2, c2400);
    wire[0:0] s5834, in5834_1, in5834_2;
    wire c5834;
    assign in5834_1 = {c2404};
    assign in5834_2 = {c2405};
    Full_Adder FA_5834(s5834, c5834, in5834_1, in5834_2, c2403);
    wire[0:0] s5835, in5835_1, in5835_2;
    wire c5835;
    assign in5835_1 = {c2407};
    assign in5835_2 = {c2408};
    Full_Adder FA_5835(s5835, c5835, in5835_1, in5835_2, c2406);
    wire[0:0] s5836, in5836_1, in5836_2;
    wire c5836;
    assign in5836_1 = {s2410[0]};
    assign in5836_2 = {s2411[0]};
    Full_Adder FA_5836(s5836, c5836, in5836_1, in5836_2, s2409[0]);
    wire[0:0] s5837, in5837_1, in5837_2;
    wire c5837;
    assign in5837_1 = {s2413[0]};
    assign in5837_2 = {s2414[0]};
    Full_Adder FA_5837(s5837, c5837, in5837_1, in5837_2, s2412[0]);
    wire[0:0] s5838, in5838_1, in5838_2;
    wire c5838;
    assign in5838_1 = {s2416[0]};
    assign in5838_2 = {s2417[0]};
    Full_Adder FA_5838(s5838, c5838, in5838_1, in5838_2, s2415[0]);
    wire[0:0] s5839, in5839_1, in5839_2;
    wire c5839;
    assign in5839_1 = {s2419[0]};
    assign in5839_2 = {s2420[0]};
    Full_Adder FA_5839(s5839, c5839, in5839_1, in5839_2, s2418[0]);
    wire[0:0] s5840, in5840_1, in5840_2;
    wire c5840;
    assign in5840_1 = {s2422[0]};
    assign in5840_2 = {s2423[0]};
    Full_Adder FA_5840(s5840, c5840, in5840_1, in5840_2, s2421[0]);
    wire[0:0] s5841, in5841_1, in5841_2;
    wire c5841;
    assign in5841_1 = {s2425[0]};
    assign in5841_2 = {s2426[0]};
    Full_Adder FA_5841(s5841, c5841, in5841_1, in5841_2, s2424[0]);
    wire[0:0] s5842, in5842_1, in5842_2;
    wire c5842;
    assign in5842_1 = {s2428[0]};
    assign in5842_2 = {s2429[0]};
    Full_Adder FA_5842(s5842, c5842, in5842_1, in5842_2, s2427[0]);
    wire[0:0] s5843, in5843_1, in5843_2;
    wire c5843;
    assign in5843_1 = {s2431[0]};
    assign in5843_2 = {s2432[0]};
    Full_Adder FA_5843(s5843, c5843, in5843_1, in5843_2, s2430[0]);
    wire[0:0] s5844, in5844_1, in5844_2;
    wire c5844;
    assign in5844_1 = {s2434[0]};
    assign in5844_2 = {s2435[0]};
    Full_Adder FA_5844(s5844, c5844, in5844_1, in5844_2, s2433[0]);
    wire[0:0] s5845, in5845_1, in5845_2;
    wire c5845;
    assign in5845_1 = {s45[0]};
    assign in5845_2 = {c2409};
    Full_Adder FA_5845(s5845, c5845, in5845_1, in5845_2, s44[0]);
    wire[0:0] s5846, in5846_1, in5846_2;
    wire c5846;
    assign in5846_1 = {c2411};
    assign in5846_2 = {c2412};
    Full_Adder FA_5846(s5846, c5846, in5846_1, in5846_2, c2410);
    wire[0:0] s5847, in5847_1, in5847_2;
    wire c5847;
    assign in5847_1 = {c2414};
    assign in5847_2 = {c2415};
    Full_Adder FA_5847(s5847, c5847, in5847_1, in5847_2, c2413);
    wire[0:0] s5848, in5848_1, in5848_2;
    wire c5848;
    assign in5848_1 = {c2417};
    assign in5848_2 = {c2418};
    Full_Adder FA_5848(s5848, c5848, in5848_1, in5848_2, c2416);
    wire[0:0] s5849, in5849_1, in5849_2;
    wire c5849;
    assign in5849_1 = {c2420};
    assign in5849_2 = {c2421};
    Full_Adder FA_5849(s5849, c5849, in5849_1, in5849_2, c2419);
    wire[0:0] s5850, in5850_1, in5850_2;
    wire c5850;
    assign in5850_1 = {c2423};
    assign in5850_2 = {c2424};
    Full_Adder FA_5850(s5850, c5850, in5850_1, in5850_2, c2422);
    wire[0:0] s5851, in5851_1, in5851_2;
    wire c5851;
    assign in5851_1 = {c2426};
    assign in5851_2 = {c2427};
    Full_Adder FA_5851(s5851, c5851, in5851_1, in5851_2, c2425);
    wire[0:0] s5852, in5852_1, in5852_2;
    wire c5852;
    assign in5852_1 = {c2429};
    assign in5852_2 = {c2430};
    Full_Adder FA_5852(s5852, c5852, in5852_1, in5852_2, c2428);
    wire[0:0] s5853, in5853_1, in5853_2;
    wire c5853;
    assign in5853_1 = {c2432};
    assign in5853_2 = {c2433};
    Full_Adder FA_5853(s5853, c5853, in5853_1, in5853_2, c2431);
    wire[0:0] s5854, in5854_1, in5854_2;
    wire c5854;
    assign in5854_1 = {c2435};
    assign in5854_2 = {c2436};
    Full_Adder FA_5854(s5854, c5854, in5854_1, in5854_2, c2434);
    wire[0:0] s5855, in5855_1, in5855_2;
    wire c5855;
    assign in5855_1 = {s2438[0]};
    assign in5855_2 = {s2439[0]};
    Full_Adder FA_5855(s5855, c5855, in5855_1, in5855_2, s2437[0]);
    wire[0:0] s5856, in5856_1, in5856_2;
    wire c5856;
    assign in5856_1 = {s2441[0]};
    assign in5856_2 = {s2442[0]};
    Full_Adder FA_5856(s5856, c5856, in5856_1, in5856_2, s2440[0]);
    wire[0:0] s5857, in5857_1, in5857_2;
    wire c5857;
    assign in5857_1 = {s2444[0]};
    assign in5857_2 = {s2445[0]};
    Full_Adder FA_5857(s5857, c5857, in5857_1, in5857_2, s2443[0]);
    wire[0:0] s5858, in5858_1, in5858_2;
    wire c5858;
    assign in5858_1 = {s2447[0]};
    assign in5858_2 = {s2448[0]};
    Full_Adder FA_5858(s5858, c5858, in5858_1, in5858_2, s2446[0]);
    wire[0:0] s5859, in5859_1, in5859_2;
    wire c5859;
    assign in5859_1 = {s2450[0]};
    assign in5859_2 = {s2451[0]};
    Full_Adder FA_5859(s5859, c5859, in5859_1, in5859_2, s2449[0]);
    wire[0:0] s5860, in5860_1, in5860_2;
    wire c5860;
    assign in5860_1 = {s2453[0]};
    assign in5860_2 = {s2454[0]};
    Full_Adder FA_5860(s5860, c5860, in5860_1, in5860_2, s2452[0]);
    wire[0:0] s5861, in5861_1, in5861_2;
    wire c5861;
    assign in5861_1 = {s2456[0]};
    assign in5861_2 = {s2457[0]};
    Full_Adder FA_5861(s5861, c5861, in5861_1, in5861_2, s2455[0]);
    wire[0:0] s5862, in5862_1, in5862_2;
    wire c5862;
    assign in5862_1 = {s2459[0]};
    assign in5862_2 = {s2460[0]};
    Full_Adder FA_5862(s5862, c5862, in5862_1, in5862_2, s2458[0]);
    wire[0:0] s5863, in5863_1, in5863_2;
    wire c5863;
    assign in5863_1 = {s2462[0]};
    assign in5863_2 = {s2463[0]};
    Full_Adder FA_5863(s5863, c5863, in5863_1, in5863_2, s2461[0]);
    wire[0:0] s5864, in5864_1, in5864_2;
    wire c5864;
    assign in5864_1 = {s55[0]};
    assign in5864_2 = {c2437};
    Full_Adder FA_5864(s5864, c5864, in5864_1, in5864_2, s54[0]);
    wire[0:0] s5865, in5865_1, in5865_2;
    wire c5865;
    assign in5865_1 = {c2439};
    assign in5865_2 = {c2440};
    Full_Adder FA_5865(s5865, c5865, in5865_1, in5865_2, c2438);
    wire[0:0] s5866, in5866_1, in5866_2;
    wire c5866;
    assign in5866_1 = {c2442};
    assign in5866_2 = {c2443};
    Full_Adder FA_5866(s5866, c5866, in5866_1, in5866_2, c2441);
    wire[0:0] s5867, in5867_1, in5867_2;
    wire c5867;
    assign in5867_1 = {c2445};
    assign in5867_2 = {c2446};
    Full_Adder FA_5867(s5867, c5867, in5867_1, in5867_2, c2444);
    wire[0:0] s5868, in5868_1, in5868_2;
    wire c5868;
    assign in5868_1 = {c2448};
    assign in5868_2 = {c2449};
    Full_Adder FA_5868(s5868, c5868, in5868_1, in5868_2, c2447);
    wire[0:0] s5869, in5869_1, in5869_2;
    wire c5869;
    assign in5869_1 = {c2451};
    assign in5869_2 = {c2452};
    Full_Adder FA_5869(s5869, c5869, in5869_1, in5869_2, c2450);
    wire[0:0] s5870, in5870_1, in5870_2;
    wire c5870;
    assign in5870_1 = {c2454};
    assign in5870_2 = {c2455};
    Full_Adder FA_5870(s5870, c5870, in5870_1, in5870_2, c2453);
    wire[0:0] s5871, in5871_1, in5871_2;
    wire c5871;
    assign in5871_1 = {c2457};
    assign in5871_2 = {c2458};
    Full_Adder FA_5871(s5871, c5871, in5871_1, in5871_2, c2456);
    wire[0:0] s5872, in5872_1, in5872_2;
    wire c5872;
    assign in5872_1 = {c2460};
    assign in5872_2 = {c2461};
    Full_Adder FA_5872(s5872, c5872, in5872_1, in5872_2, c2459);
    wire[0:0] s5873, in5873_1, in5873_2;
    wire c5873;
    assign in5873_1 = {c2463};
    assign in5873_2 = {c2464};
    Full_Adder FA_5873(s5873, c5873, in5873_1, in5873_2, c2462);
    wire[0:0] s5874, in5874_1, in5874_2;
    wire c5874;
    assign in5874_1 = {s2466[0]};
    assign in5874_2 = {s2467[0]};
    Full_Adder FA_5874(s5874, c5874, in5874_1, in5874_2, s2465[0]);
    wire[0:0] s5875, in5875_1, in5875_2;
    wire c5875;
    assign in5875_1 = {s2469[0]};
    assign in5875_2 = {s2470[0]};
    Full_Adder FA_5875(s5875, c5875, in5875_1, in5875_2, s2468[0]);
    wire[0:0] s5876, in5876_1, in5876_2;
    wire c5876;
    assign in5876_1 = {s2472[0]};
    assign in5876_2 = {s2473[0]};
    Full_Adder FA_5876(s5876, c5876, in5876_1, in5876_2, s2471[0]);
    wire[0:0] s5877, in5877_1, in5877_2;
    wire c5877;
    assign in5877_1 = {s2475[0]};
    assign in5877_2 = {s2476[0]};
    Full_Adder FA_5877(s5877, c5877, in5877_1, in5877_2, s2474[0]);
    wire[0:0] s5878, in5878_1, in5878_2;
    wire c5878;
    assign in5878_1 = {s2478[0]};
    assign in5878_2 = {s2479[0]};
    Full_Adder FA_5878(s5878, c5878, in5878_1, in5878_2, s2477[0]);
    wire[0:0] s5879, in5879_1, in5879_2;
    wire c5879;
    assign in5879_1 = {s2481[0]};
    assign in5879_2 = {s2482[0]};
    Full_Adder FA_5879(s5879, c5879, in5879_1, in5879_2, s2480[0]);
    wire[0:0] s5880, in5880_1, in5880_2;
    wire c5880;
    assign in5880_1 = {s2484[0]};
    assign in5880_2 = {s2485[0]};
    Full_Adder FA_5880(s5880, c5880, in5880_1, in5880_2, s2483[0]);
    wire[0:0] s5881, in5881_1, in5881_2;
    wire c5881;
    assign in5881_1 = {s2487[0]};
    assign in5881_2 = {s2488[0]};
    Full_Adder FA_5881(s5881, c5881, in5881_1, in5881_2, s2486[0]);
    wire[0:0] s5882, in5882_1, in5882_2;
    wire c5882;
    assign in5882_1 = {s2490[0]};
    assign in5882_2 = {s2491[0]};
    Full_Adder FA_5882(s5882, c5882, in5882_1, in5882_2, s2489[0]);
    wire[0:0] s5883, in5883_1, in5883_2;
    wire c5883;
    assign in5883_1 = {s66[0]};
    assign in5883_2 = {c2465};
    Full_Adder FA_5883(s5883, c5883, in5883_1, in5883_2, s65[0]);
    wire[0:0] s5884, in5884_1, in5884_2;
    wire c5884;
    assign in5884_1 = {c2467};
    assign in5884_2 = {c2468};
    Full_Adder FA_5884(s5884, c5884, in5884_1, in5884_2, c2466);
    wire[0:0] s5885, in5885_1, in5885_2;
    wire c5885;
    assign in5885_1 = {c2470};
    assign in5885_2 = {c2471};
    Full_Adder FA_5885(s5885, c5885, in5885_1, in5885_2, c2469);
    wire[0:0] s5886, in5886_1, in5886_2;
    wire c5886;
    assign in5886_1 = {c2473};
    assign in5886_2 = {c2474};
    Full_Adder FA_5886(s5886, c5886, in5886_1, in5886_2, c2472);
    wire[0:0] s5887, in5887_1, in5887_2;
    wire c5887;
    assign in5887_1 = {c2476};
    assign in5887_2 = {c2477};
    Full_Adder FA_5887(s5887, c5887, in5887_1, in5887_2, c2475);
    wire[0:0] s5888, in5888_1, in5888_2;
    wire c5888;
    assign in5888_1 = {c2479};
    assign in5888_2 = {c2480};
    Full_Adder FA_5888(s5888, c5888, in5888_1, in5888_2, c2478);
    wire[0:0] s5889, in5889_1, in5889_2;
    wire c5889;
    assign in5889_1 = {c2482};
    assign in5889_2 = {c2483};
    Full_Adder FA_5889(s5889, c5889, in5889_1, in5889_2, c2481);
    wire[0:0] s5890, in5890_1, in5890_2;
    wire c5890;
    assign in5890_1 = {c2485};
    assign in5890_2 = {c2486};
    Full_Adder FA_5890(s5890, c5890, in5890_1, in5890_2, c2484);
    wire[0:0] s5891, in5891_1, in5891_2;
    wire c5891;
    assign in5891_1 = {c2488};
    assign in5891_2 = {c2489};
    Full_Adder FA_5891(s5891, c5891, in5891_1, in5891_2, c2487);
    wire[0:0] s5892, in5892_1, in5892_2;
    wire c5892;
    assign in5892_1 = {c2491};
    assign in5892_2 = {c2492};
    Full_Adder FA_5892(s5892, c5892, in5892_1, in5892_2, c2490);
    wire[0:0] s5893, in5893_1, in5893_2;
    wire c5893;
    assign in5893_1 = {s2494[0]};
    assign in5893_2 = {s2495[0]};
    Full_Adder FA_5893(s5893, c5893, in5893_1, in5893_2, s2493[0]);
    wire[0:0] s5894, in5894_1, in5894_2;
    wire c5894;
    assign in5894_1 = {s2497[0]};
    assign in5894_2 = {s2498[0]};
    Full_Adder FA_5894(s5894, c5894, in5894_1, in5894_2, s2496[0]);
    wire[0:0] s5895, in5895_1, in5895_2;
    wire c5895;
    assign in5895_1 = {s2500[0]};
    assign in5895_2 = {s2501[0]};
    Full_Adder FA_5895(s5895, c5895, in5895_1, in5895_2, s2499[0]);
    wire[0:0] s5896, in5896_1, in5896_2;
    wire c5896;
    assign in5896_1 = {s2503[0]};
    assign in5896_2 = {s2504[0]};
    Full_Adder FA_5896(s5896, c5896, in5896_1, in5896_2, s2502[0]);
    wire[0:0] s5897, in5897_1, in5897_2;
    wire c5897;
    assign in5897_1 = {s2506[0]};
    assign in5897_2 = {s2507[0]};
    Full_Adder FA_5897(s5897, c5897, in5897_1, in5897_2, s2505[0]);
    wire[0:0] s5898, in5898_1, in5898_2;
    wire c5898;
    assign in5898_1 = {s2509[0]};
    assign in5898_2 = {s2510[0]};
    Full_Adder FA_5898(s5898, c5898, in5898_1, in5898_2, s2508[0]);
    wire[0:0] s5899, in5899_1, in5899_2;
    wire c5899;
    assign in5899_1 = {s2512[0]};
    assign in5899_2 = {s2513[0]};
    Full_Adder FA_5899(s5899, c5899, in5899_1, in5899_2, s2511[0]);
    wire[0:0] s5900, in5900_1, in5900_2;
    wire c5900;
    assign in5900_1 = {s2515[0]};
    assign in5900_2 = {s2516[0]};
    Full_Adder FA_5900(s5900, c5900, in5900_1, in5900_2, s2514[0]);
    wire[0:0] s5901, in5901_1, in5901_2;
    wire c5901;
    assign in5901_1 = {s2518[0]};
    assign in5901_2 = {s2519[0]};
    Full_Adder FA_5901(s5901, c5901, in5901_1, in5901_2, s2517[0]);
    wire[0:0] s5902, in5902_1, in5902_2;
    wire c5902;
    assign in5902_1 = {s78[0]};
    assign in5902_2 = {c2493};
    Full_Adder FA_5902(s5902, c5902, in5902_1, in5902_2, s77[0]);
    wire[0:0] s5903, in5903_1, in5903_2;
    wire c5903;
    assign in5903_1 = {c2495};
    assign in5903_2 = {c2496};
    Full_Adder FA_5903(s5903, c5903, in5903_1, in5903_2, c2494);
    wire[0:0] s5904, in5904_1, in5904_2;
    wire c5904;
    assign in5904_1 = {c2498};
    assign in5904_2 = {c2499};
    Full_Adder FA_5904(s5904, c5904, in5904_1, in5904_2, c2497);
    wire[0:0] s5905, in5905_1, in5905_2;
    wire c5905;
    assign in5905_1 = {c2501};
    assign in5905_2 = {c2502};
    Full_Adder FA_5905(s5905, c5905, in5905_1, in5905_2, c2500);
    wire[0:0] s5906, in5906_1, in5906_2;
    wire c5906;
    assign in5906_1 = {c2504};
    assign in5906_2 = {c2505};
    Full_Adder FA_5906(s5906, c5906, in5906_1, in5906_2, c2503);
    wire[0:0] s5907, in5907_1, in5907_2;
    wire c5907;
    assign in5907_1 = {c2507};
    assign in5907_2 = {c2508};
    Full_Adder FA_5907(s5907, c5907, in5907_1, in5907_2, c2506);
    wire[0:0] s5908, in5908_1, in5908_2;
    wire c5908;
    assign in5908_1 = {c2510};
    assign in5908_2 = {c2511};
    Full_Adder FA_5908(s5908, c5908, in5908_1, in5908_2, c2509);
    wire[0:0] s5909, in5909_1, in5909_2;
    wire c5909;
    assign in5909_1 = {c2513};
    assign in5909_2 = {c2514};
    Full_Adder FA_5909(s5909, c5909, in5909_1, in5909_2, c2512);
    wire[0:0] s5910, in5910_1, in5910_2;
    wire c5910;
    assign in5910_1 = {c2516};
    assign in5910_2 = {c2517};
    Full_Adder FA_5910(s5910, c5910, in5910_1, in5910_2, c2515);
    wire[0:0] s5911, in5911_1, in5911_2;
    wire c5911;
    assign in5911_1 = {c2519};
    assign in5911_2 = {c2520};
    Full_Adder FA_5911(s5911, c5911, in5911_1, in5911_2, c2518);
    wire[0:0] s5912, in5912_1, in5912_2;
    wire c5912;
    assign in5912_1 = {s2522[0]};
    assign in5912_2 = {s2523[0]};
    Full_Adder FA_5912(s5912, c5912, in5912_1, in5912_2, s2521[0]);
    wire[0:0] s5913, in5913_1, in5913_2;
    wire c5913;
    assign in5913_1 = {s2525[0]};
    assign in5913_2 = {s2526[0]};
    Full_Adder FA_5913(s5913, c5913, in5913_1, in5913_2, s2524[0]);
    wire[0:0] s5914, in5914_1, in5914_2;
    wire c5914;
    assign in5914_1 = {s2528[0]};
    assign in5914_2 = {s2529[0]};
    Full_Adder FA_5914(s5914, c5914, in5914_1, in5914_2, s2527[0]);
    wire[0:0] s5915, in5915_1, in5915_2;
    wire c5915;
    assign in5915_1 = {s2531[0]};
    assign in5915_2 = {s2532[0]};
    Full_Adder FA_5915(s5915, c5915, in5915_1, in5915_2, s2530[0]);
    wire[0:0] s5916, in5916_1, in5916_2;
    wire c5916;
    assign in5916_1 = {s2534[0]};
    assign in5916_2 = {s2535[0]};
    Full_Adder FA_5916(s5916, c5916, in5916_1, in5916_2, s2533[0]);
    wire[0:0] s5917, in5917_1, in5917_2;
    wire c5917;
    assign in5917_1 = {s2537[0]};
    assign in5917_2 = {s2538[0]};
    Full_Adder FA_5917(s5917, c5917, in5917_1, in5917_2, s2536[0]);
    wire[0:0] s5918, in5918_1, in5918_2;
    wire c5918;
    assign in5918_1 = {s2540[0]};
    assign in5918_2 = {s2541[0]};
    Full_Adder FA_5918(s5918, c5918, in5918_1, in5918_2, s2539[0]);
    wire[0:0] s5919, in5919_1, in5919_2;
    wire c5919;
    assign in5919_1 = {s2543[0]};
    assign in5919_2 = {s2544[0]};
    Full_Adder FA_5919(s5919, c5919, in5919_1, in5919_2, s2542[0]);
    wire[0:0] s5920, in5920_1, in5920_2;
    wire c5920;
    assign in5920_1 = {s2546[0]};
    assign in5920_2 = {s2547[0]};
    Full_Adder FA_5920(s5920, c5920, in5920_1, in5920_2, s2545[0]);
    wire[0:0] s5921, in5921_1, in5921_2;
    wire c5921;
    assign in5921_1 = {s91[0]};
    assign in5921_2 = {c2521};
    Full_Adder FA_5921(s5921, c5921, in5921_1, in5921_2, s90[0]);
    wire[0:0] s5922, in5922_1, in5922_2;
    wire c5922;
    assign in5922_1 = {c2523};
    assign in5922_2 = {c2524};
    Full_Adder FA_5922(s5922, c5922, in5922_1, in5922_2, c2522);
    wire[0:0] s5923, in5923_1, in5923_2;
    wire c5923;
    assign in5923_1 = {c2526};
    assign in5923_2 = {c2527};
    Full_Adder FA_5923(s5923, c5923, in5923_1, in5923_2, c2525);
    wire[0:0] s5924, in5924_1, in5924_2;
    wire c5924;
    assign in5924_1 = {c2529};
    assign in5924_2 = {c2530};
    Full_Adder FA_5924(s5924, c5924, in5924_1, in5924_2, c2528);
    wire[0:0] s5925, in5925_1, in5925_2;
    wire c5925;
    assign in5925_1 = {c2532};
    assign in5925_2 = {c2533};
    Full_Adder FA_5925(s5925, c5925, in5925_1, in5925_2, c2531);
    wire[0:0] s5926, in5926_1, in5926_2;
    wire c5926;
    assign in5926_1 = {c2535};
    assign in5926_2 = {c2536};
    Full_Adder FA_5926(s5926, c5926, in5926_1, in5926_2, c2534);
    wire[0:0] s5927, in5927_1, in5927_2;
    wire c5927;
    assign in5927_1 = {c2538};
    assign in5927_2 = {c2539};
    Full_Adder FA_5927(s5927, c5927, in5927_1, in5927_2, c2537);
    wire[0:0] s5928, in5928_1, in5928_2;
    wire c5928;
    assign in5928_1 = {c2541};
    assign in5928_2 = {c2542};
    Full_Adder FA_5928(s5928, c5928, in5928_1, in5928_2, c2540);
    wire[0:0] s5929, in5929_1, in5929_2;
    wire c5929;
    assign in5929_1 = {c2544};
    assign in5929_2 = {c2545};
    Full_Adder FA_5929(s5929, c5929, in5929_1, in5929_2, c2543);
    wire[0:0] s5930, in5930_1, in5930_2;
    wire c5930;
    assign in5930_1 = {c2547};
    assign in5930_2 = {c2548};
    Full_Adder FA_5930(s5930, c5930, in5930_1, in5930_2, c2546);
    wire[0:0] s5931, in5931_1, in5931_2;
    wire c5931;
    assign in5931_1 = {s2550[0]};
    assign in5931_2 = {s2551[0]};
    Full_Adder FA_5931(s5931, c5931, in5931_1, in5931_2, s2549[0]);
    wire[0:0] s5932, in5932_1, in5932_2;
    wire c5932;
    assign in5932_1 = {s2553[0]};
    assign in5932_2 = {s2554[0]};
    Full_Adder FA_5932(s5932, c5932, in5932_1, in5932_2, s2552[0]);
    wire[0:0] s5933, in5933_1, in5933_2;
    wire c5933;
    assign in5933_1 = {s2556[0]};
    assign in5933_2 = {s2557[0]};
    Full_Adder FA_5933(s5933, c5933, in5933_1, in5933_2, s2555[0]);
    wire[0:0] s5934, in5934_1, in5934_2;
    wire c5934;
    assign in5934_1 = {s2559[0]};
    assign in5934_2 = {s2560[0]};
    Full_Adder FA_5934(s5934, c5934, in5934_1, in5934_2, s2558[0]);
    wire[0:0] s5935, in5935_1, in5935_2;
    wire c5935;
    assign in5935_1 = {s2562[0]};
    assign in5935_2 = {s2563[0]};
    Full_Adder FA_5935(s5935, c5935, in5935_1, in5935_2, s2561[0]);
    wire[0:0] s5936, in5936_1, in5936_2;
    wire c5936;
    assign in5936_1 = {s2565[0]};
    assign in5936_2 = {s2566[0]};
    Full_Adder FA_5936(s5936, c5936, in5936_1, in5936_2, s2564[0]);
    wire[0:0] s5937, in5937_1, in5937_2;
    wire c5937;
    assign in5937_1 = {s2568[0]};
    assign in5937_2 = {s2569[0]};
    Full_Adder FA_5937(s5937, c5937, in5937_1, in5937_2, s2567[0]);
    wire[0:0] s5938, in5938_1, in5938_2;
    wire c5938;
    assign in5938_1 = {s2571[0]};
    assign in5938_2 = {s2572[0]};
    Full_Adder FA_5938(s5938, c5938, in5938_1, in5938_2, s2570[0]);
    wire[0:0] s5939, in5939_1, in5939_2;
    wire c5939;
    assign in5939_1 = {s2574[0]};
    assign in5939_2 = {s2575[0]};
    Full_Adder FA_5939(s5939, c5939, in5939_1, in5939_2, s2573[0]);
    wire[0:0] s5940, in5940_1, in5940_2;
    wire c5940;
    assign in5940_1 = {s105[0]};
    assign in5940_2 = {c2549};
    Full_Adder FA_5940(s5940, c5940, in5940_1, in5940_2, s104[0]);
    wire[0:0] s5941, in5941_1, in5941_2;
    wire c5941;
    assign in5941_1 = {c2551};
    assign in5941_2 = {c2552};
    Full_Adder FA_5941(s5941, c5941, in5941_1, in5941_2, c2550);
    wire[0:0] s5942, in5942_1, in5942_2;
    wire c5942;
    assign in5942_1 = {c2554};
    assign in5942_2 = {c2555};
    Full_Adder FA_5942(s5942, c5942, in5942_1, in5942_2, c2553);
    wire[0:0] s5943, in5943_1, in5943_2;
    wire c5943;
    assign in5943_1 = {c2557};
    assign in5943_2 = {c2558};
    Full_Adder FA_5943(s5943, c5943, in5943_1, in5943_2, c2556);
    wire[0:0] s5944, in5944_1, in5944_2;
    wire c5944;
    assign in5944_1 = {c2560};
    assign in5944_2 = {c2561};
    Full_Adder FA_5944(s5944, c5944, in5944_1, in5944_2, c2559);
    wire[0:0] s5945, in5945_1, in5945_2;
    wire c5945;
    assign in5945_1 = {c2563};
    assign in5945_2 = {c2564};
    Full_Adder FA_5945(s5945, c5945, in5945_1, in5945_2, c2562);
    wire[0:0] s5946, in5946_1, in5946_2;
    wire c5946;
    assign in5946_1 = {c2566};
    assign in5946_2 = {c2567};
    Full_Adder FA_5946(s5946, c5946, in5946_1, in5946_2, c2565);
    wire[0:0] s5947, in5947_1, in5947_2;
    wire c5947;
    assign in5947_1 = {c2569};
    assign in5947_2 = {c2570};
    Full_Adder FA_5947(s5947, c5947, in5947_1, in5947_2, c2568);
    wire[0:0] s5948, in5948_1, in5948_2;
    wire c5948;
    assign in5948_1 = {c2572};
    assign in5948_2 = {c2573};
    Full_Adder FA_5948(s5948, c5948, in5948_1, in5948_2, c2571);
    wire[0:0] s5949, in5949_1, in5949_2;
    wire c5949;
    assign in5949_1 = {c2575};
    assign in5949_2 = {c2576};
    Full_Adder FA_5949(s5949, c5949, in5949_1, in5949_2, c2574);
    wire[0:0] s5950, in5950_1, in5950_2;
    wire c5950;
    assign in5950_1 = {s2578[0]};
    assign in5950_2 = {s2579[0]};
    Full_Adder FA_5950(s5950, c5950, in5950_1, in5950_2, s2577[0]);
    wire[0:0] s5951, in5951_1, in5951_2;
    wire c5951;
    assign in5951_1 = {s2581[0]};
    assign in5951_2 = {s2582[0]};
    Full_Adder FA_5951(s5951, c5951, in5951_1, in5951_2, s2580[0]);
    wire[0:0] s5952, in5952_1, in5952_2;
    wire c5952;
    assign in5952_1 = {s2584[0]};
    assign in5952_2 = {s2585[0]};
    Full_Adder FA_5952(s5952, c5952, in5952_1, in5952_2, s2583[0]);
    wire[0:0] s5953, in5953_1, in5953_2;
    wire c5953;
    assign in5953_1 = {s2587[0]};
    assign in5953_2 = {s2588[0]};
    Full_Adder FA_5953(s5953, c5953, in5953_1, in5953_2, s2586[0]);
    wire[0:0] s5954, in5954_1, in5954_2;
    wire c5954;
    assign in5954_1 = {s2590[0]};
    assign in5954_2 = {s2591[0]};
    Full_Adder FA_5954(s5954, c5954, in5954_1, in5954_2, s2589[0]);
    wire[0:0] s5955, in5955_1, in5955_2;
    wire c5955;
    assign in5955_1 = {s2593[0]};
    assign in5955_2 = {s2594[0]};
    Full_Adder FA_5955(s5955, c5955, in5955_1, in5955_2, s2592[0]);
    wire[0:0] s5956, in5956_1, in5956_2;
    wire c5956;
    assign in5956_1 = {s2596[0]};
    assign in5956_2 = {s2597[0]};
    Full_Adder FA_5956(s5956, c5956, in5956_1, in5956_2, s2595[0]);
    wire[0:0] s5957, in5957_1, in5957_2;
    wire c5957;
    assign in5957_1 = {s2599[0]};
    assign in5957_2 = {s2600[0]};
    Full_Adder FA_5957(s5957, c5957, in5957_1, in5957_2, s2598[0]);
    wire[0:0] s5958, in5958_1, in5958_2;
    wire c5958;
    assign in5958_1 = {s2602[0]};
    assign in5958_2 = {s2603[0]};
    Full_Adder FA_5958(s5958, c5958, in5958_1, in5958_2, s2601[0]);
    wire[0:0] s5959, in5959_1, in5959_2;
    wire c5959;
    assign in5959_1 = {s120[0]};
    assign in5959_2 = {c2577};
    Full_Adder FA_5959(s5959, c5959, in5959_1, in5959_2, s119[0]);
    wire[0:0] s5960, in5960_1, in5960_2;
    wire c5960;
    assign in5960_1 = {c2579};
    assign in5960_2 = {c2580};
    Full_Adder FA_5960(s5960, c5960, in5960_1, in5960_2, c2578);
    wire[0:0] s5961, in5961_1, in5961_2;
    wire c5961;
    assign in5961_1 = {c2582};
    assign in5961_2 = {c2583};
    Full_Adder FA_5961(s5961, c5961, in5961_1, in5961_2, c2581);
    wire[0:0] s5962, in5962_1, in5962_2;
    wire c5962;
    assign in5962_1 = {c2585};
    assign in5962_2 = {c2586};
    Full_Adder FA_5962(s5962, c5962, in5962_1, in5962_2, c2584);
    wire[0:0] s5963, in5963_1, in5963_2;
    wire c5963;
    assign in5963_1 = {c2588};
    assign in5963_2 = {c2589};
    Full_Adder FA_5963(s5963, c5963, in5963_1, in5963_2, c2587);
    wire[0:0] s5964, in5964_1, in5964_2;
    wire c5964;
    assign in5964_1 = {c2591};
    assign in5964_2 = {c2592};
    Full_Adder FA_5964(s5964, c5964, in5964_1, in5964_2, c2590);
    wire[0:0] s5965, in5965_1, in5965_2;
    wire c5965;
    assign in5965_1 = {c2594};
    assign in5965_2 = {c2595};
    Full_Adder FA_5965(s5965, c5965, in5965_1, in5965_2, c2593);
    wire[0:0] s5966, in5966_1, in5966_2;
    wire c5966;
    assign in5966_1 = {c2597};
    assign in5966_2 = {c2598};
    Full_Adder FA_5966(s5966, c5966, in5966_1, in5966_2, c2596);
    wire[0:0] s5967, in5967_1, in5967_2;
    wire c5967;
    assign in5967_1 = {c2600};
    assign in5967_2 = {c2601};
    Full_Adder FA_5967(s5967, c5967, in5967_1, in5967_2, c2599);
    wire[0:0] s5968, in5968_1, in5968_2;
    wire c5968;
    assign in5968_1 = {c2603};
    assign in5968_2 = {c2604};
    Full_Adder FA_5968(s5968, c5968, in5968_1, in5968_2, c2602);
    wire[0:0] s5969, in5969_1, in5969_2;
    wire c5969;
    assign in5969_1 = {s2606[0]};
    assign in5969_2 = {s2607[0]};
    Full_Adder FA_5969(s5969, c5969, in5969_1, in5969_2, s2605[0]);
    wire[0:0] s5970, in5970_1, in5970_2;
    wire c5970;
    assign in5970_1 = {s2609[0]};
    assign in5970_2 = {s2610[0]};
    Full_Adder FA_5970(s5970, c5970, in5970_1, in5970_2, s2608[0]);
    wire[0:0] s5971, in5971_1, in5971_2;
    wire c5971;
    assign in5971_1 = {s2612[0]};
    assign in5971_2 = {s2613[0]};
    Full_Adder FA_5971(s5971, c5971, in5971_1, in5971_2, s2611[0]);
    wire[0:0] s5972, in5972_1, in5972_2;
    wire c5972;
    assign in5972_1 = {s2615[0]};
    assign in5972_2 = {s2616[0]};
    Full_Adder FA_5972(s5972, c5972, in5972_1, in5972_2, s2614[0]);
    wire[0:0] s5973, in5973_1, in5973_2;
    wire c5973;
    assign in5973_1 = {s2618[0]};
    assign in5973_2 = {s2619[0]};
    Full_Adder FA_5973(s5973, c5973, in5973_1, in5973_2, s2617[0]);
    wire[0:0] s5974, in5974_1, in5974_2;
    wire c5974;
    assign in5974_1 = {s2621[0]};
    assign in5974_2 = {s2622[0]};
    Full_Adder FA_5974(s5974, c5974, in5974_1, in5974_2, s2620[0]);
    wire[0:0] s5975, in5975_1, in5975_2;
    wire c5975;
    assign in5975_1 = {s2624[0]};
    assign in5975_2 = {s2625[0]};
    Full_Adder FA_5975(s5975, c5975, in5975_1, in5975_2, s2623[0]);
    wire[0:0] s5976, in5976_1, in5976_2;
    wire c5976;
    assign in5976_1 = {s2627[0]};
    assign in5976_2 = {s2628[0]};
    Full_Adder FA_5976(s5976, c5976, in5976_1, in5976_2, s2626[0]);
    wire[0:0] s5977, in5977_1, in5977_2;
    wire c5977;
    assign in5977_1 = {s2630[0]};
    assign in5977_2 = {s2631[0]};
    Full_Adder FA_5977(s5977, c5977, in5977_1, in5977_2, s2629[0]);
    wire[0:0] s5978, in5978_1, in5978_2;
    wire c5978;
    assign in5978_1 = {s136[0]};
    assign in5978_2 = {c2605};
    Full_Adder FA_5978(s5978, c5978, in5978_1, in5978_2, s135[0]);
    wire[0:0] s5979, in5979_1, in5979_2;
    wire c5979;
    assign in5979_1 = {c2607};
    assign in5979_2 = {c2608};
    Full_Adder FA_5979(s5979, c5979, in5979_1, in5979_2, c2606);
    wire[0:0] s5980, in5980_1, in5980_2;
    wire c5980;
    assign in5980_1 = {c2610};
    assign in5980_2 = {c2611};
    Full_Adder FA_5980(s5980, c5980, in5980_1, in5980_2, c2609);
    wire[0:0] s5981, in5981_1, in5981_2;
    wire c5981;
    assign in5981_1 = {c2613};
    assign in5981_2 = {c2614};
    Full_Adder FA_5981(s5981, c5981, in5981_1, in5981_2, c2612);
    wire[0:0] s5982, in5982_1, in5982_2;
    wire c5982;
    assign in5982_1 = {c2616};
    assign in5982_2 = {c2617};
    Full_Adder FA_5982(s5982, c5982, in5982_1, in5982_2, c2615);
    wire[0:0] s5983, in5983_1, in5983_2;
    wire c5983;
    assign in5983_1 = {c2619};
    assign in5983_2 = {c2620};
    Full_Adder FA_5983(s5983, c5983, in5983_1, in5983_2, c2618);
    wire[0:0] s5984, in5984_1, in5984_2;
    wire c5984;
    assign in5984_1 = {c2622};
    assign in5984_2 = {c2623};
    Full_Adder FA_5984(s5984, c5984, in5984_1, in5984_2, c2621);
    wire[0:0] s5985, in5985_1, in5985_2;
    wire c5985;
    assign in5985_1 = {c2625};
    assign in5985_2 = {c2626};
    Full_Adder FA_5985(s5985, c5985, in5985_1, in5985_2, c2624);
    wire[0:0] s5986, in5986_1, in5986_2;
    wire c5986;
    assign in5986_1 = {c2628};
    assign in5986_2 = {c2629};
    Full_Adder FA_5986(s5986, c5986, in5986_1, in5986_2, c2627);
    wire[0:0] s5987, in5987_1, in5987_2;
    wire c5987;
    assign in5987_1 = {c2631};
    assign in5987_2 = {c2632};
    Full_Adder FA_5987(s5987, c5987, in5987_1, in5987_2, c2630);
    wire[0:0] s5988, in5988_1, in5988_2;
    wire c5988;
    assign in5988_1 = {s2634[0]};
    assign in5988_2 = {s2635[0]};
    Full_Adder FA_5988(s5988, c5988, in5988_1, in5988_2, s2633[0]);
    wire[0:0] s5989, in5989_1, in5989_2;
    wire c5989;
    assign in5989_1 = {s2637[0]};
    assign in5989_2 = {s2638[0]};
    Full_Adder FA_5989(s5989, c5989, in5989_1, in5989_2, s2636[0]);
    wire[0:0] s5990, in5990_1, in5990_2;
    wire c5990;
    assign in5990_1 = {s2640[0]};
    assign in5990_2 = {s2641[0]};
    Full_Adder FA_5990(s5990, c5990, in5990_1, in5990_2, s2639[0]);
    wire[0:0] s5991, in5991_1, in5991_2;
    wire c5991;
    assign in5991_1 = {s2643[0]};
    assign in5991_2 = {s2644[0]};
    Full_Adder FA_5991(s5991, c5991, in5991_1, in5991_2, s2642[0]);
    wire[0:0] s5992, in5992_1, in5992_2;
    wire c5992;
    assign in5992_1 = {s2646[0]};
    assign in5992_2 = {s2647[0]};
    Full_Adder FA_5992(s5992, c5992, in5992_1, in5992_2, s2645[0]);
    wire[0:0] s5993, in5993_1, in5993_2;
    wire c5993;
    assign in5993_1 = {s2649[0]};
    assign in5993_2 = {s2650[0]};
    Full_Adder FA_5993(s5993, c5993, in5993_1, in5993_2, s2648[0]);
    wire[0:0] s5994, in5994_1, in5994_2;
    wire c5994;
    assign in5994_1 = {s2652[0]};
    assign in5994_2 = {s2653[0]};
    Full_Adder FA_5994(s5994, c5994, in5994_1, in5994_2, s2651[0]);
    wire[0:0] s5995, in5995_1, in5995_2;
    wire c5995;
    assign in5995_1 = {s2655[0]};
    assign in5995_2 = {s2656[0]};
    Full_Adder FA_5995(s5995, c5995, in5995_1, in5995_2, s2654[0]);
    wire[0:0] s5996, in5996_1, in5996_2;
    wire c5996;
    assign in5996_1 = {s2658[0]};
    assign in5996_2 = {s2659[0]};
    Full_Adder FA_5996(s5996, c5996, in5996_1, in5996_2, s2657[0]);
    wire[0:0] s5997, in5997_1, in5997_2;
    wire c5997;
    assign in5997_1 = {s153[0]};
    assign in5997_2 = {c2633};
    Full_Adder FA_5997(s5997, c5997, in5997_1, in5997_2, s152[0]);
    wire[0:0] s5998, in5998_1, in5998_2;
    wire c5998;
    assign in5998_1 = {c2635};
    assign in5998_2 = {c2636};
    Full_Adder FA_5998(s5998, c5998, in5998_1, in5998_2, c2634);
    wire[0:0] s5999, in5999_1, in5999_2;
    wire c5999;
    assign in5999_1 = {c2638};
    assign in5999_2 = {c2639};
    Full_Adder FA_5999(s5999, c5999, in5999_1, in5999_2, c2637);
    wire[0:0] s6000, in6000_1, in6000_2;
    wire c6000;
    assign in6000_1 = {c2641};
    assign in6000_2 = {c2642};
    Full_Adder FA_6000(s6000, c6000, in6000_1, in6000_2, c2640);
    wire[0:0] s6001, in6001_1, in6001_2;
    wire c6001;
    assign in6001_1 = {c2644};
    assign in6001_2 = {c2645};
    Full_Adder FA_6001(s6001, c6001, in6001_1, in6001_2, c2643);
    wire[0:0] s6002, in6002_1, in6002_2;
    wire c6002;
    assign in6002_1 = {c2647};
    assign in6002_2 = {c2648};
    Full_Adder FA_6002(s6002, c6002, in6002_1, in6002_2, c2646);
    wire[0:0] s6003, in6003_1, in6003_2;
    wire c6003;
    assign in6003_1 = {c2650};
    assign in6003_2 = {c2651};
    Full_Adder FA_6003(s6003, c6003, in6003_1, in6003_2, c2649);
    wire[0:0] s6004, in6004_1, in6004_2;
    wire c6004;
    assign in6004_1 = {c2653};
    assign in6004_2 = {c2654};
    Full_Adder FA_6004(s6004, c6004, in6004_1, in6004_2, c2652);
    wire[0:0] s6005, in6005_1, in6005_2;
    wire c6005;
    assign in6005_1 = {c2656};
    assign in6005_2 = {c2657};
    Full_Adder FA_6005(s6005, c6005, in6005_1, in6005_2, c2655);
    wire[0:0] s6006, in6006_1, in6006_2;
    wire c6006;
    assign in6006_1 = {c2659};
    assign in6006_2 = {c2660};
    Full_Adder FA_6006(s6006, c6006, in6006_1, in6006_2, c2658);
    wire[0:0] s6007, in6007_1, in6007_2;
    wire c6007;
    assign in6007_1 = {s2662[0]};
    assign in6007_2 = {s2663[0]};
    Full_Adder FA_6007(s6007, c6007, in6007_1, in6007_2, s2661[0]);
    wire[0:0] s6008, in6008_1, in6008_2;
    wire c6008;
    assign in6008_1 = {s2665[0]};
    assign in6008_2 = {s2666[0]};
    Full_Adder FA_6008(s6008, c6008, in6008_1, in6008_2, s2664[0]);
    wire[0:0] s6009, in6009_1, in6009_2;
    wire c6009;
    assign in6009_1 = {s2668[0]};
    assign in6009_2 = {s2669[0]};
    Full_Adder FA_6009(s6009, c6009, in6009_1, in6009_2, s2667[0]);
    wire[0:0] s6010, in6010_1, in6010_2;
    wire c6010;
    assign in6010_1 = {s2671[0]};
    assign in6010_2 = {s2672[0]};
    Full_Adder FA_6010(s6010, c6010, in6010_1, in6010_2, s2670[0]);
    wire[0:0] s6011, in6011_1, in6011_2;
    wire c6011;
    assign in6011_1 = {s2674[0]};
    assign in6011_2 = {s2675[0]};
    Full_Adder FA_6011(s6011, c6011, in6011_1, in6011_2, s2673[0]);
    wire[0:0] s6012, in6012_1, in6012_2;
    wire c6012;
    assign in6012_1 = {s2677[0]};
    assign in6012_2 = {s2678[0]};
    Full_Adder FA_6012(s6012, c6012, in6012_1, in6012_2, s2676[0]);
    wire[0:0] s6013, in6013_1, in6013_2;
    wire c6013;
    assign in6013_1 = {s2680[0]};
    assign in6013_2 = {s2681[0]};
    Full_Adder FA_6013(s6013, c6013, in6013_1, in6013_2, s2679[0]);
    wire[0:0] s6014, in6014_1, in6014_2;
    wire c6014;
    assign in6014_1 = {s2683[0]};
    assign in6014_2 = {s2684[0]};
    Full_Adder FA_6014(s6014, c6014, in6014_1, in6014_2, s2682[0]);
    wire[0:0] s6015, in6015_1, in6015_2;
    wire c6015;
    assign in6015_1 = {s2686[0]};
    assign in6015_2 = {s2687[0]};
    Full_Adder FA_6015(s6015, c6015, in6015_1, in6015_2, s2685[0]);
    wire[0:0] s6016, in6016_1, in6016_2;
    wire c6016;
    assign in6016_1 = {s171[0]};
    assign in6016_2 = {c2661};
    Full_Adder FA_6016(s6016, c6016, in6016_1, in6016_2, s170[0]);
    wire[0:0] s6017, in6017_1, in6017_2;
    wire c6017;
    assign in6017_1 = {c2663};
    assign in6017_2 = {c2664};
    Full_Adder FA_6017(s6017, c6017, in6017_1, in6017_2, c2662);
    wire[0:0] s6018, in6018_1, in6018_2;
    wire c6018;
    assign in6018_1 = {c2666};
    assign in6018_2 = {c2667};
    Full_Adder FA_6018(s6018, c6018, in6018_1, in6018_2, c2665);
    wire[0:0] s6019, in6019_1, in6019_2;
    wire c6019;
    assign in6019_1 = {c2669};
    assign in6019_2 = {c2670};
    Full_Adder FA_6019(s6019, c6019, in6019_1, in6019_2, c2668);
    wire[0:0] s6020, in6020_1, in6020_2;
    wire c6020;
    assign in6020_1 = {c2672};
    assign in6020_2 = {c2673};
    Full_Adder FA_6020(s6020, c6020, in6020_1, in6020_2, c2671);
    wire[0:0] s6021, in6021_1, in6021_2;
    wire c6021;
    assign in6021_1 = {c2675};
    assign in6021_2 = {c2676};
    Full_Adder FA_6021(s6021, c6021, in6021_1, in6021_2, c2674);
    wire[0:0] s6022, in6022_1, in6022_2;
    wire c6022;
    assign in6022_1 = {c2678};
    assign in6022_2 = {c2679};
    Full_Adder FA_6022(s6022, c6022, in6022_1, in6022_2, c2677);
    wire[0:0] s6023, in6023_1, in6023_2;
    wire c6023;
    assign in6023_1 = {c2681};
    assign in6023_2 = {c2682};
    Full_Adder FA_6023(s6023, c6023, in6023_1, in6023_2, c2680);
    wire[0:0] s6024, in6024_1, in6024_2;
    wire c6024;
    assign in6024_1 = {c2684};
    assign in6024_2 = {c2685};
    Full_Adder FA_6024(s6024, c6024, in6024_1, in6024_2, c2683);
    wire[0:0] s6025, in6025_1, in6025_2;
    wire c6025;
    assign in6025_1 = {c2687};
    assign in6025_2 = {c2688};
    Full_Adder FA_6025(s6025, c6025, in6025_1, in6025_2, c2686);
    wire[0:0] s6026, in6026_1, in6026_2;
    wire c6026;
    assign in6026_1 = {s2690[0]};
    assign in6026_2 = {s2691[0]};
    Full_Adder FA_6026(s6026, c6026, in6026_1, in6026_2, s2689[0]);
    wire[0:0] s6027, in6027_1, in6027_2;
    wire c6027;
    assign in6027_1 = {s2693[0]};
    assign in6027_2 = {s2694[0]};
    Full_Adder FA_6027(s6027, c6027, in6027_1, in6027_2, s2692[0]);
    wire[0:0] s6028, in6028_1, in6028_2;
    wire c6028;
    assign in6028_1 = {s2696[0]};
    assign in6028_2 = {s2697[0]};
    Full_Adder FA_6028(s6028, c6028, in6028_1, in6028_2, s2695[0]);
    wire[0:0] s6029, in6029_1, in6029_2;
    wire c6029;
    assign in6029_1 = {s2699[0]};
    assign in6029_2 = {s2700[0]};
    Full_Adder FA_6029(s6029, c6029, in6029_1, in6029_2, s2698[0]);
    wire[0:0] s6030, in6030_1, in6030_2;
    wire c6030;
    assign in6030_1 = {s2702[0]};
    assign in6030_2 = {s2703[0]};
    Full_Adder FA_6030(s6030, c6030, in6030_1, in6030_2, s2701[0]);
    wire[0:0] s6031, in6031_1, in6031_2;
    wire c6031;
    assign in6031_1 = {s2705[0]};
    assign in6031_2 = {s2706[0]};
    Full_Adder FA_6031(s6031, c6031, in6031_1, in6031_2, s2704[0]);
    wire[0:0] s6032, in6032_1, in6032_2;
    wire c6032;
    assign in6032_1 = {s2708[0]};
    assign in6032_2 = {s2709[0]};
    Full_Adder FA_6032(s6032, c6032, in6032_1, in6032_2, s2707[0]);
    wire[0:0] s6033, in6033_1, in6033_2;
    wire c6033;
    assign in6033_1 = {s2711[0]};
    assign in6033_2 = {s2712[0]};
    Full_Adder FA_6033(s6033, c6033, in6033_1, in6033_2, s2710[0]);
    wire[0:0] s6034, in6034_1, in6034_2;
    wire c6034;
    assign in6034_1 = {s2714[0]};
    assign in6034_2 = {s2715[0]};
    Full_Adder FA_6034(s6034, c6034, in6034_1, in6034_2, s2713[0]);
    wire[0:0] s6035, in6035_1, in6035_2;
    wire c6035;
    assign in6035_1 = {s190[0]};
    assign in6035_2 = {c2689};
    Full_Adder FA_6035(s6035, c6035, in6035_1, in6035_2, s189[0]);
    wire[0:0] s6036, in6036_1, in6036_2;
    wire c6036;
    assign in6036_1 = {c2691};
    assign in6036_2 = {c2692};
    Full_Adder FA_6036(s6036, c6036, in6036_1, in6036_2, c2690);
    wire[0:0] s6037, in6037_1, in6037_2;
    wire c6037;
    assign in6037_1 = {c2694};
    assign in6037_2 = {c2695};
    Full_Adder FA_6037(s6037, c6037, in6037_1, in6037_2, c2693);
    wire[0:0] s6038, in6038_1, in6038_2;
    wire c6038;
    assign in6038_1 = {c2697};
    assign in6038_2 = {c2698};
    Full_Adder FA_6038(s6038, c6038, in6038_1, in6038_2, c2696);
    wire[0:0] s6039, in6039_1, in6039_2;
    wire c6039;
    assign in6039_1 = {c2700};
    assign in6039_2 = {c2701};
    Full_Adder FA_6039(s6039, c6039, in6039_1, in6039_2, c2699);
    wire[0:0] s6040, in6040_1, in6040_2;
    wire c6040;
    assign in6040_1 = {c2703};
    assign in6040_2 = {c2704};
    Full_Adder FA_6040(s6040, c6040, in6040_1, in6040_2, c2702);
    wire[0:0] s6041, in6041_1, in6041_2;
    wire c6041;
    assign in6041_1 = {c2706};
    assign in6041_2 = {c2707};
    Full_Adder FA_6041(s6041, c6041, in6041_1, in6041_2, c2705);
    wire[0:0] s6042, in6042_1, in6042_2;
    wire c6042;
    assign in6042_1 = {c2709};
    assign in6042_2 = {c2710};
    Full_Adder FA_6042(s6042, c6042, in6042_1, in6042_2, c2708);
    wire[0:0] s6043, in6043_1, in6043_2;
    wire c6043;
    assign in6043_1 = {c2712};
    assign in6043_2 = {c2713};
    Full_Adder FA_6043(s6043, c6043, in6043_1, in6043_2, c2711);
    wire[0:0] s6044, in6044_1, in6044_2;
    wire c6044;
    assign in6044_1 = {c2715};
    assign in6044_2 = {c2716};
    Full_Adder FA_6044(s6044, c6044, in6044_1, in6044_2, c2714);
    wire[0:0] s6045, in6045_1, in6045_2;
    wire c6045;
    assign in6045_1 = {s2718[0]};
    assign in6045_2 = {s2719[0]};
    Full_Adder FA_6045(s6045, c6045, in6045_1, in6045_2, s2717[0]);
    wire[0:0] s6046, in6046_1, in6046_2;
    wire c6046;
    assign in6046_1 = {s2721[0]};
    assign in6046_2 = {s2722[0]};
    Full_Adder FA_6046(s6046, c6046, in6046_1, in6046_2, s2720[0]);
    wire[0:0] s6047, in6047_1, in6047_2;
    wire c6047;
    assign in6047_1 = {s2724[0]};
    assign in6047_2 = {s2725[0]};
    Full_Adder FA_6047(s6047, c6047, in6047_1, in6047_2, s2723[0]);
    wire[0:0] s6048, in6048_1, in6048_2;
    wire c6048;
    assign in6048_1 = {s2727[0]};
    assign in6048_2 = {s2728[0]};
    Full_Adder FA_6048(s6048, c6048, in6048_1, in6048_2, s2726[0]);
    wire[0:0] s6049, in6049_1, in6049_2;
    wire c6049;
    assign in6049_1 = {s2730[0]};
    assign in6049_2 = {s2731[0]};
    Full_Adder FA_6049(s6049, c6049, in6049_1, in6049_2, s2729[0]);
    wire[0:0] s6050, in6050_1, in6050_2;
    wire c6050;
    assign in6050_1 = {s2733[0]};
    assign in6050_2 = {s2734[0]};
    Full_Adder FA_6050(s6050, c6050, in6050_1, in6050_2, s2732[0]);
    wire[0:0] s6051, in6051_1, in6051_2;
    wire c6051;
    assign in6051_1 = {s2736[0]};
    assign in6051_2 = {s2737[0]};
    Full_Adder FA_6051(s6051, c6051, in6051_1, in6051_2, s2735[0]);
    wire[0:0] s6052, in6052_1, in6052_2;
    wire c6052;
    assign in6052_1 = {s2739[0]};
    assign in6052_2 = {s2740[0]};
    Full_Adder FA_6052(s6052, c6052, in6052_1, in6052_2, s2738[0]);
    wire[0:0] s6053, in6053_1, in6053_2;
    wire c6053;
    assign in6053_1 = {s2742[0]};
    assign in6053_2 = {s2743[0]};
    Full_Adder FA_6053(s6053, c6053, in6053_1, in6053_2, s2741[0]);
    wire[0:0] s6054, in6054_1, in6054_2;
    wire c6054;
    assign in6054_1 = {s210[0]};
    assign in6054_2 = {c2717};
    Full_Adder FA_6054(s6054, c6054, in6054_1, in6054_2, s209[0]);
    wire[0:0] s6055, in6055_1, in6055_2;
    wire c6055;
    assign in6055_1 = {c2719};
    assign in6055_2 = {c2720};
    Full_Adder FA_6055(s6055, c6055, in6055_1, in6055_2, c2718);
    wire[0:0] s6056, in6056_1, in6056_2;
    wire c6056;
    assign in6056_1 = {c2722};
    assign in6056_2 = {c2723};
    Full_Adder FA_6056(s6056, c6056, in6056_1, in6056_2, c2721);
    wire[0:0] s6057, in6057_1, in6057_2;
    wire c6057;
    assign in6057_1 = {c2725};
    assign in6057_2 = {c2726};
    Full_Adder FA_6057(s6057, c6057, in6057_1, in6057_2, c2724);
    wire[0:0] s6058, in6058_1, in6058_2;
    wire c6058;
    assign in6058_1 = {c2728};
    assign in6058_2 = {c2729};
    Full_Adder FA_6058(s6058, c6058, in6058_1, in6058_2, c2727);
    wire[0:0] s6059, in6059_1, in6059_2;
    wire c6059;
    assign in6059_1 = {c2731};
    assign in6059_2 = {c2732};
    Full_Adder FA_6059(s6059, c6059, in6059_1, in6059_2, c2730);
    wire[0:0] s6060, in6060_1, in6060_2;
    wire c6060;
    assign in6060_1 = {c2734};
    assign in6060_2 = {c2735};
    Full_Adder FA_6060(s6060, c6060, in6060_1, in6060_2, c2733);
    wire[0:0] s6061, in6061_1, in6061_2;
    wire c6061;
    assign in6061_1 = {c2737};
    assign in6061_2 = {c2738};
    Full_Adder FA_6061(s6061, c6061, in6061_1, in6061_2, c2736);
    wire[0:0] s6062, in6062_1, in6062_2;
    wire c6062;
    assign in6062_1 = {c2740};
    assign in6062_2 = {c2741};
    Full_Adder FA_6062(s6062, c6062, in6062_1, in6062_2, c2739);
    wire[0:0] s6063, in6063_1, in6063_2;
    wire c6063;
    assign in6063_1 = {c2743};
    assign in6063_2 = {c2744};
    Full_Adder FA_6063(s6063, c6063, in6063_1, in6063_2, c2742);
    wire[0:0] s6064, in6064_1, in6064_2;
    wire c6064;
    assign in6064_1 = {s2746[0]};
    assign in6064_2 = {s2747[0]};
    Full_Adder FA_6064(s6064, c6064, in6064_1, in6064_2, s2745[0]);
    wire[0:0] s6065, in6065_1, in6065_2;
    wire c6065;
    assign in6065_1 = {s2749[0]};
    assign in6065_2 = {s2750[0]};
    Full_Adder FA_6065(s6065, c6065, in6065_1, in6065_2, s2748[0]);
    wire[0:0] s6066, in6066_1, in6066_2;
    wire c6066;
    assign in6066_1 = {s2752[0]};
    assign in6066_2 = {s2753[0]};
    Full_Adder FA_6066(s6066, c6066, in6066_1, in6066_2, s2751[0]);
    wire[0:0] s6067, in6067_1, in6067_2;
    wire c6067;
    assign in6067_1 = {s2755[0]};
    assign in6067_2 = {s2756[0]};
    Full_Adder FA_6067(s6067, c6067, in6067_1, in6067_2, s2754[0]);
    wire[0:0] s6068, in6068_1, in6068_2;
    wire c6068;
    assign in6068_1 = {s2758[0]};
    assign in6068_2 = {s2759[0]};
    Full_Adder FA_6068(s6068, c6068, in6068_1, in6068_2, s2757[0]);
    wire[0:0] s6069, in6069_1, in6069_2;
    wire c6069;
    assign in6069_1 = {s2761[0]};
    assign in6069_2 = {s2762[0]};
    Full_Adder FA_6069(s6069, c6069, in6069_1, in6069_2, s2760[0]);
    wire[0:0] s6070, in6070_1, in6070_2;
    wire c6070;
    assign in6070_1 = {s2764[0]};
    assign in6070_2 = {s2765[0]};
    Full_Adder FA_6070(s6070, c6070, in6070_1, in6070_2, s2763[0]);
    wire[0:0] s6071, in6071_1, in6071_2;
    wire c6071;
    assign in6071_1 = {s2767[0]};
    assign in6071_2 = {s2768[0]};
    Full_Adder FA_6071(s6071, c6071, in6071_1, in6071_2, s2766[0]);
    wire[0:0] s6072, in6072_1, in6072_2;
    wire c6072;
    assign in6072_1 = {s2770[0]};
    assign in6072_2 = {s2771[0]};
    Full_Adder FA_6072(s6072, c6072, in6072_1, in6072_2, s2769[0]);
    wire[0:0] s6073, in6073_1, in6073_2;
    wire c6073;
    assign in6073_1 = {s231[0]};
    assign in6073_2 = {c2745};
    Full_Adder FA_6073(s6073, c6073, in6073_1, in6073_2, s230[0]);
    wire[0:0] s6074, in6074_1, in6074_2;
    wire c6074;
    assign in6074_1 = {c2747};
    assign in6074_2 = {c2748};
    Full_Adder FA_6074(s6074, c6074, in6074_1, in6074_2, c2746);
    wire[0:0] s6075, in6075_1, in6075_2;
    wire c6075;
    assign in6075_1 = {c2750};
    assign in6075_2 = {c2751};
    Full_Adder FA_6075(s6075, c6075, in6075_1, in6075_2, c2749);
    wire[0:0] s6076, in6076_1, in6076_2;
    wire c6076;
    assign in6076_1 = {c2753};
    assign in6076_2 = {c2754};
    Full_Adder FA_6076(s6076, c6076, in6076_1, in6076_2, c2752);
    wire[0:0] s6077, in6077_1, in6077_2;
    wire c6077;
    assign in6077_1 = {c2756};
    assign in6077_2 = {c2757};
    Full_Adder FA_6077(s6077, c6077, in6077_1, in6077_2, c2755);
    wire[0:0] s6078, in6078_1, in6078_2;
    wire c6078;
    assign in6078_1 = {c2759};
    assign in6078_2 = {c2760};
    Full_Adder FA_6078(s6078, c6078, in6078_1, in6078_2, c2758);
    wire[0:0] s6079, in6079_1, in6079_2;
    wire c6079;
    assign in6079_1 = {c2762};
    assign in6079_2 = {c2763};
    Full_Adder FA_6079(s6079, c6079, in6079_1, in6079_2, c2761);
    wire[0:0] s6080, in6080_1, in6080_2;
    wire c6080;
    assign in6080_1 = {c2765};
    assign in6080_2 = {c2766};
    Full_Adder FA_6080(s6080, c6080, in6080_1, in6080_2, c2764);
    wire[0:0] s6081, in6081_1, in6081_2;
    wire c6081;
    assign in6081_1 = {c2768};
    assign in6081_2 = {c2769};
    Full_Adder FA_6081(s6081, c6081, in6081_1, in6081_2, c2767);
    wire[0:0] s6082, in6082_1, in6082_2;
    wire c6082;
    assign in6082_1 = {c2771};
    assign in6082_2 = {c2772};
    Full_Adder FA_6082(s6082, c6082, in6082_1, in6082_2, c2770);
    wire[0:0] s6083, in6083_1, in6083_2;
    wire c6083;
    assign in6083_1 = {s2774[0]};
    assign in6083_2 = {s2775[0]};
    Full_Adder FA_6083(s6083, c6083, in6083_1, in6083_2, s2773[0]);
    wire[0:0] s6084, in6084_1, in6084_2;
    wire c6084;
    assign in6084_1 = {s2777[0]};
    assign in6084_2 = {s2778[0]};
    Full_Adder FA_6084(s6084, c6084, in6084_1, in6084_2, s2776[0]);
    wire[0:0] s6085, in6085_1, in6085_2;
    wire c6085;
    assign in6085_1 = {s2780[0]};
    assign in6085_2 = {s2781[0]};
    Full_Adder FA_6085(s6085, c6085, in6085_1, in6085_2, s2779[0]);
    wire[0:0] s6086, in6086_1, in6086_2;
    wire c6086;
    assign in6086_1 = {s2783[0]};
    assign in6086_2 = {s2784[0]};
    Full_Adder FA_6086(s6086, c6086, in6086_1, in6086_2, s2782[0]);
    wire[0:0] s6087, in6087_1, in6087_2;
    wire c6087;
    assign in6087_1 = {s2786[0]};
    assign in6087_2 = {s2787[0]};
    Full_Adder FA_6087(s6087, c6087, in6087_1, in6087_2, s2785[0]);
    wire[0:0] s6088, in6088_1, in6088_2;
    wire c6088;
    assign in6088_1 = {s2789[0]};
    assign in6088_2 = {s2790[0]};
    Full_Adder FA_6088(s6088, c6088, in6088_1, in6088_2, s2788[0]);
    wire[0:0] s6089, in6089_1, in6089_2;
    wire c6089;
    assign in6089_1 = {s2792[0]};
    assign in6089_2 = {s2793[0]};
    Full_Adder FA_6089(s6089, c6089, in6089_1, in6089_2, s2791[0]);
    wire[0:0] s6090, in6090_1, in6090_2;
    wire c6090;
    assign in6090_1 = {s2795[0]};
    assign in6090_2 = {s2796[0]};
    Full_Adder FA_6090(s6090, c6090, in6090_1, in6090_2, s2794[0]);
    wire[0:0] s6091, in6091_1, in6091_2;
    wire c6091;
    assign in6091_1 = {s2798[0]};
    assign in6091_2 = {s2799[0]};
    Full_Adder FA_6091(s6091, c6091, in6091_1, in6091_2, s2797[0]);
    wire[0:0] s6092, in6092_1, in6092_2;
    wire c6092;
    assign in6092_1 = {s253[0]};
    assign in6092_2 = {c2773};
    Full_Adder FA_6092(s6092, c6092, in6092_1, in6092_2, s252[0]);
    wire[0:0] s6093, in6093_1, in6093_2;
    wire c6093;
    assign in6093_1 = {c2775};
    assign in6093_2 = {c2776};
    Full_Adder FA_6093(s6093, c6093, in6093_1, in6093_2, c2774);
    wire[0:0] s6094, in6094_1, in6094_2;
    wire c6094;
    assign in6094_1 = {c2778};
    assign in6094_2 = {c2779};
    Full_Adder FA_6094(s6094, c6094, in6094_1, in6094_2, c2777);
    wire[0:0] s6095, in6095_1, in6095_2;
    wire c6095;
    assign in6095_1 = {c2781};
    assign in6095_2 = {c2782};
    Full_Adder FA_6095(s6095, c6095, in6095_1, in6095_2, c2780);
    wire[0:0] s6096, in6096_1, in6096_2;
    wire c6096;
    assign in6096_1 = {c2784};
    assign in6096_2 = {c2785};
    Full_Adder FA_6096(s6096, c6096, in6096_1, in6096_2, c2783);
    wire[0:0] s6097, in6097_1, in6097_2;
    wire c6097;
    assign in6097_1 = {c2787};
    assign in6097_2 = {c2788};
    Full_Adder FA_6097(s6097, c6097, in6097_1, in6097_2, c2786);
    wire[0:0] s6098, in6098_1, in6098_2;
    wire c6098;
    assign in6098_1 = {c2790};
    assign in6098_2 = {c2791};
    Full_Adder FA_6098(s6098, c6098, in6098_1, in6098_2, c2789);
    wire[0:0] s6099, in6099_1, in6099_2;
    wire c6099;
    assign in6099_1 = {c2793};
    assign in6099_2 = {c2794};
    Full_Adder FA_6099(s6099, c6099, in6099_1, in6099_2, c2792);
    wire[0:0] s6100, in6100_1, in6100_2;
    wire c6100;
    assign in6100_1 = {c2796};
    assign in6100_2 = {c2797};
    Full_Adder FA_6100(s6100, c6100, in6100_1, in6100_2, c2795);
    wire[0:0] s6101, in6101_1, in6101_2;
    wire c6101;
    assign in6101_1 = {c2799};
    assign in6101_2 = {c2800};
    Full_Adder FA_6101(s6101, c6101, in6101_1, in6101_2, c2798);
    wire[0:0] s6102, in6102_1, in6102_2;
    wire c6102;
    assign in6102_1 = {s2802[0]};
    assign in6102_2 = {s2803[0]};
    Full_Adder FA_6102(s6102, c6102, in6102_1, in6102_2, s2801[0]);
    wire[0:0] s6103, in6103_1, in6103_2;
    wire c6103;
    assign in6103_1 = {s2805[0]};
    assign in6103_2 = {s2806[0]};
    Full_Adder FA_6103(s6103, c6103, in6103_1, in6103_2, s2804[0]);
    wire[0:0] s6104, in6104_1, in6104_2;
    wire c6104;
    assign in6104_1 = {s2808[0]};
    assign in6104_2 = {s2809[0]};
    Full_Adder FA_6104(s6104, c6104, in6104_1, in6104_2, s2807[0]);
    wire[0:0] s6105, in6105_1, in6105_2;
    wire c6105;
    assign in6105_1 = {s2811[0]};
    assign in6105_2 = {s2812[0]};
    Full_Adder FA_6105(s6105, c6105, in6105_1, in6105_2, s2810[0]);
    wire[0:0] s6106, in6106_1, in6106_2;
    wire c6106;
    assign in6106_1 = {s2814[0]};
    assign in6106_2 = {s2815[0]};
    Full_Adder FA_6106(s6106, c6106, in6106_1, in6106_2, s2813[0]);
    wire[0:0] s6107, in6107_1, in6107_2;
    wire c6107;
    assign in6107_1 = {s2817[0]};
    assign in6107_2 = {s2818[0]};
    Full_Adder FA_6107(s6107, c6107, in6107_1, in6107_2, s2816[0]);
    wire[0:0] s6108, in6108_1, in6108_2;
    wire c6108;
    assign in6108_1 = {s2820[0]};
    assign in6108_2 = {s2821[0]};
    Full_Adder FA_6108(s6108, c6108, in6108_1, in6108_2, s2819[0]);
    wire[0:0] s6109, in6109_1, in6109_2;
    wire c6109;
    assign in6109_1 = {s2823[0]};
    assign in6109_2 = {s2824[0]};
    Full_Adder FA_6109(s6109, c6109, in6109_1, in6109_2, s2822[0]);
    wire[0:0] s6110, in6110_1, in6110_2;
    wire c6110;
    assign in6110_1 = {s2826[0]};
    assign in6110_2 = {s2827[0]};
    Full_Adder FA_6110(s6110, c6110, in6110_1, in6110_2, s2825[0]);
    wire[0:0] s6111, in6111_1, in6111_2;
    wire c6111;
    assign in6111_1 = {s276[0]};
    assign in6111_2 = {c2801};
    Full_Adder FA_6111(s6111, c6111, in6111_1, in6111_2, s275[0]);
    wire[0:0] s6112, in6112_1, in6112_2;
    wire c6112;
    assign in6112_1 = {c2803};
    assign in6112_2 = {c2804};
    Full_Adder FA_6112(s6112, c6112, in6112_1, in6112_2, c2802);
    wire[0:0] s6113, in6113_1, in6113_2;
    wire c6113;
    assign in6113_1 = {c2806};
    assign in6113_2 = {c2807};
    Full_Adder FA_6113(s6113, c6113, in6113_1, in6113_2, c2805);
    wire[0:0] s6114, in6114_1, in6114_2;
    wire c6114;
    assign in6114_1 = {c2809};
    assign in6114_2 = {c2810};
    Full_Adder FA_6114(s6114, c6114, in6114_1, in6114_2, c2808);
    wire[0:0] s6115, in6115_1, in6115_2;
    wire c6115;
    assign in6115_1 = {c2812};
    assign in6115_2 = {c2813};
    Full_Adder FA_6115(s6115, c6115, in6115_1, in6115_2, c2811);
    wire[0:0] s6116, in6116_1, in6116_2;
    wire c6116;
    assign in6116_1 = {c2815};
    assign in6116_2 = {c2816};
    Full_Adder FA_6116(s6116, c6116, in6116_1, in6116_2, c2814);
    wire[0:0] s6117, in6117_1, in6117_2;
    wire c6117;
    assign in6117_1 = {c2818};
    assign in6117_2 = {c2819};
    Full_Adder FA_6117(s6117, c6117, in6117_1, in6117_2, c2817);
    wire[0:0] s6118, in6118_1, in6118_2;
    wire c6118;
    assign in6118_1 = {c2821};
    assign in6118_2 = {c2822};
    Full_Adder FA_6118(s6118, c6118, in6118_1, in6118_2, c2820);
    wire[0:0] s6119, in6119_1, in6119_2;
    wire c6119;
    assign in6119_1 = {c2824};
    assign in6119_2 = {c2825};
    Full_Adder FA_6119(s6119, c6119, in6119_1, in6119_2, c2823);
    wire[0:0] s6120, in6120_1, in6120_2;
    wire c6120;
    assign in6120_1 = {c2827};
    assign in6120_2 = {c2828};
    Full_Adder FA_6120(s6120, c6120, in6120_1, in6120_2, c2826);
    wire[0:0] s6121, in6121_1, in6121_2;
    wire c6121;
    assign in6121_1 = {s2830[0]};
    assign in6121_2 = {s2831[0]};
    Full_Adder FA_6121(s6121, c6121, in6121_1, in6121_2, s2829[0]);
    wire[0:0] s6122, in6122_1, in6122_2;
    wire c6122;
    assign in6122_1 = {s2833[0]};
    assign in6122_2 = {s2834[0]};
    Full_Adder FA_6122(s6122, c6122, in6122_1, in6122_2, s2832[0]);
    wire[0:0] s6123, in6123_1, in6123_2;
    wire c6123;
    assign in6123_1 = {s2836[0]};
    assign in6123_2 = {s2837[0]};
    Full_Adder FA_6123(s6123, c6123, in6123_1, in6123_2, s2835[0]);
    wire[0:0] s6124, in6124_1, in6124_2;
    wire c6124;
    assign in6124_1 = {s2839[0]};
    assign in6124_2 = {s2840[0]};
    Full_Adder FA_6124(s6124, c6124, in6124_1, in6124_2, s2838[0]);
    wire[0:0] s6125, in6125_1, in6125_2;
    wire c6125;
    assign in6125_1 = {s2842[0]};
    assign in6125_2 = {s2843[0]};
    Full_Adder FA_6125(s6125, c6125, in6125_1, in6125_2, s2841[0]);
    wire[0:0] s6126, in6126_1, in6126_2;
    wire c6126;
    assign in6126_1 = {s2845[0]};
    assign in6126_2 = {s2846[0]};
    Full_Adder FA_6126(s6126, c6126, in6126_1, in6126_2, s2844[0]);
    wire[0:0] s6127, in6127_1, in6127_2;
    wire c6127;
    assign in6127_1 = {s2848[0]};
    assign in6127_2 = {s2849[0]};
    Full_Adder FA_6127(s6127, c6127, in6127_1, in6127_2, s2847[0]);
    wire[0:0] s6128, in6128_1, in6128_2;
    wire c6128;
    assign in6128_1 = {s2851[0]};
    assign in6128_2 = {s2852[0]};
    Full_Adder FA_6128(s6128, c6128, in6128_1, in6128_2, s2850[0]);
    wire[0:0] s6129, in6129_1, in6129_2;
    wire c6129;
    assign in6129_1 = {s2854[0]};
    assign in6129_2 = {s2855[0]};
    Full_Adder FA_6129(s6129, c6129, in6129_1, in6129_2, s2853[0]);
    wire[0:0] s6130, in6130_1, in6130_2;
    wire c6130;
    assign in6130_1 = {s300[0]};
    assign in6130_2 = {c2829};
    Full_Adder FA_6130(s6130, c6130, in6130_1, in6130_2, s299[0]);
    wire[0:0] s6131, in6131_1, in6131_2;
    wire c6131;
    assign in6131_1 = {c2831};
    assign in6131_2 = {c2832};
    Full_Adder FA_6131(s6131, c6131, in6131_1, in6131_2, c2830);
    wire[0:0] s6132, in6132_1, in6132_2;
    wire c6132;
    assign in6132_1 = {c2834};
    assign in6132_2 = {c2835};
    Full_Adder FA_6132(s6132, c6132, in6132_1, in6132_2, c2833);
    wire[0:0] s6133, in6133_1, in6133_2;
    wire c6133;
    assign in6133_1 = {c2837};
    assign in6133_2 = {c2838};
    Full_Adder FA_6133(s6133, c6133, in6133_1, in6133_2, c2836);
    wire[0:0] s6134, in6134_1, in6134_2;
    wire c6134;
    assign in6134_1 = {c2840};
    assign in6134_2 = {c2841};
    Full_Adder FA_6134(s6134, c6134, in6134_1, in6134_2, c2839);
    wire[0:0] s6135, in6135_1, in6135_2;
    wire c6135;
    assign in6135_1 = {c2843};
    assign in6135_2 = {c2844};
    Full_Adder FA_6135(s6135, c6135, in6135_1, in6135_2, c2842);
    wire[0:0] s6136, in6136_1, in6136_2;
    wire c6136;
    assign in6136_1 = {c2846};
    assign in6136_2 = {c2847};
    Full_Adder FA_6136(s6136, c6136, in6136_1, in6136_2, c2845);
    wire[0:0] s6137, in6137_1, in6137_2;
    wire c6137;
    assign in6137_1 = {c2849};
    assign in6137_2 = {c2850};
    Full_Adder FA_6137(s6137, c6137, in6137_1, in6137_2, c2848);
    wire[0:0] s6138, in6138_1, in6138_2;
    wire c6138;
    assign in6138_1 = {c2852};
    assign in6138_2 = {c2853};
    Full_Adder FA_6138(s6138, c6138, in6138_1, in6138_2, c2851);
    wire[0:0] s6139, in6139_1, in6139_2;
    wire c6139;
    assign in6139_1 = {c2855};
    assign in6139_2 = {c2856};
    Full_Adder FA_6139(s6139, c6139, in6139_1, in6139_2, c2854);
    wire[0:0] s6140, in6140_1, in6140_2;
    wire c6140;
    assign in6140_1 = {s2858[0]};
    assign in6140_2 = {s2859[0]};
    Full_Adder FA_6140(s6140, c6140, in6140_1, in6140_2, s2857[0]);
    wire[0:0] s6141, in6141_1, in6141_2;
    wire c6141;
    assign in6141_1 = {s2861[0]};
    assign in6141_2 = {s2862[0]};
    Full_Adder FA_6141(s6141, c6141, in6141_1, in6141_2, s2860[0]);
    wire[0:0] s6142, in6142_1, in6142_2;
    wire c6142;
    assign in6142_1 = {s2864[0]};
    assign in6142_2 = {s2865[0]};
    Full_Adder FA_6142(s6142, c6142, in6142_1, in6142_2, s2863[0]);
    wire[0:0] s6143, in6143_1, in6143_2;
    wire c6143;
    assign in6143_1 = {s2867[0]};
    assign in6143_2 = {s2868[0]};
    Full_Adder FA_6143(s6143, c6143, in6143_1, in6143_2, s2866[0]);
    wire[0:0] s6144, in6144_1, in6144_2;
    wire c6144;
    assign in6144_1 = {s2870[0]};
    assign in6144_2 = {s2871[0]};
    Full_Adder FA_6144(s6144, c6144, in6144_1, in6144_2, s2869[0]);
    wire[0:0] s6145, in6145_1, in6145_2;
    wire c6145;
    assign in6145_1 = {s2873[0]};
    assign in6145_2 = {s2874[0]};
    Full_Adder FA_6145(s6145, c6145, in6145_1, in6145_2, s2872[0]);
    wire[0:0] s6146, in6146_1, in6146_2;
    wire c6146;
    assign in6146_1 = {s2876[0]};
    assign in6146_2 = {s2877[0]};
    Full_Adder FA_6146(s6146, c6146, in6146_1, in6146_2, s2875[0]);
    wire[0:0] s6147, in6147_1, in6147_2;
    wire c6147;
    assign in6147_1 = {s2879[0]};
    assign in6147_2 = {s2880[0]};
    Full_Adder FA_6147(s6147, c6147, in6147_1, in6147_2, s2878[0]);
    wire[0:0] s6148, in6148_1, in6148_2;
    wire c6148;
    assign in6148_1 = {s2882[0]};
    assign in6148_2 = {s2883[0]};
    Full_Adder FA_6148(s6148, c6148, in6148_1, in6148_2, s2881[0]);
    wire[0:0] s6149, in6149_1, in6149_2;
    wire c6149;
    assign in6149_1 = {s325[0]};
    assign in6149_2 = {c2857};
    Full_Adder FA_6149(s6149, c6149, in6149_1, in6149_2, s324[0]);
    wire[0:0] s6150, in6150_1, in6150_2;
    wire c6150;
    assign in6150_1 = {c2859};
    assign in6150_2 = {c2860};
    Full_Adder FA_6150(s6150, c6150, in6150_1, in6150_2, c2858);
    wire[0:0] s6151, in6151_1, in6151_2;
    wire c6151;
    assign in6151_1 = {c2862};
    assign in6151_2 = {c2863};
    Full_Adder FA_6151(s6151, c6151, in6151_1, in6151_2, c2861);
    wire[0:0] s6152, in6152_1, in6152_2;
    wire c6152;
    assign in6152_1 = {c2865};
    assign in6152_2 = {c2866};
    Full_Adder FA_6152(s6152, c6152, in6152_1, in6152_2, c2864);
    wire[0:0] s6153, in6153_1, in6153_2;
    wire c6153;
    assign in6153_1 = {c2868};
    assign in6153_2 = {c2869};
    Full_Adder FA_6153(s6153, c6153, in6153_1, in6153_2, c2867);
    wire[0:0] s6154, in6154_1, in6154_2;
    wire c6154;
    assign in6154_1 = {c2871};
    assign in6154_2 = {c2872};
    Full_Adder FA_6154(s6154, c6154, in6154_1, in6154_2, c2870);
    wire[0:0] s6155, in6155_1, in6155_2;
    wire c6155;
    assign in6155_1 = {c2874};
    assign in6155_2 = {c2875};
    Full_Adder FA_6155(s6155, c6155, in6155_1, in6155_2, c2873);
    wire[0:0] s6156, in6156_1, in6156_2;
    wire c6156;
    assign in6156_1 = {c2877};
    assign in6156_2 = {c2878};
    Full_Adder FA_6156(s6156, c6156, in6156_1, in6156_2, c2876);
    wire[0:0] s6157, in6157_1, in6157_2;
    wire c6157;
    assign in6157_1 = {c2880};
    assign in6157_2 = {c2881};
    Full_Adder FA_6157(s6157, c6157, in6157_1, in6157_2, c2879);
    wire[0:0] s6158, in6158_1, in6158_2;
    wire c6158;
    assign in6158_1 = {c2883};
    assign in6158_2 = {c2884};
    Full_Adder FA_6158(s6158, c6158, in6158_1, in6158_2, c2882);
    wire[0:0] s6159, in6159_1, in6159_2;
    wire c6159;
    assign in6159_1 = {s2886[0]};
    assign in6159_2 = {s2887[0]};
    Full_Adder FA_6159(s6159, c6159, in6159_1, in6159_2, s2885[0]);
    wire[0:0] s6160, in6160_1, in6160_2;
    wire c6160;
    assign in6160_1 = {s2889[0]};
    assign in6160_2 = {s2890[0]};
    Full_Adder FA_6160(s6160, c6160, in6160_1, in6160_2, s2888[0]);
    wire[0:0] s6161, in6161_1, in6161_2;
    wire c6161;
    assign in6161_1 = {s2892[0]};
    assign in6161_2 = {s2893[0]};
    Full_Adder FA_6161(s6161, c6161, in6161_1, in6161_2, s2891[0]);
    wire[0:0] s6162, in6162_1, in6162_2;
    wire c6162;
    assign in6162_1 = {s2895[0]};
    assign in6162_2 = {s2896[0]};
    Full_Adder FA_6162(s6162, c6162, in6162_1, in6162_2, s2894[0]);
    wire[0:0] s6163, in6163_1, in6163_2;
    wire c6163;
    assign in6163_1 = {s2898[0]};
    assign in6163_2 = {s2899[0]};
    Full_Adder FA_6163(s6163, c6163, in6163_1, in6163_2, s2897[0]);
    wire[0:0] s6164, in6164_1, in6164_2;
    wire c6164;
    assign in6164_1 = {s2901[0]};
    assign in6164_2 = {s2902[0]};
    Full_Adder FA_6164(s6164, c6164, in6164_1, in6164_2, s2900[0]);
    wire[0:0] s6165, in6165_1, in6165_2;
    wire c6165;
    assign in6165_1 = {s2904[0]};
    assign in6165_2 = {s2905[0]};
    Full_Adder FA_6165(s6165, c6165, in6165_1, in6165_2, s2903[0]);
    wire[0:0] s6166, in6166_1, in6166_2;
    wire c6166;
    assign in6166_1 = {s2907[0]};
    assign in6166_2 = {s2908[0]};
    Full_Adder FA_6166(s6166, c6166, in6166_1, in6166_2, s2906[0]);
    wire[0:0] s6167, in6167_1, in6167_2;
    wire c6167;
    assign in6167_1 = {s2910[0]};
    assign in6167_2 = {s2911[0]};
    Full_Adder FA_6167(s6167, c6167, in6167_1, in6167_2, s2909[0]);
    wire[0:0] s6168, in6168_1, in6168_2;
    wire c6168;
    assign in6168_1 = {s351[0]};
    assign in6168_2 = {c2885};
    Full_Adder FA_6168(s6168, c6168, in6168_1, in6168_2, s350[0]);
    wire[0:0] s6169, in6169_1, in6169_2;
    wire c6169;
    assign in6169_1 = {c2887};
    assign in6169_2 = {c2888};
    Full_Adder FA_6169(s6169, c6169, in6169_1, in6169_2, c2886);
    wire[0:0] s6170, in6170_1, in6170_2;
    wire c6170;
    assign in6170_1 = {c2890};
    assign in6170_2 = {c2891};
    Full_Adder FA_6170(s6170, c6170, in6170_1, in6170_2, c2889);
    wire[0:0] s6171, in6171_1, in6171_2;
    wire c6171;
    assign in6171_1 = {c2893};
    assign in6171_2 = {c2894};
    Full_Adder FA_6171(s6171, c6171, in6171_1, in6171_2, c2892);
    wire[0:0] s6172, in6172_1, in6172_2;
    wire c6172;
    assign in6172_1 = {c2896};
    assign in6172_2 = {c2897};
    Full_Adder FA_6172(s6172, c6172, in6172_1, in6172_2, c2895);
    wire[0:0] s6173, in6173_1, in6173_2;
    wire c6173;
    assign in6173_1 = {c2899};
    assign in6173_2 = {c2900};
    Full_Adder FA_6173(s6173, c6173, in6173_1, in6173_2, c2898);
    wire[0:0] s6174, in6174_1, in6174_2;
    wire c6174;
    assign in6174_1 = {c2902};
    assign in6174_2 = {c2903};
    Full_Adder FA_6174(s6174, c6174, in6174_1, in6174_2, c2901);
    wire[0:0] s6175, in6175_1, in6175_2;
    wire c6175;
    assign in6175_1 = {c2905};
    assign in6175_2 = {c2906};
    Full_Adder FA_6175(s6175, c6175, in6175_1, in6175_2, c2904);
    wire[0:0] s6176, in6176_1, in6176_2;
    wire c6176;
    assign in6176_1 = {c2908};
    assign in6176_2 = {c2909};
    Full_Adder FA_6176(s6176, c6176, in6176_1, in6176_2, c2907);
    wire[0:0] s6177, in6177_1, in6177_2;
    wire c6177;
    assign in6177_1 = {c2911};
    assign in6177_2 = {c2912};
    Full_Adder FA_6177(s6177, c6177, in6177_1, in6177_2, c2910);
    wire[0:0] s6178, in6178_1, in6178_2;
    wire c6178;
    assign in6178_1 = {s2914[0]};
    assign in6178_2 = {s2915[0]};
    Full_Adder FA_6178(s6178, c6178, in6178_1, in6178_2, s2913[0]);
    wire[0:0] s6179, in6179_1, in6179_2;
    wire c6179;
    assign in6179_1 = {s2917[0]};
    assign in6179_2 = {s2918[0]};
    Full_Adder FA_6179(s6179, c6179, in6179_1, in6179_2, s2916[0]);
    wire[0:0] s6180, in6180_1, in6180_2;
    wire c6180;
    assign in6180_1 = {s2920[0]};
    assign in6180_2 = {s2921[0]};
    Full_Adder FA_6180(s6180, c6180, in6180_1, in6180_2, s2919[0]);
    wire[0:0] s6181, in6181_1, in6181_2;
    wire c6181;
    assign in6181_1 = {s2923[0]};
    assign in6181_2 = {s2924[0]};
    Full_Adder FA_6181(s6181, c6181, in6181_1, in6181_2, s2922[0]);
    wire[0:0] s6182, in6182_1, in6182_2;
    wire c6182;
    assign in6182_1 = {s2926[0]};
    assign in6182_2 = {s2927[0]};
    Full_Adder FA_6182(s6182, c6182, in6182_1, in6182_2, s2925[0]);
    wire[0:0] s6183, in6183_1, in6183_2;
    wire c6183;
    assign in6183_1 = {s2929[0]};
    assign in6183_2 = {s2930[0]};
    Full_Adder FA_6183(s6183, c6183, in6183_1, in6183_2, s2928[0]);
    wire[0:0] s6184, in6184_1, in6184_2;
    wire c6184;
    assign in6184_1 = {s2932[0]};
    assign in6184_2 = {s2933[0]};
    Full_Adder FA_6184(s6184, c6184, in6184_1, in6184_2, s2931[0]);
    wire[0:0] s6185, in6185_1, in6185_2;
    wire c6185;
    assign in6185_1 = {s2935[0]};
    assign in6185_2 = {s2936[0]};
    Full_Adder FA_6185(s6185, c6185, in6185_1, in6185_2, s2934[0]);
    wire[0:0] s6186, in6186_1, in6186_2;
    wire c6186;
    assign in6186_1 = {s2938[0]};
    assign in6186_2 = {s2939[0]};
    Full_Adder FA_6186(s6186, c6186, in6186_1, in6186_2, s2937[0]);
    wire[0:0] s6187, in6187_1, in6187_2;
    wire c6187;
    assign in6187_1 = {s378[0]};
    assign in6187_2 = {c2913};
    Full_Adder FA_6187(s6187, c6187, in6187_1, in6187_2, s377[0]);
    wire[0:0] s6188, in6188_1, in6188_2;
    wire c6188;
    assign in6188_1 = {c2915};
    assign in6188_2 = {c2916};
    Full_Adder FA_6188(s6188, c6188, in6188_1, in6188_2, c2914);
    wire[0:0] s6189, in6189_1, in6189_2;
    wire c6189;
    assign in6189_1 = {c2918};
    assign in6189_2 = {c2919};
    Full_Adder FA_6189(s6189, c6189, in6189_1, in6189_2, c2917);
    wire[0:0] s6190, in6190_1, in6190_2;
    wire c6190;
    assign in6190_1 = {c2921};
    assign in6190_2 = {c2922};
    Full_Adder FA_6190(s6190, c6190, in6190_1, in6190_2, c2920);
    wire[0:0] s6191, in6191_1, in6191_2;
    wire c6191;
    assign in6191_1 = {c2924};
    assign in6191_2 = {c2925};
    Full_Adder FA_6191(s6191, c6191, in6191_1, in6191_2, c2923);
    wire[0:0] s6192, in6192_1, in6192_2;
    wire c6192;
    assign in6192_1 = {c2927};
    assign in6192_2 = {c2928};
    Full_Adder FA_6192(s6192, c6192, in6192_1, in6192_2, c2926);
    wire[0:0] s6193, in6193_1, in6193_2;
    wire c6193;
    assign in6193_1 = {c2930};
    assign in6193_2 = {c2931};
    Full_Adder FA_6193(s6193, c6193, in6193_1, in6193_2, c2929);
    wire[0:0] s6194, in6194_1, in6194_2;
    wire c6194;
    assign in6194_1 = {c2933};
    assign in6194_2 = {c2934};
    Full_Adder FA_6194(s6194, c6194, in6194_1, in6194_2, c2932);
    wire[0:0] s6195, in6195_1, in6195_2;
    wire c6195;
    assign in6195_1 = {c2936};
    assign in6195_2 = {c2937};
    Full_Adder FA_6195(s6195, c6195, in6195_1, in6195_2, c2935);
    wire[0:0] s6196, in6196_1, in6196_2;
    wire c6196;
    assign in6196_1 = {c2939};
    assign in6196_2 = {c2940};
    Full_Adder FA_6196(s6196, c6196, in6196_1, in6196_2, c2938);
    wire[0:0] s6197, in6197_1, in6197_2;
    wire c6197;
    assign in6197_1 = {s2942[0]};
    assign in6197_2 = {s2943[0]};
    Full_Adder FA_6197(s6197, c6197, in6197_1, in6197_2, s2941[0]);
    wire[0:0] s6198, in6198_1, in6198_2;
    wire c6198;
    assign in6198_1 = {s2945[0]};
    assign in6198_2 = {s2946[0]};
    Full_Adder FA_6198(s6198, c6198, in6198_1, in6198_2, s2944[0]);
    wire[0:0] s6199, in6199_1, in6199_2;
    wire c6199;
    assign in6199_1 = {s2948[0]};
    assign in6199_2 = {s2949[0]};
    Full_Adder FA_6199(s6199, c6199, in6199_1, in6199_2, s2947[0]);
    wire[0:0] s6200, in6200_1, in6200_2;
    wire c6200;
    assign in6200_1 = {s2951[0]};
    assign in6200_2 = {s2952[0]};
    Full_Adder FA_6200(s6200, c6200, in6200_1, in6200_2, s2950[0]);
    wire[0:0] s6201, in6201_1, in6201_2;
    wire c6201;
    assign in6201_1 = {s2954[0]};
    assign in6201_2 = {s2955[0]};
    Full_Adder FA_6201(s6201, c6201, in6201_1, in6201_2, s2953[0]);
    wire[0:0] s6202, in6202_1, in6202_2;
    wire c6202;
    assign in6202_1 = {s2957[0]};
    assign in6202_2 = {s2958[0]};
    Full_Adder FA_6202(s6202, c6202, in6202_1, in6202_2, s2956[0]);
    wire[0:0] s6203, in6203_1, in6203_2;
    wire c6203;
    assign in6203_1 = {s2960[0]};
    assign in6203_2 = {s2961[0]};
    Full_Adder FA_6203(s6203, c6203, in6203_1, in6203_2, s2959[0]);
    wire[0:0] s6204, in6204_1, in6204_2;
    wire c6204;
    assign in6204_1 = {s2963[0]};
    assign in6204_2 = {s2964[0]};
    Full_Adder FA_6204(s6204, c6204, in6204_1, in6204_2, s2962[0]);
    wire[0:0] s6205, in6205_1, in6205_2;
    wire c6205;
    assign in6205_1 = {s2966[0]};
    assign in6205_2 = {s2967[0]};
    Full_Adder FA_6205(s6205, c6205, in6205_1, in6205_2, s2965[0]);
    wire[0:0] s6206, in6206_1, in6206_2;
    wire c6206;
    assign in6206_1 = {s406[0]};
    assign in6206_2 = {c2941};
    Full_Adder FA_6206(s6206, c6206, in6206_1, in6206_2, s405[0]);
    wire[0:0] s6207, in6207_1, in6207_2;
    wire c6207;
    assign in6207_1 = {c2943};
    assign in6207_2 = {c2944};
    Full_Adder FA_6207(s6207, c6207, in6207_1, in6207_2, c2942);
    wire[0:0] s6208, in6208_1, in6208_2;
    wire c6208;
    assign in6208_1 = {c2946};
    assign in6208_2 = {c2947};
    Full_Adder FA_6208(s6208, c6208, in6208_1, in6208_2, c2945);
    wire[0:0] s6209, in6209_1, in6209_2;
    wire c6209;
    assign in6209_1 = {c2949};
    assign in6209_2 = {c2950};
    Full_Adder FA_6209(s6209, c6209, in6209_1, in6209_2, c2948);
    wire[0:0] s6210, in6210_1, in6210_2;
    wire c6210;
    assign in6210_1 = {c2952};
    assign in6210_2 = {c2953};
    Full_Adder FA_6210(s6210, c6210, in6210_1, in6210_2, c2951);
    wire[0:0] s6211, in6211_1, in6211_2;
    wire c6211;
    assign in6211_1 = {c2955};
    assign in6211_2 = {c2956};
    Full_Adder FA_6211(s6211, c6211, in6211_1, in6211_2, c2954);
    wire[0:0] s6212, in6212_1, in6212_2;
    wire c6212;
    assign in6212_1 = {c2958};
    assign in6212_2 = {c2959};
    Full_Adder FA_6212(s6212, c6212, in6212_1, in6212_2, c2957);
    wire[0:0] s6213, in6213_1, in6213_2;
    wire c6213;
    assign in6213_1 = {c2961};
    assign in6213_2 = {c2962};
    Full_Adder FA_6213(s6213, c6213, in6213_1, in6213_2, c2960);
    wire[0:0] s6214, in6214_1, in6214_2;
    wire c6214;
    assign in6214_1 = {c2964};
    assign in6214_2 = {c2965};
    Full_Adder FA_6214(s6214, c6214, in6214_1, in6214_2, c2963);
    wire[0:0] s6215, in6215_1, in6215_2;
    wire c6215;
    assign in6215_1 = {c2967};
    assign in6215_2 = {c2968};
    Full_Adder FA_6215(s6215, c6215, in6215_1, in6215_2, c2966);
    wire[0:0] s6216, in6216_1, in6216_2;
    wire c6216;
    assign in6216_1 = {s2970[0]};
    assign in6216_2 = {s2971[0]};
    Full_Adder FA_6216(s6216, c6216, in6216_1, in6216_2, s2969[0]);
    wire[0:0] s6217, in6217_1, in6217_2;
    wire c6217;
    assign in6217_1 = {s2973[0]};
    assign in6217_2 = {s2974[0]};
    Full_Adder FA_6217(s6217, c6217, in6217_1, in6217_2, s2972[0]);
    wire[0:0] s6218, in6218_1, in6218_2;
    wire c6218;
    assign in6218_1 = {s2976[0]};
    assign in6218_2 = {s2977[0]};
    Full_Adder FA_6218(s6218, c6218, in6218_1, in6218_2, s2975[0]);
    wire[0:0] s6219, in6219_1, in6219_2;
    wire c6219;
    assign in6219_1 = {s2979[0]};
    assign in6219_2 = {s2980[0]};
    Full_Adder FA_6219(s6219, c6219, in6219_1, in6219_2, s2978[0]);
    wire[0:0] s6220, in6220_1, in6220_2;
    wire c6220;
    assign in6220_1 = {s2982[0]};
    assign in6220_2 = {s2983[0]};
    Full_Adder FA_6220(s6220, c6220, in6220_1, in6220_2, s2981[0]);
    wire[0:0] s6221, in6221_1, in6221_2;
    wire c6221;
    assign in6221_1 = {s2985[0]};
    assign in6221_2 = {s2986[0]};
    Full_Adder FA_6221(s6221, c6221, in6221_1, in6221_2, s2984[0]);
    wire[0:0] s6222, in6222_1, in6222_2;
    wire c6222;
    assign in6222_1 = {s2988[0]};
    assign in6222_2 = {s2989[0]};
    Full_Adder FA_6222(s6222, c6222, in6222_1, in6222_2, s2987[0]);
    wire[0:0] s6223, in6223_1, in6223_2;
    wire c6223;
    assign in6223_1 = {s2991[0]};
    assign in6223_2 = {s2992[0]};
    Full_Adder FA_6223(s6223, c6223, in6223_1, in6223_2, s2990[0]);
    wire[0:0] s6224, in6224_1, in6224_2;
    wire c6224;
    assign in6224_1 = {s2994[0]};
    assign in6224_2 = {s2995[0]};
    Full_Adder FA_6224(s6224, c6224, in6224_1, in6224_2, s2993[0]);
    wire[0:0] s6225, in6225_1, in6225_2;
    wire c6225;
    assign in6225_1 = {s435[0]};
    assign in6225_2 = {c2969};
    Full_Adder FA_6225(s6225, c6225, in6225_1, in6225_2, s434[0]);
    wire[0:0] s6226, in6226_1, in6226_2;
    wire c6226;
    assign in6226_1 = {c2971};
    assign in6226_2 = {c2972};
    Full_Adder FA_6226(s6226, c6226, in6226_1, in6226_2, c2970);
    wire[0:0] s6227, in6227_1, in6227_2;
    wire c6227;
    assign in6227_1 = {c2974};
    assign in6227_2 = {c2975};
    Full_Adder FA_6227(s6227, c6227, in6227_1, in6227_2, c2973);
    wire[0:0] s6228, in6228_1, in6228_2;
    wire c6228;
    assign in6228_1 = {c2977};
    assign in6228_2 = {c2978};
    Full_Adder FA_6228(s6228, c6228, in6228_1, in6228_2, c2976);
    wire[0:0] s6229, in6229_1, in6229_2;
    wire c6229;
    assign in6229_1 = {c2980};
    assign in6229_2 = {c2981};
    Full_Adder FA_6229(s6229, c6229, in6229_1, in6229_2, c2979);
    wire[0:0] s6230, in6230_1, in6230_2;
    wire c6230;
    assign in6230_1 = {c2983};
    assign in6230_2 = {c2984};
    Full_Adder FA_6230(s6230, c6230, in6230_1, in6230_2, c2982);
    wire[0:0] s6231, in6231_1, in6231_2;
    wire c6231;
    assign in6231_1 = {c2986};
    assign in6231_2 = {c2987};
    Full_Adder FA_6231(s6231, c6231, in6231_1, in6231_2, c2985);
    wire[0:0] s6232, in6232_1, in6232_2;
    wire c6232;
    assign in6232_1 = {c2989};
    assign in6232_2 = {c2990};
    Full_Adder FA_6232(s6232, c6232, in6232_1, in6232_2, c2988);
    wire[0:0] s6233, in6233_1, in6233_2;
    wire c6233;
    assign in6233_1 = {c2992};
    assign in6233_2 = {c2993};
    Full_Adder FA_6233(s6233, c6233, in6233_1, in6233_2, c2991);
    wire[0:0] s6234, in6234_1, in6234_2;
    wire c6234;
    assign in6234_1 = {c2995};
    assign in6234_2 = {c2996};
    Full_Adder FA_6234(s6234, c6234, in6234_1, in6234_2, c2994);
    wire[0:0] s6235, in6235_1, in6235_2;
    wire c6235;
    assign in6235_1 = {s2998[0]};
    assign in6235_2 = {s2999[0]};
    Full_Adder FA_6235(s6235, c6235, in6235_1, in6235_2, s2997[0]);
    wire[0:0] s6236, in6236_1, in6236_2;
    wire c6236;
    assign in6236_1 = {s3001[0]};
    assign in6236_2 = {s3002[0]};
    Full_Adder FA_6236(s6236, c6236, in6236_1, in6236_2, s3000[0]);
    wire[0:0] s6237, in6237_1, in6237_2;
    wire c6237;
    assign in6237_1 = {s3004[0]};
    assign in6237_2 = {s3005[0]};
    Full_Adder FA_6237(s6237, c6237, in6237_1, in6237_2, s3003[0]);
    wire[0:0] s6238, in6238_1, in6238_2;
    wire c6238;
    assign in6238_1 = {s3007[0]};
    assign in6238_2 = {s3008[0]};
    Full_Adder FA_6238(s6238, c6238, in6238_1, in6238_2, s3006[0]);
    wire[0:0] s6239, in6239_1, in6239_2;
    wire c6239;
    assign in6239_1 = {s3010[0]};
    assign in6239_2 = {s3011[0]};
    Full_Adder FA_6239(s6239, c6239, in6239_1, in6239_2, s3009[0]);
    wire[0:0] s6240, in6240_1, in6240_2;
    wire c6240;
    assign in6240_1 = {s3013[0]};
    assign in6240_2 = {s3014[0]};
    Full_Adder FA_6240(s6240, c6240, in6240_1, in6240_2, s3012[0]);
    wire[0:0] s6241, in6241_1, in6241_2;
    wire c6241;
    assign in6241_1 = {s3016[0]};
    assign in6241_2 = {s3017[0]};
    Full_Adder FA_6241(s6241, c6241, in6241_1, in6241_2, s3015[0]);
    wire[0:0] s6242, in6242_1, in6242_2;
    wire c6242;
    assign in6242_1 = {s3019[0]};
    assign in6242_2 = {s3020[0]};
    Full_Adder FA_6242(s6242, c6242, in6242_1, in6242_2, s3018[0]);
    wire[0:0] s6243, in6243_1, in6243_2;
    wire c6243;
    assign in6243_1 = {s3022[0]};
    assign in6243_2 = {s3023[0]};
    Full_Adder FA_6243(s6243, c6243, in6243_1, in6243_2, s3021[0]);
    wire[0:0] s6244, in6244_1, in6244_2;
    wire c6244;
    assign in6244_1 = {s465[0]};
    assign in6244_2 = {c2997};
    Full_Adder FA_6244(s6244, c6244, in6244_1, in6244_2, s464[0]);
    wire[0:0] s6245, in6245_1, in6245_2;
    wire c6245;
    assign in6245_1 = {c2999};
    assign in6245_2 = {c3000};
    Full_Adder FA_6245(s6245, c6245, in6245_1, in6245_2, c2998);
    wire[0:0] s6246, in6246_1, in6246_2;
    wire c6246;
    assign in6246_1 = {c3002};
    assign in6246_2 = {c3003};
    Full_Adder FA_6246(s6246, c6246, in6246_1, in6246_2, c3001);
    wire[0:0] s6247, in6247_1, in6247_2;
    wire c6247;
    assign in6247_1 = {c3005};
    assign in6247_2 = {c3006};
    Full_Adder FA_6247(s6247, c6247, in6247_1, in6247_2, c3004);
    wire[0:0] s6248, in6248_1, in6248_2;
    wire c6248;
    assign in6248_1 = {c3008};
    assign in6248_2 = {c3009};
    Full_Adder FA_6248(s6248, c6248, in6248_1, in6248_2, c3007);
    wire[0:0] s6249, in6249_1, in6249_2;
    wire c6249;
    assign in6249_1 = {c3011};
    assign in6249_2 = {c3012};
    Full_Adder FA_6249(s6249, c6249, in6249_1, in6249_2, c3010);
    wire[0:0] s6250, in6250_1, in6250_2;
    wire c6250;
    assign in6250_1 = {c3014};
    assign in6250_2 = {c3015};
    Full_Adder FA_6250(s6250, c6250, in6250_1, in6250_2, c3013);
    wire[0:0] s6251, in6251_1, in6251_2;
    wire c6251;
    assign in6251_1 = {c3017};
    assign in6251_2 = {c3018};
    Full_Adder FA_6251(s6251, c6251, in6251_1, in6251_2, c3016);
    wire[0:0] s6252, in6252_1, in6252_2;
    wire c6252;
    assign in6252_1 = {c3020};
    assign in6252_2 = {c3021};
    Full_Adder FA_6252(s6252, c6252, in6252_1, in6252_2, c3019);
    wire[0:0] s6253, in6253_1, in6253_2;
    wire c6253;
    assign in6253_1 = {c3023};
    assign in6253_2 = {c3024};
    Full_Adder FA_6253(s6253, c6253, in6253_1, in6253_2, c3022);
    wire[0:0] s6254, in6254_1, in6254_2;
    wire c6254;
    assign in6254_1 = {s3026[0]};
    assign in6254_2 = {s3027[0]};
    Full_Adder FA_6254(s6254, c6254, in6254_1, in6254_2, s3025[0]);
    wire[0:0] s6255, in6255_1, in6255_2;
    wire c6255;
    assign in6255_1 = {s3029[0]};
    assign in6255_2 = {s3030[0]};
    Full_Adder FA_6255(s6255, c6255, in6255_1, in6255_2, s3028[0]);
    wire[0:0] s6256, in6256_1, in6256_2;
    wire c6256;
    assign in6256_1 = {s3032[0]};
    assign in6256_2 = {s3033[0]};
    Full_Adder FA_6256(s6256, c6256, in6256_1, in6256_2, s3031[0]);
    wire[0:0] s6257, in6257_1, in6257_2;
    wire c6257;
    assign in6257_1 = {s3035[0]};
    assign in6257_2 = {s3036[0]};
    Full_Adder FA_6257(s6257, c6257, in6257_1, in6257_2, s3034[0]);
    wire[0:0] s6258, in6258_1, in6258_2;
    wire c6258;
    assign in6258_1 = {s3038[0]};
    assign in6258_2 = {s3039[0]};
    Full_Adder FA_6258(s6258, c6258, in6258_1, in6258_2, s3037[0]);
    wire[0:0] s6259, in6259_1, in6259_2;
    wire c6259;
    assign in6259_1 = {s3041[0]};
    assign in6259_2 = {s3042[0]};
    Full_Adder FA_6259(s6259, c6259, in6259_1, in6259_2, s3040[0]);
    wire[0:0] s6260, in6260_1, in6260_2;
    wire c6260;
    assign in6260_1 = {s3044[0]};
    assign in6260_2 = {s3045[0]};
    Full_Adder FA_6260(s6260, c6260, in6260_1, in6260_2, s3043[0]);
    wire[0:0] s6261, in6261_1, in6261_2;
    wire c6261;
    assign in6261_1 = {s3047[0]};
    assign in6261_2 = {s3048[0]};
    Full_Adder FA_6261(s6261, c6261, in6261_1, in6261_2, s3046[0]);
    wire[0:0] s6262, in6262_1, in6262_2;
    wire c6262;
    assign in6262_1 = {s3050[0]};
    assign in6262_2 = {s3051[0]};
    Full_Adder FA_6262(s6262, c6262, in6262_1, in6262_2, s3049[0]);
    wire[0:0] s6263, in6263_1, in6263_2;
    wire c6263;
    assign in6263_1 = {s496[0]};
    assign in6263_2 = {c3025};
    Full_Adder FA_6263(s6263, c6263, in6263_1, in6263_2, s495[0]);
    wire[0:0] s6264, in6264_1, in6264_2;
    wire c6264;
    assign in6264_1 = {c3027};
    assign in6264_2 = {c3028};
    Full_Adder FA_6264(s6264, c6264, in6264_1, in6264_2, c3026);
    wire[0:0] s6265, in6265_1, in6265_2;
    wire c6265;
    assign in6265_1 = {c3030};
    assign in6265_2 = {c3031};
    Full_Adder FA_6265(s6265, c6265, in6265_1, in6265_2, c3029);
    wire[0:0] s6266, in6266_1, in6266_2;
    wire c6266;
    assign in6266_1 = {c3033};
    assign in6266_2 = {c3034};
    Full_Adder FA_6266(s6266, c6266, in6266_1, in6266_2, c3032);
    wire[0:0] s6267, in6267_1, in6267_2;
    wire c6267;
    assign in6267_1 = {c3036};
    assign in6267_2 = {c3037};
    Full_Adder FA_6267(s6267, c6267, in6267_1, in6267_2, c3035);
    wire[0:0] s6268, in6268_1, in6268_2;
    wire c6268;
    assign in6268_1 = {c3039};
    assign in6268_2 = {c3040};
    Full_Adder FA_6268(s6268, c6268, in6268_1, in6268_2, c3038);
    wire[0:0] s6269, in6269_1, in6269_2;
    wire c6269;
    assign in6269_1 = {c3042};
    assign in6269_2 = {c3043};
    Full_Adder FA_6269(s6269, c6269, in6269_1, in6269_2, c3041);
    wire[0:0] s6270, in6270_1, in6270_2;
    wire c6270;
    assign in6270_1 = {c3045};
    assign in6270_2 = {c3046};
    Full_Adder FA_6270(s6270, c6270, in6270_1, in6270_2, c3044);
    wire[0:0] s6271, in6271_1, in6271_2;
    wire c6271;
    assign in6271_1 = {c3048};
    assign in6271_2 = {c3049};
    Full_Adder FA_6271(s6271, c6271, in6271_1, in6271_2, c3047);
    wire[0:0] s6272, in6272_1, in6272_2;
    wire c6272;
    assign in6272_1 = {c3051};
    assign in6272_2 = {c3052};
    Full_Adder FA_6272(s6272, c6272, in6272_1, in6272_2, c3050);
    wire[0:0] s6273, in6273_1, in6273_2;
    wire c6273;
    assign in6273_1 = {s3054[0]};
    assign in6273_2 = {s3055[0]};
    Full_Adder FA_6273(s6273, c6273, in6273_1, in6273_2, s3053[0]);
    wire[0:0] s6274, in6274_1, in6274_2;
    wire c6274;
    assign in6274_1 = {s3057[0]};
    assign in6274_2 = {s3058[0]};
    Full_Adder FA_6274(s6274, c6274, in6274_1, in6274_2, s3056[0]);
    wire[0:0] s6275, in6275_1, in6275_2;
    wire c6275;
    assign in6275_1 = {s3060[0]};
    assign in6275_2 = {s3061[0]};
    Full_Adder FA_6275(s6275, c6275, in6275_1, in6275_2, s3059[0]);
    wire[0:0] s6276, in6276_1, in6276_2;
    wire c6276;
    assign in6276_1 = {s3063[0]};
    assign in6276_2 = {s3064[0]};
    Full_Adder FA_6276(s6276, c6276, in6276_1, in6276_2, s3062[0]);
    wire[0:0] s6277, in6277_1, in6277_2;
    wire c6277;
    assign in6277_1 = {s3066[0]};
    assign in6277_2 = {s3067[0]};
    Full_Adder FA_6277(s6277, c6277, in6277_1, in6277_2, s3065[0]);
    wire[0:0] s6278, in6278_1, in6278_2;
    wire c6278;
    assign in6278_1 = {s3069[0]};
    assign in6278_2 = {s3070[0]};
    Full_Adder FA_6278(s6278, c6278, in6278_1, in6278_2, s3068[0]);
    wire[0:0] s6279, in6279_1, in6279_2;
    wire c6279;
    assign in6279_1 = {s3072[0]};
    assign in6279_2 = {s3073[0]};
    Full_Adder FA_6279(s6279, c6279, in6279_1, in6279_2, s3071[0]);
    wire[0:0] s6280, in6280_1, in6280_2;
    wire c6280;
    assign in6280_1 = {s3075[0]};
    assign in6280_2 = {s3076[0]};
    Full_Adder FA_6280(s6280, c6280, in6280_1, in6280_2, s3074[0]);
    wire[0:0] s6281, in6281_1, in6281_2;
    wire c6281;
    assign in6281_1 = {s3078[0]};
    assign in6281_2 = {s3079[0]};
    Full_Adder FA_6281(s6281, c6281, in6281_1, in6281_2, s3077[0]);
    wire[0:0] s6282, in6282_1, in6282_2;
    wire c6282;
    assign in6282_1 = {s528[0]};
    assign in6282_2 = {c3053};
    Full_Adder FA_6282(s6282, c6282, in6282_1, in6282_2, s527[0]);
    wire[0:0] s6283, in6283_1, in6283_2;
    wire c6283;
    assign in6283_1 = {c3055};
    assign in6283_2 = {c3056};
    Full_Adder FA_6283(s6283, c6283, in6283_1, in6283_2, c3054);
    wire[0:0] s6284, in6284_1, in6284_2;
    wire c6284;
    assign in6284_1 = {c3058};
    assign in6284_2 = {c3059};
    Full_Adder FA_6284(s6284, c6284, in6284_1, in6284_2, c3057);
    wire[0:0] s6285, in6285_1, in6285_2;
    wire c6285;
    assign in6285_1 = {c3061};
    assign in6285_2 = {c3062};
    Full_Adder FA_6285(s6285, c6285, in6285_1, in6285_2, c3060);
    wire[0:0] s6286, in6286_1, in6286_2;
    wire c6286;
    assign in6286_1 = {c3064};
    assign in6286_2 = {c3065};
    Full_Adder FA_6286(s6286, c6286, in6286_1, in6286_2, c3063);
    wire[0:0] s6287, in6287_1, in6287_2;
    wire c6287;
    assign in6287_1 = {c3067};
    assign in6287_2 = {c3068};
    Full_Adder FA_6287(s6287, c6287, in6287_1, in6287_2, c3066);
    wire[0:0] s6288, in6288_1, in6288_2;
    wire c6288;
    assign in6288_1 = {c3070};
    assign in6288_2 = {c3071};
    Full_Adder FA_6288(s6288, c6288, in6288_1, in6288_2, c3069);
    wire[0:0] s6289, in6289_1, in6289_2;
    wire c6289;
    assign in6289_1 = {c3073};
    assign in6289_2 = {c3074};
    Full_Adder FA_6289(s6289, c6289, in6289_1, in6289_2, c3072);
    wire[0:0] s6290, in6290_1, in6290_2;
    wire c6290;
    assign in6290_1 = {c3076};
    assign in6290_2 = {c3077};
    Full_Adder FA_6290(s6290, c6290, in6290_1, in6290_2, c3075);
    wire[0:0] s6291, in6291_1, in6291_2;
    wire c6291;
    assign in6291_1 = {c3079};
    assign in6291_2 = {c3080};
    Full_Adder FA_6291(s6291, c6291, in6291_1, in6291_2, c3078);
    wire[0:0] s6292, in6292_1, in6292_2;
    wire c6292;
    assign in6292_1 = {s3082[0]};
    assign in6292_2 = {s3083[0]};
    Full_Adder FA_6292(s6292, c6292, in6292_1, in6292_2, s3081[0]);
    wire[0:0] s6293, in6293_1, in6293_2;
    wire c6293;
    assign in6293_1 = {s3085[0]};
    assign in6293_2 = {s3086[0]};
    Full_Adder FA_6293(s6293, c6293, in6293_1, in6293_2, s3084[0]);
    wire[0:0] s6294, in6294_1, in6294_2;
    wire c6294;
    assign in6294_1 = {s3088[0]};
    assign in6294_2 = {s3089[0]};
    Full_Adder FA_6294(s6294, c6294, in6294_1, in6294_2, s3087[0]);
    wire[0:0] s6295, in6295_1, in6295_2;
    wire c6295;
    assign in6295_1 = {s3091[0]};
    assign in6295_2 = {s3092[0]};
    Full_Adder FA_6295(s6295, c6295, in6295_1, in6295_2, s3090[0]);
    wire[0:0] s6296, in6296_1, in6296_2;
    wire c6296;
    assign in6296_1 = {s3094[0]};
    assign in6296_2 = {s3095[0]};
    Full_Adder FA_6296(s6296, c6296, in6296_1, in6296_2, s3093[0]);
    wire[0:0] s6297, in6297_1, in6297_2;
    wire c6297;
    assign in6297_1 = {s3097[0]};
    assign in6297_2 = {s3098[0]};
    Full_Adder FA_6297(s6297, c6297, in6297_1, in6297_2, s3096[0]);
    wire[0:0] s6298, in6298_1, in6298_2;
    wire c6298;
    assign in6298_1 = {s3100[0]};
    assign in6298_2 = {s3101[0]};
    Full_Adder FA_6298(s6298, c6298, in6298_1, in6298_2, s3099[0]);
    wire[0:0] s6299, in6299_1, in6299_2;
    wire c6299;
    assign in6299_1 = {s3103[0]};
    assign in6299_2 = {s3104[0]};
    Full_Adder FA_6299(s6299, c6299, in6299_1, in6299_2, s3102[0]);
    wire[0:0] s6300, in6300_1, in6300_2;
    wire c6300;
    assign in6300_1 = {s3106[0]};
    assign in6300_2 = {s3107[0]};
    Full_Adder FA_6300(s6300, c6300, in6300_1, in6300_2, s3105[0]);
    wire[0:0] s6301, in6301_1, in6301_2;
    wire c6301;
    assign in6301_1 = {s561[0]};
    assign in6301_2 = {c3081};
    Full_Adder FA_6301(s6301, c6301, in6301_1, in6301_2, s560[0]);
    wire[0:0] s6302, in6302_1, in6302_2;
    wire c6302;
    assign in6302_1 = {c3083};
    assign in6302_2 = {c3084};
    Full_Adder FA_6302(s6302, c6302, in6302_1, in6302_2, c3082);
    wire[0:0] s6303, in6303_1, in6303_2;
    wire c6303;
    assign in6303_1 = {c3086};
    assign in6303_2 = {c3087};
    Full_Adder FA_6303(s6303, c6303, in6303_1, in6303_2, c3085);
    wire[0:0] s6304, in6304_1, in6304_2;
    wire c6304;
    assign in6304_1 = {c3089};
    assign in6304_2 = {c3090};
    Full_Adder FA_6304(s6304, c6304, in6304_1, in6304_2, c3088);
    wire[0:0] s6305, in6305_1, in6305_2;
    wire c6305;
    assign in6305_1 = {c3092};
    assign in6305_2 = {c3093};
    Full_Adder FA_6305(s6305, c6305, in6305_1, in6305_2, c3091);
    wire[0:0] s6306, in6306_1, in6306_2;
    wire c6306;
    assign in6306_1 = {c3095};
    assign in6306_2 = {c3096};
    Full_Adder FA_6306(s6306, c6306, in6306_1, in6306_2, c3094);
    wire[0:0] s6307, in6307_1, in6307_2;
    wire c6307;
    assign in6307_1 = {c3098};
    assign in6307_2 = {c3099};
    Full_Adder FA_6307(s6307, c6307, in6307_1, in6307_2, c3097);
    wire[0:0] s6308, in6308_1, in6308_2;
    wire c6308;
    assign in6308_1 = {c3101};
    assign in6308_2 = {c3102};
    Full_Adder FA_6308(s6308, c6308, in6308_1, in6308_2, c3100);
    wire[0:0] s6309, in6309_1, in6309_2;
    wire c6309;
    assign in6309_1 = {c3104};
    assign in6309_2 = {c3105};
    Full_Adder FA_6309(s6309, c6309, in6309_1, in6309_2, c3103);
    wire[0:0] s6310, in6310_1, in6310_2;
    wire c6310;
    assign in6310_1 = {c3107};
    assign in6310_2 = {c3108};
    Full_Adder FA_6310(s6310, c6310, in6310_1, in6310_2, c3106);
    wire[0:0] s6311, in6311_1, in6311_2;
    wire c6311;
    assign in6311_1 = {s3110[0]};
    assign in6311_2 = {s3111[0]};
    Full_Adder FA_6311(s6311, c6311, in6311_1, in6311_2, s3109[0]);
    wire[0:0] s6312, in6312_1, in6312_2;
    wire c6312;
    assign in6312_1 = {s3113[0]};
    assign in6312_2 = {s3114[0]};
    Full_Adder FA_6312(s6312, c6312, in6312_1, in6312_2, s3112[0]);
    wire[0:0] s6313, in6313_1, in6313_2;
    wire c6313;
    assign in6313_1 = {s3116[0]};
    assign in6313_2 = {s3117[0]};
    Full_Adder FA_6313(s6313, c6313, in6313_1, in6313_2, s3115[0]);
    wire[0:0] s6314, in6314_1, in6314_2;
    wire c6314;
    assign in6314_1 = {s3119[0]};
    assign in6314_2 = {s3120[0]};
    Full_Adder FA_6314(s6314, c6314, in6314_1, in6314_2, s3118[0]);
    wire[0:0] s6315, in6315_1, in6315_2;
    wire c6315;
    assign in6315_1 = {s3122[0]};
    assign in6315_2 = {s3123[0]};
    Full_Adder FA_6315(s6315, c6315, in6315_1, in6315_2, s3121[0]);
    wire[0:0] s6316, in6316_1, in6316_2;
    wire c6316;
    assign in6316_1 = {s3125[0]};
    assign in6316_2 = {s3126[0]};
    Full_Adder FA_6316(s6316, c6316, in6316_1, in6316_2, s3124[0]);
    wire[0:0] s6317, in6317_1, in6317_2;
    wire c6317;
    assign in6317_1 = {s3128[0]};
    assign in6317_2 = {s3129[0]};
    Full_Adder FA_6317(s6317, c6317, in6317_1, in6317_2, s3127[0]);
    wire[0:0] s6318, in6318_1, in6318_2;
    wire c6318;
    assign in6318_1 = {s3131[0]};
    assign in6318_2 = {s3132[0]};
    Full_Adder FA_6318(s6318, c6318, in6318_1, in6318_2, s3130[0]);
    wire[0:0] s6319, in6319_1, in6319_2;
    wire c6319;
    assign in6319_1 = {s3134[0]};
    assign in6319_2 = {s3135[0]};
    Full_Adder FA_6319(s6319, c6319, in6319_1, in6319_2, s3133[0]);
    wire[0:0] s6320, in6320_1, in6320_2;
    wire c6320;
    assign in6320_1 = {s595[0]};
    assign in6320_2 = {c3109};
    Full_Adder FA_6320(s6320, c6320, in6320_1, in6320_2, s594[0]);
    wire[0:0] s6321, in6321_1, in6321_2;
    wire c6321;
    assign in6321_1 = {c3111};
    assign in6321_2 = {c3112};
    Full_Adder FA_6321(s6321, c6321, in6321_1, in6321_2, c3110);
    wire[0:0] s6322, in6322_1, in6322_2;
    wire c6322;
    assign in6322_1 = {c3114};
    assign in6322_2 = {c3115};
    Full_Adder FA_6322(s6322, c6322, in6322_1, in6322_2, c3113);
    wire[0:0] s6323, in6323_1, in6323_2;
    wire c6323;
    assign in6323_1 = {c3117};
    assign in6323_2 = {c3118};
    Full_Adder FA_6323(s6323, c6323, in6323_1, in6323_2, c3116);
    wire[0:0] s6324, in6324_1, in6324_2;
    wire c6324;
    assign in6324_1 = {c3120};
    assign in6324_2 = {c3121};
    Full_Adder FA_6324(s6324, c6324, in6324_1, in6324_2, c3119);
    wire[0:0] s6325, in6325_1, in6325_2;
    wire c6325;
    assign in6325_1 = {c3123};
    assign in6325_2 = {c3124};
    Full_Adder FA_6325(s6325, c6325, in6325_1, in6325_2, c3122);
    wire[0:0] s6326, in6326_1, in6326_2;
    wire c6326;
    assign in6326_1 = {c3126};
    assign in6326_2 = {c3127};
    Full_Adder FA_6326(s6326, c6326, in6326_1, in6326_2, c3125);
    wire[0:0] s6327, in6327_1, in6327_2;
    wire c6327;
    assign in6327_1 = {c3129};
    assign in6327_2 = {c3130};
    Full_Adder FA_6327(s6327, c6327, in6327_1, in6327_2, c3128);
    wire[0:0] s6328, in6328_1, in6328_2;
    wire c6328;
    assign in6328_1 = {c3132};
    assign in6328_2 = {c3133};
    Full_Adder FA_6328(s6328, c6328, in6328_1, in6328_2, c3131);
    wire[0:0] s6329, in6329_1, in6329_2;
    wire c6329;
    assign in6329_1 = {c3135};
    assign in6329_2 = {c3136};
    Full_Adder FA_6329(s6329, c6329, in6329_1, in6329_2, c3134);
    wire[0:0] s6330, in6330_1, in6330_2;
    wire c6330;
    assign in6330_1 = {s3138[0]};
    assign in6330_2 = {s3139[0]};
    Full_Adder FA_6330(s6330, c6330, in6330_1, in6330_2, s3137[0]);
    wire[0:0] s6331, in6331_1, in6331_2;
    wire c6331;
    assign in6331_1 = {s3141[0]};
    assign in6331_2 = {s3142[0]};
    Full_Adder FA_6331(s6331, c6331, in6331_1, in6331_2, s3140[0]);
    wire[0:0] s6332, in6332_1, in6332_2;
    wire c6332;
    assign in6332_1 = {s3144[0]};
    assign in6332_2 = {s3145[0]};
    Full_Adder FA_6332(s6332, c6332, in6332_1, in6332_2, s3143[0]);
    wire[0:0] s6333, in6333_1, in6333_2;
    wire c6333;
    assign in6333_1 = {s3147[0]};
    assign in6333_2 = {s3148[0]};
    Full_Adder FA_6333(s6333, c6333, in6333_1, in6333_2, s3146[0]);
    wire[0:0] s6334, in6334_1, in6334_2;
    wire c6334;
    assign in6334_1 = {s3150[0]};
    assign in6334_2 = {s3151[0]};
    Full_Adder FA_6334(s6334, c6334, in6334_1, in6334_2, s3149[0]);
    wire[0:0] s6335, in6335_1, in6335_2;
    wire c6335;
    assign in6335_1 = {s3153[0]};
    assign in6335_2 = {s3154[0]};
    Full_Adder FA_6335(s6335, c6335, in6335_1, in6335_2, s3152[0]);
    wire[0:0] s6336, in6336_1, in6336_2;
    wire c6336;
    assign in6336_1 = {s3156[0]};
    assign in6336_2 = {s3157[0]};
    Full_Adder FA_6336(s6336, c6336, in6336_1, in6336_2, s3155[0]);
    wire[0:0] s6337, in6337_1, in6337_2;
    wire c6337;
    assign in6337_1 = {s3159[0]};
    assign in6337_2 = {s3160[0]};
    Full_Adder FA_6337(s6337, c6337, in6337_1, in6337_2, s3158[0]);
    wire[0:0] s6338, in6338_1, in6338_2;
    wire c6338;
    assign in6338_1 = {s3162[0]};
    assign in6338_2 = {s3163[0]};
    Full_Adder FA_6338(s6338, c6338, in6338_1, in6338_2, s3161[0]);
    wire[0:0] s6339, in6339_1, in6339_2;
    wire c6339;
    assign in6339_1 = {s630[0]};
    assign in6339_2 = {c3137};
    Full_Adder FA_6339(s6339, c6339, in6339_1, in6339_2, s629[0]);
    wire[0:0] s6340, in6340_1, in6340_2;
    wire c6340;
    assign in6340_1 = {c3139};
    assign in6340_2 = {c3140};
    Full_Adder FA_6340(s6340, c6340, in6340_1, in6340_2, c3138);
    wire[0:0] s6341, in6341_1, in6341_2;
    wire c6341;
    assign in6341_1 = {c3142};
    assign in6341_2 = {c3143};
    Full_Adder FA_6341(s6341, c6341, in6341_1, in6341_2, c3141);
    wire[0:0] s6342, in6342_1, in6342_2;
    wire c6342;
    assign in6342_1 = {c3145};
    assign in6342_2 = {c3146};
    Full_Adder FA_6342(s6342, c6342, in6342_1, in6342_2, c3144);
    wire[0:0] s6343, in6343_1, in6343_2;
    wire c6343;
    assign in6343_1 = {c3148};
    assign in6343_2 = {c3149};
    Full_Adder FA_6343(s6343, c6343, in6343_1, in6343_2, c3147);
    wire[0:0] s6344, in6344_1, in6344_2;
    wire c6344;
    assign in6344_1 = {c3151};
    assign in6344_2 = {c3152};
    Full_Adder FA_6344(s6344, c6344, in6344_1, in6344_2, c3150);
    wire[0:0] s6345, in6345_1, in6345_2;
    wire c6345;
    assign in6345_1 = {c3154};
    assign in6345_2 = {c3155};
    Full_Adder FA_6345(s6345, c6345, in6345_1, in6345_2, c3153);
    wire[0:0] s6346, in6346_1, in6346_2;
    wire c6346;
    assign in6346_1 = {c3157};
    assign in6346_2 = {c3158};
    Full_Adder FA_6346(s6346, c6346, in6346_1, in6346_2, c3156);
    wire[0:0] s6347, in6347_1, in6347_2;
    wire c6347;
    assign in6347_1 = {c3160};
    assign in6347_2 = {c3161};
    Full_Adder FA_6347(s6347, c6347, in6347_1, in6347_2, c3159);
    wire[0:0] s6348, in6348_1, in6348_2;
    wire c6348;
    assign in6348_1 = {c3163};
    assign in6348_2 = {c3164};
    Full_Adder FA_6348(s6348, c6348, in6348_1, in6348_2, c3162);
    wire[0:0] s6349, in6349_1, in6349_2;
    wire c6349;
    assign in6349_1 = {s3166[0]};
    assign in6349_2 = {s3167[0]};
    Full_Adder FA_6349(s6349, c6349, in6349_1, in6349_2, s3165[0]);
    wire[0:0] s6350, in6350_1, in6350_2;
    wire c6350;
    assign in6350_1 = {s3169[0]};
    assign in6350_2 = {s3170[0]};
    Full_Adder FA_6350(s6350, c6350, in6350_1, in6350_2, s3168[0]);
    wire[0:0] s6351, in6351_1, in6351_2;
    wire c6351;
    assign in6351_1 = {s3172[0]};
    assign in6351_2 = {s3173[0]};
    Full_Adder FA_6351(s6351, c6351, in6351_1, in6351_2, s3171[0]);
    wire[0:0] s6352, in6352_1, in6352_2;
    wire c6352;
    assign in6352_1 = {s3175[0]};
    assign in6352_2 = {s3176[0]};
    Full_Adder FA_6352(s6352, c6352, in6352_1, in6352_2, s3174[0]);
    wire[0:0] s6353, in6353_1, in6353_2;
    wire c6353;
    assign in6353_1 = {s3178[0]};
    assign in6353_2 = {s3179[0]};
    Full_Adder FA_6353(s6353, c6353, in6353_1, in6353_2, s3177[0]);
    wire[0:0] s6354, in6354_1, in6354_2;
    wire c6354;
    assign in6354_1 = {s3181[0]};
    assign in6354_2 = {s3182[0]};
    Full_Adder FA_6354(s6354, c6354, in6354_1, in6354_2, s3180[0]);
    wire[0:0] s6355, in6355_1, in6355_2;
    wire c6355;
    assign in6355_1 = {s3184[0]};
    assign in6355_2 = {s3185[0]};
    Full_Adder FA_6355(s6355, c6355, in6355_1, in6355_2, s3183[0]);
    wire[0:0] s6356, in6356_1, in6356_2;
    wire c6356;
    assign in6356_1 = {s3187[0]};
    assign in6356_2 = {s3188[0]};
    Full_Adder FA_6356(s6356, c6356, in6356_1, in6356_2, s3186[0]);
    wire[0:0] s6357, in6357_1, in6357_2;
    wire c6357;
    assign in6357_1 = {s3190[0]};
    assign in6357_2 = {s3191[0]};
    Full_Adder FA_6357(s6357, c6357, in6357_1, in6357_2, s3189[0]);
    wire[0:0] s6358, in6358_1, in6358_2;
    wire c6358;
    assign in6358_1 = {s666[0]};
    assign in6358_2 = {c3165};
    Full_Adder FA_6358(s6358, c6358, in6358_1, in6358_2, s665[0]);
    wire[0:0] s6359, in6359_1, in6359_2;
    wire c6359;
    assign in6359_1 = {c3167};
    assign in6359_2 = {c3168};
    Full_Adder FA_6359(s6359, c6359, in6359_1, in6359_2, c3166);
    wire[0:0] s6360, in6360_1, in6360_2;
    wire c6360;
    assign in6360_1 = {c3170};
    assign in6360_2 = {c3171};
    Full_Adder FA_6360(s6360, c6360, in6360_1, in6360_2, c3169);
    wire[0:0] s6361, in6361_1, in6361_2;
    wire c6361;
    assign in6361_1 = {c3173};
    assign in6361_2 = {c3174};
    Full_Adder FA_6361(s6361, c6361, in6361_1, in6361_2, c3172);
    wire[0:0] s6362, in6362_1, in6362_2;
    wire c6362;
    assign in6362_1 = {c3176};
    assign in6362_2 = {c3177};
    Full_Adder FA_6362(s6362, c6362, in6362_1, in6362_2, c3175);
    wire[0:0] s6363, in6363_1, in6363_2;
    wire c6363;
    assign in6363_1 = {c3179};
    assign in6363_2 = {c3180};
    Full_Adder FA_6363(s6363, c6363, in6363_1, in6363_2, c3178);
    wire[0:0] s6364, in6364_1, in6364_2;
    wire c6364;
    assign in6364_1 = {c3182};
    assign in6364_2 = {c3183};
    Full_Adder FA_6364(s6364, c6364, in6364_1, in6364_2, c3181);
    wire[0:0] s6365, in6365_1, in6365_2;
    wire c6365;
    assign in6365_1 = {c3185};
    assign in6365_2 = {c3186};
    Full_Adder FA_6365(s6365, c6365, in6365_1, in6365_2, c3184);
    wire[0:0] s6366, in6366_1, in6366_2;
    wire c6366;
    assign in6366_1 = {c3188};
    assign in6366_2 = {c3189};
    Full_Adder FA_6366(s6366, c6366, in6366_1, in6366_2, c3187);
    wire[0:0] s6367, in6367_1, in6367_2;
    wire c6367;
    assign in6367_1 = {c3191};
    assign in6367_2 = {c3192};
    Full_Adder FA_6367(s6367, c6367, in6367_1, in6367_2, c3190);
    wire[0:0] s6368, in6368_1, in6368_2;
    wire c6368;
    assign in6368_1 = {s3194[0]};
    assign in6368_2 = {s3195[0]};
    Full_Adder FA_6368(s6368, c6368, in6368_1, in6368_2, s3193[0]);
    wire[0:0] s6369, in6369_1, in6369_2;
    wire c6369;
    assign in6369_1 = {s3197[0]};
    assign in6369_2 = {s3198[0]};
    Full_Adder FA_6369(s6369, c6369, in6369_1, in6369_2, s3196[0]);
    wire[0:0] s6370, in6370_1, in6370_2;
    wire c6370;
    assign in6370_1 = {s3200[0]};
    assign in6370_2 = {s3201[0]};
    Full_Adder FA_6370(s6370, c6370, in6370_1, in6370_2, s3199[0]);
    wire[0:0] s6371, in6371_1, in6371_2;
    wire c6371;
    assign in6371_1 = {s3203[0]};
    assign in6371_2 = {s3204[0]};
    Full_Adder FA_6371(s6371, c6371, in6371_1, in6371_2, s3202[0]);
    wire[0:0] s6372, in6372_1, in6372_2;
    wire c6372;
    assign in6372_1 = {s3206[0]};
    assign in6372_2 = {s3207[0]};
    Full_Adder FA_6372(s6372, c6372, in6372_1, in6372_2, s3205[0]);
    wire[0:0] s6373, in6373_1, in6373_2;
    wire c6373;
    assign in6373_1 = {s3209[0]};
    assign in6373_2 = {s3210[0]};
    Full_Adder FA_6373(s6373, c6373, in6373_1, in6373_2, s3208[0]);
    wire[0:0] s6374, in6374_1, in6374_2;
    wire c6374;
    assign in6374_1 = {s3212[0]};
    assign in6374_2 = {s3213[0]};
    Full_Adder FA_6374(s6374, c6374, in6374_1, in6374_2, s3211[0]);
    wire[0:0] s6375, in6375_1, in6375_2;
    wire c6375;
    assign in6375_1 = {s3215[0]};
    assign in6375_2 = {s3216[0]};
    Full_Adder FA_6375(s6375, c6375, in6375_1, in6375_2, s3214[0]);
    wire[0:0] s6376, in6376_1, in6376_2;
    wire c6376;
    assign in6376_1 = {s3218[0]};
    assign in6376_2 = {s3219[0]};
    Full_Adder FA_6376(s6376, c6376, in6376_1, in6376_2, s3217[0]);
    wire[0:0] s6377, in6377_1, in6377_2;
    wire c6377;
    assign in6377_1 = {s703[0]};
    assign in6377_2 = {c3193};
    Full_Adder FA_6377(s6377, c6377, in6377_1, in6377_2, s702[0]);
    wire[0:0] s6378, in6378_1, in6378_2;
    wire c6378;
    assign in6378_1 = {c3195};
    assign in6378_2 = {c3196};
    Full_Adder FA_6378(s6378, c6378, in6378_1, in6378_2, c3194);
    wire[0:0] s6379, in6379_1, in6379_2;
    wire c6379;
    assign in6379_1 = {c3198};
    assign in6379_2 = {c3199};
    Full_Adder FA_6379(s6379, c6379, in6379_1, in6379_2, c3197);
    wire[0:0] s6380, in6380_1, in6380_2;
    wire c6380;
    assign in6380_1 = {c3201};
    assign in6380_2 = {c3202};
    Full_Adder FA_6380(s6380, c6380, in6380_1, in6380_2, c3200);
    wire[0:0] s6381, in6381_1, in6381_2;
    wire c6381;
    assign in6381_1 = {c3204};
    assign in6381_2 = {c3205};
    Full_Adder FA_6381(s6381, c6381, in6381_1, in6381_2, c3203);
    wire[0:0] s6382, in6382_1, in6382_2;
    wire c6382;
    assign in6382_1 = {c3207};
    assign in6382_2 = {c3208};
    Full_Adder FA_6382(s6382, c6382, in6382_1, in6382_2, c3206);
    wire[0:0] s6383, in6383_1, in6383_2;
    wire c6383;
    assign in6383_1 = {c3210};
    assign in6383_2 = {c3211};
    Full_Adder FA_6383(s6383, c6383, in6383_1, in6383_2, c3209);
    wire[0:0] s6384, in6384_1, in6384_2;
    wire c6384;
    assign in6384_1 = {c3213};
    assign in6384_2 = {c3214};
    Full_Adder FA_6384(s6384, c6384, in6384_1, in6384_2, c3212);
    wire[0:0] s6385, in6385_1, in6385_2;
    wire c6385;
    assign in6385_1 = {c3216};
    assign in6385_2 = {c3217};
    Full_Adder FA_6385(s6385, c6385, in6385_1, in6385_2, c3215);
    wire[0:0] s6386, in6386_1, in6386_2;
    wire c6386;
    assign in6386_1 = {c3219};
    assign in6386_2 = {c3220};
    Full_Adder FA_6386(s6386, c6386, in6386_1, in6386_2, c3218);
    wire[0:0] s6387, in6387_1, in6387_2;
    wire c6387;
    assign in6387_1 = {s3222[0]};
    assign in6387_2 = {s3223[0]};
    Full_Adder FA_6387(s6387, c6387, in6387_1, in6387_2, s3221[0]);
    wire[0:0] s6388, in6388_1, in6388_2;
    wire c6388;
    assign in6388_1 = {s3225[0]};
    assign in6388_2 = {s3226[0]};
    Full_Adder FA_6388(s6388, c6388, in6388_1, in6388_2, s3224[0]);
    wire[0:0] s6389, in6389_1, in6389_2;
    wire c6389;
    assign in6389_1 = {s3228[0]};
    assign in6389_2 = {s3229[0]};
    Full_Adder FA_6389(s6389, c6389, in6389_1, in6389_2, s3227[0]);
    wire[0:0] s6390, in6390_1, in6390_2;
    wire c6390;
    assign in6390_1 = {s3231[0]};
    assign in6390_2 = {s3232[0]};
    Full_Adder FA_6390(s6390, c6390, in6390_1, in6390_2, s3230[0]);
    wire[0:0] s6391, in6391_1, in6391_2;
    wire c6391;
    assign in6391_1 = {s3234[0]};
    assign in6391_2 = {s3235[0]};
    Full_Adder FA_6391(s6391, c6391, in6391_1, in6391_2, s3233[0]);
    wire[0:0] s6392, in6392_1, in6392_2;
    wire c6392;
    assign in6392_1 = {s3237[0]};
    assign in6392_2 = {s3238[0]};
    Full_Adder FA_6392(s6392, c6392, in6392_1, in6392_2, s3236[0]);
    wire[0:0] s6393, in6393_1, in6393_2;
    wire c6393;
    assign in6393_1 = {s3240[0]};
    assign in6393_2 = {s3241[0]};
    Full_Adder FA_6393(s6393, c6393, in6393_1, in6393_2, s3239[0]);
    wire[0:0] s6394, in6394_1, in6394_2;
    wire c6394;
    assign in6394_1 = {s3243[0]};
    assign in6394_2 = {s3244[0]};
    Full_Adder FA_6394(s6394, c6394, in6394_1, in6394_2, s3242[0]);
    wire[0:0] s6395, in6395_1, in6395_2;
    wire c6395;
    assign in6395_1 = {s3246[0]};
    assign in6395_2 = {s3247[0]};
    Full_Adder FA_6395(s6395, c6395, in6395_1, in6395_2, s3245[0]);
    wire[0:0] s6396, in6396_1, in6396_2;
    wire c6396;
    assign in6396_1 = {s741[0]};
    assign in6396_2 = {c3221};
    Full_Adder FA_6396(s6396, c6396, in6396_1, in6396_2, s740[0]);
    wire[0:0] s6397, in6397_1, in6397_2;
    wire c6397;
    assign in6397_1 = {c3223};
    assign in6397_2 = {c3224};
    Full_Adder FA_6397(s6397, c6397, in6397_1, in6397_2, c3222);
    wire[0:0] s6398, in6398_1, in6398_2;
    wire c6398;
    assign in6398_1 = {c3226};
    assign in6398_2 = {c3227};
    Full_Adder FA_6398(s6398, c6398, in6398_1, in6398_2, c3225);
    wire[0:0] s6399, in6399_1, in6399_2;
    wire c6399;
    assign in6399_1 = {c3229};
    assign in6399_2 = {c3230};
    Full_Adder FA_6399(s6399, c6399, in6399_1, in6399_2, c3228);
    wire[0:0] s6400, in6400_1, in6400_2;
    wire c6400;
    assign in6400_1 = {c3232};
    assign in6400_2 = {c3233};
    Full_Adder FA_6400(s6400, c6400, in6400_1, in6400_2, c3231);
    wire[0:0] s6401, in6401_1, in6401_2;
    wire c6401;
    assign in6401_1 = {c3235};
    assign in6401_2 = {c3236};
    Full_Adder FA_6401(s6401, c6401, in6401_1, in6401_2, c3234);
    wire[0:0] s6402, in6402_1, in6402_2;
    wire c6402;
    assign in6402_1 = {c3238};
    assign in6402_2 = {c3239};
    Full_Adder FA_6402(s6402, c6402, in6402_1, in6402_2, c3237);
    wire[0:0] s6403, in6403_1, in6403_2;
    wire c6403;
    assign in6403_1 = {c3241};
    assign in6403_2 = {c3242};
    Full_Adder FA_6403(s6403, c6403, in6403_1, in6403_2, c3240);
    wire[0:0] s6404, in6404_1, in6404_2;
    wire c6404;
    assign in6404_1 = {c3244};
    assign in6404_2 = {c3245};
    Full_Adder FA_6404(s6404, c6404, in6404_1, in6404_2, c3243);
    wire[0:0] s6405, in6405_1, in6405_2;
    wire c6405;
    assign in6405_1 = {c3247};
    assign in6405_2 = {c3248};
    Full_Adder FA_6405(s6405, c6405, in6405_1, in6405_2, c3246);
    wire[0:0] s6406, in6406_1, in6406_2;
    wire c6406;
    assign in6406_1 = {s3250[0]};
    assign in6406_2 = {s3251[0]};
    Full_Adder FA_6406(s6406, c6406, in6406_1, in6406_2, s3249[0]);
    wire[0:0] s6407, in6407_1, in6407_2;
    wire c6407;
    assign in6407_1 = {s3253[0]};
    assign in6407_2 = {s3254[0]};
    Full_Adder FA_6407(s6407, c6407, in6407_1, in6407_2, s3252[0]);
    wire[0:0] s6408, in6408_1, in6408_2;
    wire c6408;
    assign in6408_1 = {s3256[0]};
    assign in6408_2 = {s3257[0]};
    Full_Adder FA_6408(s6408, c6408, in6408_1, in6408_2, s3255[0]);
    wire[0:0] s6409, in6409_1, in6409_2;
    wire c6409;
    assign in6409_1 = {s3259[0]};
    assign in6409_2 = {s3260[0]};
    Full_Adder FA_6409(s6409, c6409, in6409_1, in6409_2, s3258[0]);
    wire[0:0] s6410, in6410_1, in6410_2;
    wire c6410;
    assign in6410_1 = {s3262[0]};
    assign in6410_2 = {s3263[0]};
    Full_Adder FA_6410(s6410, c6410, in6410_1, in6410_2, s3261[0]);
    wire[0:0] s6411, in6411_1, in6411_2;
    wire c6411;
    assign in6411_1 = {s3265[0]};
    assign in6411_2 = {s3266[0]};
    Full_Adder FA_6411(s6411, c6411, in6411_1, in6411_2, s3264[0]);
    wire[0:0] s6412, in6412_1, in6412_2;
    wire c6412;
    assign in6412_1 = {s3268[0]};
    assign in6412_2 = {s3269[0]};
    Full_Adder FA_6412(s6412, c6412, in6412_1, in6412_2, s3267[0]);
    wire[0:0] s6413, in6413_1, in6413_2;
    wire c6413;
    assign in6413_1 = {s3271[0]};
    assign in6413_2 = {s3272[0]};
    Full_Adder FA_6413(s6413, c6413, in6413_1, in6413_2, s3270[0]);
    wire[0:0] s6414, in6414_1, in6414_2;
    wire c6414;
    assign in6414_1 = {s3274[0]};
    assign in6414_2 = {s3275[0]};
    Full_Adder FA_6414(s6414, c6414, in6414_1, in6414_2, s3273[0]);
    wire[0:0] s6415, in6415_1, in6415_2;
    wire c6415;
    assign in6415_1 = {s780[0]};
    assign in6415_2 = {c3249};
    Full_Adder FA_6415(s6415, c6415, in6415_1, in6415_2, s779[0]);
    wire[0:0] s6416, in6416_1, in6416_2;
    wire c6416;
    assign in6416_1 = {c3251};
    assign in6416_2 = {c3252};
    Full_Adder FA_6416(s6416, c6416, in6416_1, in6416_2, c3250);
    wire[0:0] s6417, in6417_1, in6417_2;
    wire c6417;
    assign in6417_1 = {c3254};
    assign in6417_2 = {c3255};
    Full_Adder FA_6417(s6417, c6417, in6417_1, in6417_2, c3253);
    wire[0:0] s6418, in6418_1, in6418_2;
    wire c6418;
    assign in6418_1 = {c3257};
    assign in6418_2 = {c3258};
    Full_Adder FA_6418(s6418, c6418, in6418_1, in6418_2, c3256);
    wire[0:0] s6419, in6419_1, in6419_2;
    wire c6419;
    assign in6419_1 = {c3260};
    assign in6419_2 = {c3261};
    Full_Adder FA_6419(s6419, c6419, in6419_1, in6419_2, c3259);
    wire[0:0] s6420, in6420_1, in6420_2;
    wire c6420;
    assign in6420_1 = {c3263};
    assign in6420_2 = {c3264};
    Full_Adder FA_6420(s6420, c6420, in6420_1, in6420_2, c3262);
    wire[0:0] s6421, in6421_1, in6421_2;
    wire c6421;
    assign in6421_1 = {c3266};
    assign in6421_2 = {c3267};
    Full_Adder FA_6421(s6421, c6421, in6421_1, in6421_2, c3265);
    wire[0:0] s6422, in6422_1, in6422_2;
    wire c6422;
    assign in6422_1 = {c3269};
    assign in6422_2 = {c3270};
    Full_Adder FA_6422(s6422, c6422, in6422_1, in6422_2, c3268);
    wire[0:0] s6423, in6423_1, in6423_2;
    wire c6423;
    assign in6423_1 = {c3272};
    assign in6423_2 = {c3273};
    Full_Adder FA_6423(s6423, c6423, in6423_1, in6423_2, c3271);
    wire[0:0] s6424, in6424_1, in6424_2;
    wire c6424;
    assign in6424_1 = {c3275};
    assign in6424_2 = {c3276};
    Full_Adder FA_6424(s6424, c6424, in6424_1, in6424_2, c3274);
    wire[0:0] s6425, in6425_1, in6425_2;
    wire c6425;
    assign in6425_1 = {s3278[0]};
    assign in6425_2 = {s3279[0]};
    Full_Adder FA_6425(s6425, c6425, in6425_1, in6425_2, s3277[0]);
    wire[0:0] s6426, in6426_1, in6426_2;
    wire c6426;
    assign in6426_1 = {s3281[0]};
    assign in6426_2 = {s3282[0]};
    Full_Adder FA_6426(s6426, c6426, in6426_1, in6426_2, s3280[0]);
    wire[0:0] s6427, in6427_1, in6427_2;
    wire c6427;
    assign in6427_1 = {s3284[0]};
    assign in6427_2 = {s3285[0]};
    Full_Adder FA_6427(s6427, c6427, in6427_1, in6427_2, s3283[0]);
    wire[0:0] s6428, in6428_1, in6428_2;
    wire c6428;
    assign in6428_1 = {s3287[0]};
    assign in6428_2 = {s3288[0]};
    Full_Adder FA_6428(s6428, c6428, in6428_1, in6428_2, s3286[0]);
    wire[0:0] s6429, in6429_1, in6429_2;
    wire c6429;
    assign in6429_1 = {s3290[0]};
    assign in6429_2 = {s3291[0]};
    Full_Adder FA_6429(s6429, c6429, in6429_1, in6429_2, s3289[0]);
    wire[0:0] s6430, in6430_1, in6430_2;
    wire c6430;
    assign in6430_1 = {s3293[0]};
    assign in6430_2 = {s3294[0]};
    Full_Adder FA_6430(s6430, c6430, in6430_1, in6430_2, s3292[0]);
    wire[0:0] s6431, in6431_1, in6431_2;
    wire c6431;
    assign in6431_1 = {s3296[0]};
    assign in6431_2 = {s3297[0]};
    Full_Adder FA_6431(s6431, c6431, in6431_1, in6431_2, s3295[0]);
    wire[0:0] s6432, in6432_1, in6432_2;
    wire c6432;
    assign in6432_1 = {s3299[0]};
    assign in6432_2 = {s3300[0]};
    Full_Adder FA_6432(s6432, c6432, in6432_1, in6432_2, s3298[0]);
    wire[0:0] s6433, in6433_1, in6433_2;
    wire c6433;
    assign in6433_1 = {s3302[0]};
    assign in6433_2 = {s3303[0]};
    Full_Adder FA_6433(s6433, c6433, in6433_1, in6433_2, s3301[0]);
    wire[0:0] s6434, in6434_1, in6434_2;
    wire c6434;
    assign in6434_1 = {s820[0]};
    assign in6434_2 = {c3277};
    Full_Adder FA_6434(s6434, c6434, in6434_1, in6434_2, s819[0]);
    wire[0:0] s6435, in6435_1, in6435_2;
    wire c6435;
    assign in6435_1 = {c3279};
    assign in6435_2 = {c3280};
    Full_Adder FA_6435(s6435, c6435, in6435_1, in6435_2, c3278);
    wire[0:0] s6436, in6436_1, in6436_2;
    wire c6436;
    assign in6436_1 = {c3282};
    assign in6436_2 = {c3283};
    Full_Adder FA_6436(s6436, c6436, in6436_1, in6436_2, c3281);
    wire[0:0] s6437, in6437_1, in6437_2;
    wire c6437;
    assign in6437_1 = {c3285};
    assign in6437_2 = {c3286};
    Full_Adder FA_6437(s6437, c6437, in6437_1, in6437_2, c3284);
    wire[0:0] s6438, in6438_1, in6438_2;
    wire c6438;
    assign in6438_1 = {c3288};
    assign in6438_2 = {c3289};
    Full_Adder FA_6438(s6438, c6438, in6438_1, in6438_2, c3287);
    wire[0:0] s6439, in6439_1, in6439_2;
    wire c6439;
    assign in6439_1 = {c3291};
    assign in6439_2 = {c3292};
    Full_Adder FA_6439(s6439, c6439, in6439_1, in6439_2, c3290);
    wire[0:0] s6440, in6440_1, in6440_2;
    wire c6440;
    assign in6440_1 = {c3294};
    assign in6440_2 = {c3295};
    Full_Adder FA_6440(s6440, c6440, in6440_1, in6440_2, c3293);
    wire[0:0] s6441, in6441_1, in6441_2;
    wire c6441;
    assign in6441_1 = {c3297};
    assign in6441_2 = {c3298};
    Full_Adder FA_6441(s6441, c6441, in6441_1, in6441_2, c3296);
    wire[0:0] s6442, in6442_1, in6442_2;
    wire c6442;
    assign in6442_1 = {c3300};
    assign in6442_2 = {c3301};
    Full_Adder FA_6442(s6442, c6442, in6442_1, in6442_2, c3299);
    wire[0:0] s6443, in6443_1, in6443_2;
    wire c6443;
    assign in6443_1 = {c3303};
    assign in6443_2 = {c3304};
    Full_Adder FA_6443(s6443, c6443, in6443_1, in6443_2, c3302);
    wire[0:0] s6444, in6444_1, in6444_2;
    wire c6444;
    assign in6444_1 = {s3306[0]};
    assign in6444_2 = {s3307[0]};
    Full_Adder FA_6444(s6444, c6444, in6444_1, in6444_2, s3305[0]);
    wire[0:0] s6445, in6445_1, in6445_2;
    wire c6445;
    assign in6445_1 = {s3309[0]};
    assign in6445_2 = {s3310[0]};
    Full_Adder FA_6445(s6445, c6445, in6445_1, in6445_2, s3308[0]);
    wire[0:0] s6446, in6446_1, in6446_2;
    wire c6446;
    assign in6446_1 = {s3312[0]};
    assign in6446_2 = {s3313[0]};
    Full_Adder FA_6446(s6446, c6446, in6446_1, in6446_2, s3311[0]);
    wire[0:0] s6447, in6447_1, in6447_2;
    wire c6447;
    assign in6447_1 = {s3315[0]};
    assign in6447_2 = {s3316[0]};
    Full_Adder FA_6447(s6447, c6447, in6447_1, in6447_2, s3314[0]);
    wire[0:0] s6448, in6448_1, in6448_2;
    wire c6448;
    assign in6448_1 = {s3318[0]};
    assign in6448_2 = {s3319[0]};
    Full_Adder FA_6448(s6448, c6448, in6448_1, in6448_2, s3317[0]);
    wire[0:0] s6449, in6449_1, in6449_2;
    wire c6449;
    assign in6449_1 = {s3321[0]};
    assign in6449_2 = {s3322[0]};
    Full_Adder FA_6449(s6449, c6449, in6449_1, in6449_2, s3320[0]);
    wire[0:0] s6450, in6450_1, in6450_2;
    wire c6450;
    assign in6450_1 = {s3324[0]};
    assign in6450_2 = {s3325[0]};
    Full_Adder FA_6450(s6450, c6450, in6450_1, in6450_2, s3323[0]);
    wire[0:0] s6451, in6451_1, in6451_2;
    wire c6451;
    assign in6451_1 = {s3327[0]};
    assign in6451_2 = {s3328[0]};
    Full_Adder FA_6451(s6451, c6451, in6451_1, in6451_2, s3326[0]);
    wire[0:0] s6452, in6452_1, in6452_2;
    wire c6452;
    assign in6452_1 = {s3330[0]};
    assign in6452_2 = {s3331[0]};
    Full_Adder FA_6452(s6452, c6452, in6452_1, in6452_2, s3329[0]);
    wire[0:0] s6453, in6453_1, in6453_2;
    wire c6453;
    assign in6453_1 = {s861[0]};
    assign in6453_2 = {c3305};
    Full_Adder FA_6453(s6453, c6453, in6453_1, in6453_2, s860[0]);
    wire[0:0] s6454, in6454_1, in6454_2;
    wire c6454;
    assign in6454_1 = {c3307};
    assign in6454_2 = {c3308};
    Full_Adder FA_6454(s6454, c6454, in6454_1, in6454_2, c3306);
    wire[0:0] s6455, in6455_1, in6455_2;
    wire c6455;
    assign in6455_1 = {c3310};
    assign in6455_2 = {c3311};
    Full_Adder FA_6455(s6455, c6455, in6455_1, in6455_2, c3309);
    wire[0:0] s6456, in6456_1, in6456_2;
    wire c6456;
    assign in6456_1 = {c3313};
    assign in6456_2 = {c3314};
    Full_Adder FA_6456(s6456, c6456, in6456_1, in6456_2, c3312);
    wire[0:0] s6457, in6457_1, in6457_2;
    wire c6457;
    assign in6457_1 = {c3316};
    assign in6457_2 = {c3317};
    Full_Adder FA_6457(s6457, c6457, in6457_1, in6457_2, c3315);
    wire[0:0] s6458, in6458_1, in6458_2;
    wire c6458;
    assign in6458_1 = {c3319};
    assign in6458_2 = {c3320};
    Full_Adder FA_6458(s6458, c6458, in6458_1, in6458_2, c3318);
    wire[0:0] s6459, in6459_1, in6459_2;
    wire c6459;
    assign in6459_1 = {c3322};
    assign in6459_2 = {c3323};
    Full_Adder FA_6459(s6459, c6459, in6459_1, in6459_2, c3321);
    wire[0:0] s6460, in6460_1, in6460_2;
    wire c6460;
    assign in6460_1 = {c3325};
    assign in6460_2 = {c3326};
    Full_Adder FA_6460(s6460, c6460, in6460_1, in6460_2, c3324);
    wire[0:0] s6461, in6461_1, in6461_2;
    wire c6461;
    assign in6461_1 = {c3328};
    assign in6461_2 = {c3329};
    Full_Adder FA_6461(s6461, c6461, in6461_1, in6461_2, c3327);
    wire[0:0] s6462, in6462_1, in6462_2;
    wire c6462;
    assign in6462_1 = {c3331};
    assign in6462_2 = {c3332};
    Full_Adder FA_6462(s6462, c6462, in6462_1, in6462_2, c3330);
    wire[0:0] s6463, in6463_1, in6463_2;
    wire c6463;
    assign in6463_1 = {s3334[0]};
    assign in6463_2 = {s3335[0]};
    Full_Adder FA_6463(s6463, c6463, in6463_1, in6463_2, s3333[0]);
    wire[0:0] s6464, in6464_1, in6464_2;
    wire c6464;
    assign in6464_1 = {s3337[0]};
    assign in6464_2 = {s3338[0]};
    Full_Adder FA_6464(s6464, c6464, in6464_1, in6464_2, s3336[0]);
    wire[0:0] s6465, in6465_1, in6465_2;
    wire c6465;
    assign in6465_1 = {s3340[0]};
    assign in6465_2 = {s3341[0]};
    Full_Adder FA_6465(s6465, c6465, in6465_1, in6465_2, s3339[0]);
    wire[0:0] s6466, in6466_1, in6466_2;
    wire c6466;
    assign in6466_1 = {s3343[0]};
    assign in6466_2 = {s3344[0]};
    Full_Adder FA_6466(s6466, c6466, in6466_1, in6466_2, s3342[0]);
    wire[0:0] s6467, in6467_1, in6467_2;
    wire c6467;
    assign in6467_1 = {s3346[0]};
    assign in6467_2 = {s3347[0]};
    Full_Adder FA_6467(s6467, c6467, in6467_1, in6467_2, s3345[0]);
    wire[0:0] s6468, in6468_1, in6468_2;
    wire c6468;
    assign in6468_1 = {s3349[0]};
    assign in6468_2 = {s3350[0]};
    Full_Adder FA_6468(s6468, c6468, in6468_1, in6468_2, s3348[0]);
    wire[0:0] s6469, in6469_1, in6469_2;
    wire c6469;
    assign in6469_1 = {s3352[0]};
    assign in6469_2 = {s3353[0]};
    Full_Adder FA_6469(s6469, c6469, in6469_1, in6469_2, s3351[0]);
    wire[0:0] s6470, in6470_1, in6470_2;
    wire c6470;
    assign in6470_1 = {s3355[0]};
    assign in6470_2 = {s3356[0]};
    Full_Adder FA_6470(s6470, c6470, in6470_1, in6470_2, s3354[0]);
    wire[0:0] s6471, in6471_1, in6471_2;
    wire c6471;
    assign in6471_1 = {s3358[0]};
    assign in6471_2 = {s3359[0]};
    Full_Adder FA_6471(s6471, c6471, in6471_1, in6471_2, s3357[0]);
    wire[0:0] s6472, in6472_1, in6472_2;
    wire c6472;
    assign in6472_1 = {s903[0]};
    assign in6472_2 = {c3333};
    Full_Adder FA_6472(s6472, c6472, in6472_1, in6472_2, s902[0]);
    wire[0:0] s6473, in6473_1, in6473_2;
    wire c6473;
    assign in6473_1 = {c3335};
    assign in6473_2 = {c3336};
    Full_Adder FA_6473(s6473, c6473, in6473_1, in6473_2, c3334);
    wire[0:0] s6474, in6474_1, in6474_2;
    wire c6474;
    assign in6474_1 = {c3338};
    assign in6474_2 = {c3339};
    Full_Adder FA_6474(s6474, c6474, in6474_1, in6474_2, c3337);
    wire[0:0] s6475, in6475_1, in6475_2;
    wire c6475;
    assign in6475_1 = {c3341};
    assign in6475_2 = {c3342};
    Full_Adder FA_6475(s6475, c6475, in6475_1, in6475_2, c3340);
    wire[0:0] s6476, in6476_1, in6476_2;
    wire c6476;
    assign in6476_1 = {c3344};
    assign in6476_2 = {c3345};
    Full_Adder FA_6476(s6476, c6476, in6476_1, in6476_2, c3343);
    wire[0:0] s6477, in6477_1, in6477_2;
    wire c6477;
    assign in6477_1 = {c3347};
    assign in6477_2 = {c3348};
    Full_Adder FA_6477(s6477, c6477, in6477_1, in6477_2, c3346);
    wire[0:0] s6478, in6478_1, in6478_2;
    wire c6478;
    assign in6478_1 = {c3350};
    assign in6478_2 = {c3351};
    Full_Adder FA_6478(s6478, c6478, in6478_1, in6478_2, c3349);
    wire[0:0] s6479, in6479_1, in6479_2;
    wire c6479;
    assign in6479_1 = {c3353};
    assign in6479_2 = {c3354};
    Full_Adder FA_6479(s6479, c6479, in6479_1, in6479_2, c3352);
    wire[0:0] s6480, in6480_1, in6480_2;
    wire c6480;
    assign in6480_1 = {c3356};
    assign in6480_2 = {c3357};
    Full_Adder FA_6480(s6480, c6480, in6480_1, in6480_2, c3355);
    wire[0:0] s6481, in6481_1, in6481_2;
    wire c6481;
    assign in6481_1 = {c3359};
    assign in6481_2 = {c3360};
    Full_Adder FA_6481(s6481, c6481, in6481_1, in6481_2, c3358);
    wire[0:0] s6482, in6482_1, in6482_2;
    wire c6482;
    assign in6482_1 = {s3362[0]};
    assign in6482_2 = {s3363[0]};
    Full_Adder FA_6482(s6482, c6482, in6482_1, in6482_2, s3361[0]);
    wire[0:0] s6483, in6483_1, in6483_2;
    wire c6483;
    assign in6483_1 = {s3365[0]};
    assign in6483_2 = {s3366[0]};
    Full_Adder FA_6483(s6483, c6483, in6483_1, in6483_2, s3364[0]);
    wire[0:0] s6484, in6484_1, in6484_2;
    wire c6484;
    assign in6484_1 = {s3368[0]};
    assign in6484_2 = {s3369[0]};
    Full_Adder FA_6484(s6484, c6484, in6484_1, in6484_2, s3367[0]);
    wire[0:0] s6485, in6485_1, in6485_2;
    wire c6485;
    assign in6485_1 = {s3371[0]};
    assign in6485_2 = {s3372[0]};
    Full_Adder FA_6485(s6485, c6485, in6485_1, in6485_2, s3370[0]);
    wire[0:0] s6486, in6486_1, in6486_2;
    wire c6486;
    assign in6486_1 = {s3374[0]};
    assign in6486_2 = {s3375[0]};
    Full_Adder FA_6486(s6486, c6486, in6486_1, in6486_2, s3373[0]);
    wire[0:0] s6487, in6487_1, in6487_2;
    wire c6487;
    assign in6487_1 = {s3377[0]};
    assign in6487_2 = {s3378[0]};
    Full_Adder FA_6487(s6487, c6487, in6487_1, in6487_2, s3376[0]);
    wire[0:0] s6488, in6488_1, in6488_2;
    wire c6488;
    assign in6488_1 = {s3380[0]};
    assign in6488_2 = {s3381[0]};
    Full_Adder FA_6488(s6488, c6488, in6488_1, in6488_2, s3379[0]);
    wire[0:0] s6489, in6489_1, in6489_2;
    wire c6489;
    assign in6489_1 = {s3383[0]};
    assign in6489_2 = {s3384[0]};
    Full_Adder FA_6489(s6489, c6489, in6489_1, in6489_2, s3382[0]);
    wire[0:0] s6490, in6490_1, in6490_2;
    wire c6490;
    assign in6490_1 = {s3386[0]};
    assign in6490_2 = {s3387[0]};
    Full_Adder FA_6490(s6490, c6490, in6490_1, in6490_2, s3385[0]);
    wire[0:0] s6491, in6491_1, in6491_2;
    wire c6491;
    assign in6491_1 = {s945[0]};
    assign in6491_2 = {c3361};
    Full_Adder FA_6491(s6491, c6491, in6491_1, in6491_2, s944[0]);
    wire[0:0] s6492, in6492_1, in6492_2;
    wire c6492;
    assign in6492_1 = {c3363};
    assign in6492_2 = {c3364};
    Full_Adder FA_6492(s6492, c6492, in6492_1, in6492_2, c3362);
    wire[0:0] s6493, in6493_1, in6493_2;
    wire c6493;
    assign in6493_1 = {c3366};
    assign in6493_2 = {c3367};
    Full_Adder FA_6493(s6493, c6493, in6493_1, in6493_2, c3365);
    wire[0:0] s6494, in6494_1, in6494_2;
    wire c6494;
    assign in6494_1 = {c3369};
    assign in6494_2 = {c3370};
    Full_Adder FA_6494(s6494, c6494, in6494_1, in6494_2, c3368);
    wire[0:0] s6495, in6495_1, in6495_2;
    wire c6495;
    assign in6495_1 = {c3372};
    assign in6495_2 = {c3373};
    Full_Adder FA_6495(s6495, c6495, in6495_1, in6495_2, c3371);
    wire[0:0] s6496, in6496_1, in6496_2;
    wire c6496;
    assign in6496_1 = {c3375};
    assign in6496_2 = {c3376};
    Full_Adder FA_6496(s6496, c6496, in6496_1, in6496_2, c3374);
    wire[0:0] s6497, in6497_1, in6497_2;
    wire c6497;
    assign in6497_1 = {c3378};
    assign in6497_2 = {c3379};
    Full_Adder FA_6497(s6497, c6497, in6497_1, in6497_2, c3377);
    wire[0:0] s6498, in6498_1, in6498_2;
    wire c6498;
    assign in6498_1 = {c3381};
    assign in6498_2 = {c3382};
    Full_Adder FA_6498(s6498, c6498, in6498_1, in6498_2, c3380);
    wire[0:0] s6499, in6499_1, in6499_2;
    wire c6499;
    assign in6499_1 = {c3384};
    assign in6499_2 = {c3385};
    Full_Adder FA_6499(s6499, c6499, in6499_1, in6499_2, c3383);
    wire[0:0] s6500, in6500_1, in6500_2;
    wire c6500;
    assign in6500_1 = {c3387};
    assign in6500_2 = {c3388};
    Full_Adder FA_6500(s6500, c6500, in6500_1, in6500_2, c3386);
    wire[0:0] s6501, in6501_1, in6501_2;
    wire c6501;
    assign in6501_1 = {s3390[0]};
    assign in6501_2 = {s3391[0]};
    Full_Adder FA_6501(s6501, c6501, in6501_1, in6501_2, s3389[0]);
    wire[0:0] s6502, in6502_1, in6502_2;
    wire c6502;
    assign in6502_1 = {s3393[0]};
    assign in6502_2 = {s3394[0]};
    Full_Adder FA_6502(s6502, c6502, in6502_1, in6502_2, s3392[0]);
    wire[0:0] s6503, in6503_1, in6503_2;
    wire c6503;
    assign in6503_1 = {s3396[0]};
    assign in6503_2 = {s3397[0]};
    Full_Adder FA_6503(s6503, c6503, in6503_1, in6503_2, s3395[0]);
    wire[0:0] s6504, in6504_1, in6504_2;
    wire c6504;
    assign in6504_1 = {s3399[0]};
    assign in6504_2 = {s3400[0]};
    Full_Adder FA_6504(s6504, c6504, in6504_1, in6504_2, s3398[0]);
    wire[0:0] s6505, in6505_1, in6505_2;
    wire c6505;
    assign in6505_1 = {s3402[0]};
    assign in6505_2 = {s3403[0]};
    Full_Adder FA_6505(s6505, c6505, in6505_1, in6505_2, s3401[0]);
    wire[0:0] s6506, in6506_1, in6506_2;
    wire c6506;
    assign in6506_1 = {s3405[0]};
    assign in6506_2 = {s3406[0]};
    Full_Adder FA_6506(s6506, c6506, in6506_1, in6506_2, s3404[0]);
    wire[0:0] s6507, in6507_1, in6507_2;
    wire c6507;
    assign in6507_1 = {s3408[0]};
    assign in6507_2 = {s3409[0]};
    Full_Adder FA_6507(s6507, c6507, in6507_1, in6507_2, s3407[0]);
    wire[0:0] s6508, in6508_1, in6508_2;
    wire c6508;
    assign in6508_1 = {s3411[0]};
    assign in6508_2 = {s3412[0]};
    Full_Adder FA_6508(s6508, c6508, in6508_1, in6508_2, s3410[0]);
    wire[0:0] s6509, in6509_1, in6509_2;
    wire c6509;
    assign in6509_1 = {s3414[0]};
    assign in6509_2 = {s3415[0]};
    Full_Adder FA_6509(s6509, c6509, in6509_1, in6509_2, s3413[0]);
    wire[0:0] s6510, in6510_1, in6510_2;
    wire c6510;
    assign in6510_1 = {s986[0]};
    assign in6510_2 = {c3389};
    Full_Adder FA_6510(s6510, c6510, in6510_1, in6510_2, s985[0]);
    wire[0:0] s6511, in6511_1, in6511_2;
    wire c6511;
    assign in6511_1 = {c3391};
    assign in6511_2 = {c3392};
    Full_Adder FA_6511(s6511, c6511, in6511_1, in6511_2, c3390);
    wire[0:0] s6512, in6512_1, in6512_2;
    wire c6512;
    assign in6512_1 = {c3394};
    assign in6512_2 = {c3395};
    Full_Adder FA_6512(s6512, c6512, in6512_1, in6512_2, c3393);
    wire[0:0] s6513, in6513_1, in6513_2;
    wire c6513;
    assign in6513_1 = {c3397};
    assign in6513_2 = {c3398};
    Full_Adder FA_6513(s6513, c6513, in6513_1, in6513_2, c3396);
    wire[0:0] s6514, in6514_1, in6514_2;
    wire c6514;
    assign in6514_1 = {c3400};
    assign in6514_2 = {c3401};
    Full_Adder FA_6514(s6514, c6514, in6514_1, in6514_2, c3399);
    wire[0:0] s6515, in6515_1, in6515_2;
    wire c6515;
    assign in6515_1 = {c3403};
    assign in6515_2 = {c3404};
    Full_Adder FA_6515(s6515, c6515, in6515_1, in6515_2, c3402);
    wire[0:0] s6516, in6516_1, in6516_2;
    wire c6516;
    assign in6516_1 = {c3406};
    assign in6516_2 = {c3407};
    Full_Adder FA_6516(s6516, c6516, in6516_1, in6516_2, c3405);
    wire[0:0] s6517, in6517_1, in6517_2;
    wire c6517;
    assign in6517_1 = {c3409};
    assign in6517_2 = {c3410};
    Full_Adder FA_6517(s6517, c6517, in6517_1, in6517_2, c3408);
    wire[0:0] s6518, in6518_1, in6518_2;
    wire c6518;
    assign in6518_1 = {c3412};
    assign in6518_2 = {c3413};
    Full_Adder FA_6518(s6518, c6518, in6518_1, in6518_2, c3411);
    wire[0:0] s6519, in6519_1, in6519_2;
    wire c6519;
    assign in6519_1 = {c3415};
    assign in6519_2 = {c3416};
    Full_Adder FA_6519(s6519, c6519, in6519_1, in6519_2, c3414);
    wire[0:0] s6520, in6520_1, in6520_2;
    wire c6520;
    assign in6520_1 = {s3418[0]};
    assign in6520_2 = {s3419[0]};
    Full_Adder FA_6520(s6520, c6520, in6520_1, in6520_2, s3417[0]);
    wire[0:0] s6521, in6521_1, in6521_2;
    wire c6521;
    assign in6521_1 = {s3421[0]};
    assign in6521_2 = {s3422[0]};
    Full_Adder FA_6521(s6521, c6521, in6521_1, in6521_2, s3420[0]);
    wire[0:0] s6522, in6522_1, in6522_2;
    wire c6522;
    assign in6522_1 = {s3424[0]};
    assign in6522_2 = {s3425[0]};
    Full_Adder FA_6522(s6522, c6522, in6522_1, in6522_2, s3423[0]);
    wire[0:0] s6523, in6523_1, in6523_2;
    wire c6523;
    assign in6523_1 = {s3427[0]};
    assign in6523_2 = {s3428[0]};
    Full_Adder FA_6523(s6523, c6523, in6523_1, in6523_2, s3426[0]);
    wire[0:0] s6524, in6524_1, in6524_2;
    wire c6524;
    assign in6524_1 = {s3430[0]};
    assign in6524_2 = {s3431[0]};
    Full_Adder FA_6524(s6524, c6524, in6524_1, in6524_2, s3429[0]);
    wire[0:0] s6525, in6525_1, in6525_2;
    wire c6525;
    assign in6525_1 = {s3433[0]};
    assign in6525_2 = {s3434[0]};
    Full_Adder FA_6525(s6525, c6525, in6525_1, in6525_2, s3432[0]);
    wire[0:0] s6526, in6526_1, in6526_2;
    wire c6526;
    assign in6526_1 = {s3436[0]};
    assign in6526_2 = {s3437[0]};
    Full_Adder FA_6526(s6526, c6526, in6526_1, in6526_2, s3435[0]);
    wire[0:0] s6527, in6527_1, in6527_2;
    wire c6527;
    assign in6527_1 = {s3439[0]};
    assign in6527_2 = {s3440[0]};
    Full_Adder FA_6527(s6527, c6527, in6527_1, in6527_2, s3438[0]);
    wire[0:0] s6528, in6528_1, in6528_2;
    wire c6528;
    assign in6528_1 = {s3442[0]};
    assign in6528_2 = {s3443[0]};
    Full_Adder FA_6528(s6528, c6528, in6528_1, in6528_2, s3441[0]);
    wire[0:0] s6529, in6529_1, in6529_2;
    wire c6529;
    assign in6529_1 = {s1026[0]};
    assign in6529_2 = {c3417};
    Full_Adder FA_6529(s6529, c6529, in6529_1, in6529_2, s1025[0]);
    wire[0:0] s6530, in6530_1, in6530_2;
    wire c6530;
    assign in6530_1 = {c3419};
    assign in6530_2 = {c3420};
    Full_Adder FA_6530(s6530, c6530, in6530_1, in6530_2, c3418);
    wire[0:0] s6531, in6531_1, in6531_2;
    wire c6531;
    assign in6531_1 = {c3422};
    assign in6531_2 = {c3423};
    Full_Adder FA_6531(s6531, c6531, in6531_1, in6531_2, c3421);
    wire[0:0] s6532, in6532_1, in6532_2;
    wire c6532;
    assign in6532_1 = {c3425};
    assign in6532_2 = {c3426};
    Full_Adder FA_6532(s6532, c6532, in6532_1, in6532_2, c3424);
    wire[0:0] s6533, in6533_1, in6533_2;
    wire c6533;
    assign in6533_1 = {c3428};
    assign in6533_2 = {c3429};
    Full_Adder FA_6533(s6533, c6533, in6533_1, in6533_2, c3427);
    wire[0:0] s6534, in6534_1, in6534_2;
    wire c6534;
    assign in6534_1 = {c3431};
    assign in6534_2 = {c3432};
    Full_Adder FA_6534(s6534, c6534, in6534_1, in6534_2, c3430);
    wire[0:0] s6535, in6535_1, in6535_2;
    wire c6535;
    assign in6535_1 = {c3434};
    assign in6535_2 = {c3435};
    Full_Adder FA_6535(s6535, c6535, in6535_1, in6535_2, c3433);
    wire[0:0] s6536, in6536_1, in6536_2;
    wire c6536;
    assign in6536_1 = {c3437};
    assign in6536_2 = {c3438};
    Full_Adder FA_6536(s6536, c6536, in6536_1, in6536_2, c3436);
    wire[0:0] s6537, in6537_1, in6537_2;
    wire c6537;
    assign in6537_1 = {c3440};
    assign in6537_2 = {c3441};
    Full_Adder FA_6537(s6537, c6537, in6537_1, in6537_2, c3439);
    wire[0:0] s6538, in6538_1, in6538_2;
    wire c6538;
    assign in6538_1 = {c3443};
    assign in6538_2 = {c3444};
    Full_Adder FA_6538(s6538, c6538, in6538_1, in6538_2, c3442);
    wire[0:0] s6539, in6539_1, in6539_2;
    wire c6539;
    assign in6539_1 = {s3446[0]};
    assign in6539_2 = {s3447[0]};
    Full_Adder FA_6539(s6539, c6539, in6539_1, in6539_2, s3445[0]);
    wire[0:0] s6540, in6540_1, in6540_2;
    wire c6540;
    assign in6540_1 = {s3449[0]};
    assign in6540_2 = {s3450[0]};
    Full_Adder FA_6540(s6540, c6540, in6540_1, in6540_2, s3448[0]);
    wire[0:0] s6541, in6541_1, in6541_2;
    wire c6541;
    assign in6541_1 = {s3452[0]};
    assign in6541_2 = {s3453[0]};
    Full_Adder FA_6541(s6541, c6541, in6541_1, in6541_2, s3451[0]);
    wire[0:0] s6542, in6542_1, in6542_2;
    wire c6542;
    assign in6542_1 = {s3455[0]};
    assign in6542_2 = {s3456[0]};
    Full_Adder FA_6542(s6542, c6542, in6542_1, in6542_2, s3454[0]);
    wire[0:0] s6543, in6543_1, in6543_2;
    wire c6543;
    assign in6543_1 = {s3458[0]};
    assign in6543_2 = {s3459[0]};
    Full_Adder FA_6543(s6543, c6543, in6543_1, in6543_2, s3457[0]);
    wire[0:0] s6544, in6544_1, in6544_2;
    wire c6544;
    assign in6544_1 = {s3461[0]};
    assign in6544_2 = {s3462[0]};
    Full_Adder FA_6544(s6544, c6544, in6544_1, in6544_2, s3460[0]);
    wire[0:0] s6545, in6545_1, in6545_2;
    wire c6545;
    assign in6545_1 = {s3464[0]};
    assign in6545_2 = {s3465[0]};
    Full_Adder FA_6545(s6545, c6545, in6545_1, in6545_2, s3463[0]);
    wire[0:0] s6546, in6546_1, in6546_2;
    wire c6546;
    assign in6546_1 = {s3467[0]};
    assign in6546_2 = {s3468[0]};
    Full_Adder FA_6546(s6546, c6546, in6546_1, in6546_2, s3466[0]);
    wire[0:0] s6547, in6547_1, in6547_2;
    wire c6547;
    assign in6547_1 = {s3470[0]};
    assign in6547_2 = {s3471[0]};
    Full_Adder FA_6547(s6547, c6547, in6547_1, in6547_2, s3469[0]);
    wire[0:0] s6548, in6548_1, in6548_2;
    wire c6548;
    assign in6548_1 = {s1065[0]};
    assign in6548_2 = {c3445};
    Full_Adder FA_6548(s6548, c6548, in6548_1, in6548_2, s1064[0]);
    wire[0:0] s6549, in6549_1, in6549_2;
    wire c6549;
    assign in6549_1 = {c3447};
    assign in6549_2 = {c3448};
    Full_Adder FA_6549(s6549, c6549, in6549_1, in6549_2, c3446);
    wire[0:0] s6550, in6550_1, in6550_2;
    wire c6550;
    assign in6550_1 = {c3450};
    assign in6550_2 = {c3451};
    Full_Adder FA_6550(s6550, c6550, in6550_1, in6550_2, c3449);
    wire[0:0] s6551, in6551_1, in6551_2;
    wire c6551;
    assign in6551_1 = {c3453};
    assign in6551_2 = {c3454};
    Full_Adder FA_6551(s6551, c6551, in6551_1, in6551_2, c3452);
    wire[0:0] s6552, in6552_1, in6552_2;
    wire c6552;
    assign in6552_1 = {c3456};
    assign in6552_2 = {c3457};
    Full_Adder FA_6552(s6552, c6552, in6552_1, in6552_2, c3455);
    wire[0:0] s6553, in6553_1, in6553_2;
    wire c6553;
    assign in6553_1 = {c3459};
    assign in6553_2 = {c3460};
    Full_Adder FA_6553(s6553, c6553, in6553_1, in6553_2, c3458);
    wire[0:0] s6554, in6554_1, in6554_2;
    wire c6554;
    assign in6554_1 = {c3462};
    assign in6554_2 = {c3463};
    Full_Adder FA_6554(s6554, c6554, in6554_1, in6554_2, c3461);
    wire[0:0] s6555, in6555_1, in6555_2;
    wire c6555;
    assign in6555_1 = {c3465};
    assign in6555_2 = {c3466};
    Full_Adder FA_6555(s6555, c6555, in6555_1, in6555_2, c3464);
    wire[0:0] s6556, in6556_1, in6556_2;
    wire c6556;
    assign in6556_1 = {c3468};
    assign in6556_2 = {c3469};
    Full_Adder FA_6556(s6556, c6556, in6556_1, in6556_2, c3467);
    wire[0:0] s6557, in6557_1, in6557_2;
    wire c6557;
    assign in6557_1 = {c3471};
    assign in6557_2 = {c3472};
    Full_Adder FA_6557(s6557, c6557, in6557_1, in6557_2, c3470);
    wire[0:0] s6558, in6558_1, in6558_2;
    wire c6558;
    assign in6558_1 = {s3474[0]};
    assign in6558_2 = {s3475[0]};
    Full_Adder FA_6558(s6558, c6558, in6558_1, in6558_2, s3473[0]);
    wire[0:0] s6559, in6559_1, in6559_2;
    wire c6559;
    assign in6559_1 = {s3477[0]};
    assign in6559_2 = {s3478[0]};
    Full_Adder FA_6559(s6559, c6559, in6559_1, in6559_2, s3476[0]);
    wire[0:0] s6560, in6560_1, in6560_2;
    wire c6560;
    assign in6560_1 = {s3480[0]};
    assign in6560_2 = {s3481[0]};
    Full_Adder FA_6560(s6560, c6560, in6560_1, in6560_2, s3479[0]);
    wire[0:0] s6561, in6561_1, in6561_2;
    wire c6561;
    assign in6561_1 = {s3483[0]};
    assign in6561_2 = {s3484[0]};
    Full_Adder FA_6561(s6561, c6561, in6561_1, in6561_2, s3482[0]);
    wire[0:0] s6562, in6562_1, in6562_2;
    wire c6562;
    assign in6562_1 = {s3486[0]};
    assign in6562_2 = {s3487[0]};
    Full_Adder FA_6562(s6562, c6562, in6562_1, in6562_2, s3485[0]);
    wire[0:0] s6563, in6563_1, in6563_2;
    wire c6563;
    assign in6563_1 = {s3489[0]};
    assign in6563_2 = {s3490[0]};
    Full_Adder FA_6563(s6563, c6563, in6563_1, in6563_2, s3488[0]);
    wire[0:0] s6564, in6564_1, in6564_2;
    wire c6564;
    assign in6564_1 = {s3492[0]};
    assign in6564_2 = {s3493[0]};
    Full_Adder FA_6564(s6564, c6564, in6564_1, in6564_2, s3491[0]);
    wire[0:0] s6565, in6565_1, in6565_2;
    wire c6565;
    assign in6565_1 = {s3495[0]};
    assign in6565_2 = {s3496[0]};
    Full_Adder FA_6565(s6565, c6565, in6565_1, in6565_2, s3494[0]);
    wire[0:0] s6566, in6566_1, in6566_2;
    wire c6566;
    assign in6566_1 = {s3498[0]};
    assign in6566_2 = {s3499[0]};
    Full_Adder FA_6566(s6566, c6566, in6566_1, in6566_2, s3497[0]);
    wire[0:0] s6567, in6567_1, in6567_2;
    wire c6567;
    assign in6567_1 = {s1103[0]};
    assign in6567_2 = {c3473};
    Full_Adder FA_6567(s6567, c6567, in6567_1, in6567_2, s1102[0]);
    wire[0:0] s6568, in6568_1, in6568_2;
    wire c6568;
    assign in6568_1 = {c3475};
    assign in6568_2 = {c3476};
    Full_Adder FA_6568(s6568, c6568, in6568_1, in6568_2, c3474);
    wire[0:0] s6569, in6569_1, in6569_2;
    wire c6569;
    assign in6569_1 = {c3478};
    assign in6569_2 = {c3479};
    Full_Adder FA_6569(s6569, c6569, in6569_1, in6569_2, c3477);
    wire[0:0] s6570, in6570_1, in6570_2;
    wire c6570;
    assign in6570_1 = {c3481};
    assign in6570_2 = {c3482};
    Full_Adder FA_6570(s6570, c6570, in6570_1, in6570_2, c3480);
    wire[0:0] s6571, in6571_1, in6571_2;
    wire c6571;
    assign in6571_1 = {c3484};
    assign in6571_2 = {c3485};
    Full_Adder FA_6571(s6571, c6571, in6571_1, in6571_2, c3483);
    wire[0:0] s6572, in6572_1, in6572_2;
    wire c6572;
    assign in6572_1 = {c3487};
    assign in6572_2 = {c3488};
    Full_Adder FA_6572(s6572, c6572, in6572_1, in6572_2, c3486);
    wire[0:0] s6573, in6573_1, in6573_2;
    wire c6573;
    assign in6573_1 = {c3490};
    assign in6573_2 = {c3491};
    Full_Adder FA_6573(s6573, c6573, in6573_1, in6573_2, c3489);
    wire[0:0] s6574, in6574_1, in6574_2;
    wire c6574;
    assign in6574_1 = {c3493};
    assign in6574_2 = {c3494};
    Full_Adder FA_6574(s6574, c6574, in6574_1, in6574_2, c3492);
    wire[0:0] s6575, in6575_1, in6575_2;
    wire c6575;
    assign in6575_1 = {c3496};
    assign in6575_2 = {c3497};
    Full_Adder FA_6575(s6575, c6575, in6575_1, in6575_2, c3495);
    wire[0:0] s6576, in6576_1, in6576_2;
    wire c6576;
    assign in6576_1 = {c3499};
    assign in6576_2 = {c3500};
    Full_Adder FA_6576(s6576, c6576, in6576_1, in6576_2, c3498);
    wire[0:0] s6577, in6577_1, in6577_2;
    wire c6577;
    assign in6577_1 = {s3502[0]};
    assign in6577_2 = {s3503[0]};
    Full_Adder FA_6577(s6577, c6577, in6577_1, in6577_2, s3501[0]);
    wire[0:0] s6578, in6578_1, in6578_2;
    wire c6578;
    assign in6578_1 = {s3505[0]};
    assign in6578_2 = {s3506[0]};
    Full_Adder FA_6578(s6578, c6578, in6578_1, in6578_2, s3504[0]);
    wire[0:0] s6579, in6579_1, in6579_2;
    wire c6579;
    assign in6579_1 = {s3508[0]};
    assign in6579_2 = {s3509[0]};
    Full_Adder FA_6579(s6579, c6579, in6579_1, in6579_2, s3507[0]);
    wire[0:0] s6580, in6580_1, in6580_2;
    wire c6580;
    assign in6580_1 = {s3511[0]};
    assign in6580_2 = {s3512[0]};
    Full_Adder FA_6580(s6580, c6580, in6580_1, in6580_2, s3510[0]);
    wire[0:0] s6581, in6581_1, in6581_2;
    wire c6581;
    assign in6581_1 = {s3514[0]};
    assign in6581_2 = {s3515[0]};
    Full_Adder FA_6581(s6581, c6581, in6581_1, in6581_2, s3513[0]);
    wire[0:0] s6582, in6582_1, in6582_2;
    wire c6582;
    assign in6582_1 = {s3517[0]};
    assign in6582_2 = {s3518[0]};
    Full_Adder FA_6582(s6582, c6582, in6582_1, in6582_2, s3516[0]);
    wire[0:0] s6583, in6583_1, in6583_2;
    wire c6583;
    assign in6583_1 = {s3520[0]};
    assign in6583_2 = {s3521[0]};
    Full_Adder FA_6583(s6583, c6583, in6583_1, in6583_2, s3519[0]);
    wire[0:0] s6584, in6584_1, in6584_2;
    wire c6584;
    assign in6584_1 = {s3523[0]};
    assign in6584_2 = {s3524[0]};
    Full_Adder FA_6584(s6584, c6584, in6584_1, in6584_2, s3522[0]);
    wire[0:0] s6585, in6585_1, in6585_2;
    wire c6585;
    assign in6585_1 = {s3526[0]};
    assign in6585_2 = {s3527[0]};
    Full_Adder FA_6585(s6585, c6585, in6585_1, in6585_2, s3525[0]);
    wire[0:0] s6586, in6586_1, in6586_2;
    wire c6586;
    assign in6586_1 = {s1140[0]};
    assign in6586_2 = {c3501};
    Full_Adder FA_6586(s6586, c6586, in6586_1, in6586_2, s1139[0]);
    wire[0:0] s6587, in6587_1, in6587_2;
    wire c6587;
    assign in6587_1 = {c3503};
    assign in6587_2 = {c3504};
    Full_Adder FA_6587(s6587, c6587, in6587_1, in6587_2, c3502);
    wire[0:0] s6588, in6588_1, in6588_2;
    wire c6588;
    assign in6588_1 = {c3506};
    assign in6588_2 = {c3507};
    Full_Adder FA_6588(s6588, c6588, in6588_1, in6588_2, c3505);
    wire[0:0] s6589, in6589_1, in6589_2;
    wire c6589;
    assign in6589_1 = {c3509};
    assign in6589_2 = {c3510};
    Full_Adder FA_6589(s6589, c6589, in6589_1, in6589_2, c3508);
    wire[0:0] s6590, in6590_1, in6590_2;
    wire c6590;
    assign in6590_1 = {c3512};
    assign in6590_2 = {c3513};
    Full_Adder FA_6590(s6590, c6590, in6590_1, in6590_2, c3511);
    wire[0:0] s6591, in6591_1, in6591_2;
    wire c6591;
    assign in6591_1 = {c3515};
    assign in6591_2 = {c3516};
    Full_Adder FA_6591(s6591, c6591, in6591_1, in6591_2, c3514);
    wire[0:0] s6592, in6592_1, in6592_2;
    wire c6592;
    assign in6592_1 = {c3518};
    assign in6592_2 = {c3519};
    Full_Adder FA_6592(s6592, c6592, in6592_1, in6592_2, c3517);
    wire[0:0] s6593, in6593_1, in6593_2;
    wire c6593;
    assign in6593_1 = {c3521};
    assign in6593_2 = {c3522};
    Full_Adder FA_6593(s6593, c6593, in6593_1, in6593_2, c3520);
    wire[0:0] s6594, in6594_1, in6594_2;
    wire c6594;
    assign in6594_1 = {c3524};
    assign in6594_2 = {c3525};
    Full_Adder FA_6594(s6594, c6594, in6594_1, in6594_2, c3523);
    wire[0:0] s6595, in6595_1, in6595_2;
    wire c6595;
    assign in6595_1 = {c3527};
    assign in6595_2 = {c3528};
    Full_Adder FA_6595(s6595, c6595, in6595_1, in6595_2, c3526);
    wire[0:0] s6596, in6596_1, in6596_2;
    wire c6596;
    assign in6596_1 = {s3530[0]};
    assign in6596_2 = {s3531[0]};
    Full_Adder FA_6596(s6596, c6596, in6596_1, in6596_2, s3529[0]);
    wire[0:0] s6597, in6597_1, in6597_2;
    wire c6597;
    assign in6597_1 = {s3533[0]};
    assign in6597_2 = {s3534[0]};
    Full_Adder FA_6597(s6597, c6597, in6597_1, in6597_2, s3532[0]);
    wire[0:0] s6598, in6598_1, in6598_2;
    wire c6598;
    assign in6598_1 = {s3536[0]};
    assign in6598_2 = {s3537[0]};
    Full_Adder FA_6598(s6598, c6598, in6598_1, in6598_2, s3535[0]);
    wire[0:0] s6599, in6599_1, in6599_2;
    wire c6599;
    assign in6599_1 = {s3539[0]};
    assign in6599_2 = {s3540[0]};
    Full_Adder FA_6599(s6599, c6599, in6599_1, in6599_2, s3538[0]);
    wire[0:0] s6600, in6600_1, in6600_2;
    wire c6600;
    assign in6600_1 = {s3542[0]};
    assign in6600_2 = {s3543[0]};
    Full_Adder FA_6600(s6600, c6600, in6600_1, in6600_2, s3541[0]);
    wire[0:0] s6601, in6601_1, in6601_2;
    wire c6601;
    assign in6601_1 = {s3545[0]};
    assign in6601_2 = {s3546[0]};
    Full_Adder FA_6601(s6601, c6601, in6601_1, in6601_2, s3544[0]);
    wire[0:0] s6602, in6602_1, in6602_2;
    wire c6602;
    assign in6602_1 = {s3548[0]};
    assign in6602_2 = {s3549[0]};
    Full_Adder FA_6602(s6602, c6602, in6602_1, in6602_2, s3547[0]);
    wire[0:0] s6603, in6603_1, in6603_2;
    wire c6603;
    assign in6603_1 = {s3551[0]};
    assign in6603_2 = {s3552[0]};
    Full_Adder FA_6603(s6603, c6603, in6603_1, in6603_2, s3550[0]);
    wire[0:0] s6604, in6604_1, in6604_2;
    wire c6604;
    assign in6604_1 = {s3554[0]};
    assign in6604_2 = {s3555[0]};
    Full_Adder FA_6604(s6604, c6604, in6604_1, in6604_2, s3553[0]);
    wire[0:0] s6605, in6605_1, in6605_2;
    wire c6605;
    assign in6605_1 = {s1176[0]};
    assign in6605_2 = {c3529};
    Full_Adder FA_6605(s6605, c6605, in6605_1, in6605_2, s1175[0]);
    wire[0:0] s6606, in6606_1, in6606_2;
    wire c6606;
    assign in6606_1 = {c3531};
    assign in6606_2 = {c3532};
    Full_Adder FA_6606(s6606, c6606, in6606_1, in6606_2, c3530);
    wire[0:0] s6607, in6607_1, in6607_2;
    wire c6607;
    assign in6607_1 = {c3534};
    assign in6607_2 = {c3535};
    Full_Adder FA_6607(s6607, c6607, in6607_1, in6607_2, c3533);
    wire[0:0] s6608, in6608_1, in6608_2;
    wire c6608;
    assign in6608_1 = {c3537};
    assign in6608_2 = {c3538};
    Full_Adder FA_6608(s6608, c6608, in6608_1, in6608_2, c3536);
    wire[0:0] s6609, in6609_1, in6609_2;
    wire c6609;
    assign in6609_1 = {c3540};
    assign in6609_2 = {c3541};
    Full_Adder FA_6609(s6609, c6609, in6609_1, in6609_2, c3539);
    wire[0:0] s6610, in6610_1, in6610_2;
    wire c6610;
    assign in6610_1 = {c3543};
    assign in6610_2 = {c3544};
    Full_Adder FA_6610(s6610, c6610, in6610_1, in6610_2, c3542);
    wire[0:0] s6611, in6611_1, in6611_2;
    wire c6611;
    assign in6611_1 = {c3546};
    assign in6611_2 = {c3547};
    Full_Adder FA_6611(s6611, c6611, in6611_1, in6611_2, c3545);
    wire[0:0] s6612, in6612_1, in6612_2;
    wire c6612;
    assign in6612_1 = {c3549};
    assign in6612_2 = {c3550};
    Full_Adder FA_6612(s6612, c6612, in6612_1, in6612_2, c3548);
    wire[0:0] s6613, in6613_1, in6613_2;
    wire c6613;
    assign in6613_1 = {c3552};
    assign in6613_2 = {c3553};
    Full_Adder FA_6613(s6613, c6613, in6613_1, in6613_2, c3551);
    wire[0:0] s6614, in6614_1, in6614_2;
    wire c6614;
    assign in6614_1 = {c3555};
    assign in6614_2 = {c3556};
    Full_Adder FA_6614(s6614, c6614, in6614_1, in6614_2, c3554);
    wire[0:0] s6615, in6615_1, in6615_2;
    wire c6615;
    assign in6615_1 = {s3558[0]};
    assign in6615_2 = {s3559[0]};
    Full_Adder FA_6615(s6615, c6615, in6615_1, in6615_2, s3557[0]);
    wire[0:0] s6616, in6616_1, in6616_2;
    wire c6616;
    assign in6616_1 = {s3561[0]};
    assign in6616_2 = {s3562[0]};
    Full_Adder FA_6616(s6616, c6616, in6616_1, in6616_2, s3560[0]);
    wire[0:0] s6617, in6617_1, in6617_2;
    wire c6617;
    assign in6617_1 = {s3564[0]};
    assign in6617_2 = {s3565[0]};
    Full_Adder FA_6617(s6617, c6617, in6617_1, in6617_2, s3563[0]);
    wire[0:0] s6618, in6618_1, in6618_2;
    wire c6618;
    assign in6618_1 = {s3567[0]};
    assign in6618_2 = {s3568[0]};
    Full_Adder FA_6618(s6618, c6618, in6618_1, in6618_2, s3566[0]);
    wire[0:0] s6619, in6619_1, in6619_2;
    wire c6619;
    assign in6619_1 = {s3570[0]};
    assign in6619_2 = {s3571[0]};
    Full_Adder FA_6619(s6619, c6619, in6619_1, in6619_2, s3569[0]);
    wire[0:0] s6620, in6620_1, in6620_2;
    wire c6620;
    assign in6620_1 = {s3573[0]};
    assign in6620_2 = {s3574[0]};
    Full_Adder FA_6620(s6620, c6620, in6620_1, in6620_2, s3572[0]);
    wire[0:0] s6621, in6621_1, in6621_2;
    wire c6621;
    assign in6621_1 = {s3576[0]};
    assign in6621_2 = {s3577[0]};
    Full_Adder FA_6621(s6621, c6621, in6621_1, in6621_2, s3575[0]);
    wire[0:0] s6622, in6622_1, in6622_2;
    wire c6622;
    assign in6622_1 = {s3579[0]};
    assign in6622_2 = {s3580[0]};
    Full_Adder FA_6622(s6622, c6622, in6622_1, in6622_2, s3578[0]);
    wire[0:0] s6623, in6623_1, in6623_2;
    wire c6623;
    assign in6623_1 = {s3582[0]};
    assign in6623_2 = {s3583[0]};
    Full_Adder FA_6623(s6623, c6623, in6623_1, in6623_2, s3581[0]);
    wire[0:0] s6624, in6624_1, in6624_2;
    wire c6624;
    assign in6624_1 = {s1211[0]};
    assign in6624_2 = {c3557};
    Full_Adder FA_6624(s6624, c6624, in6624_1, in6624_2, s1210[0]);
    wire[0:0] s6625, in6625_1, in6625_2;
    wire c6625;
    assign in6625_1 = {c3559};
    assign in6625_2 = {c3560};
    Full_Adder FA_6625(s6625, c6625, in6625_1, in6625_2, c3558);
    wire[0:0] s6626, in6626_1, in6626_2;
    wire c6626;
    assign in6626_1 = {c3562};
    assign in6626_2 = {c3563};
    Full_Adder FA_6626(s6626, c6626, in6626_1, in6626_2, c3561);
    wire[0:0] s6627, in6627_1, in6627_2;
    wire c6627;
    assign in6627_1 = {c3565};
    assign in6627_2 = {c3566};
    Full_Adder FA_6627(s6627, c6627, in6627_1, in6627_2, c3564);
    wire[0:0] s6628, in6628_1, in6628_2;
    wire c6628;
    assign in6628_1 = {c3568};
    assign in6628_2 = {c3569};
    Full_Adder FA_6628(s6628, c6628, in6628_1, in6628_2, c3567);
    wire[0:0] s6629, in6629_1, in6629_2;
    wire c6629;
    assign in6629_1 = {c3571};
    assign in6629_2 = {c3572};
    Full_Adder FA_6629(s6629, c6629, in6629_1, in6629_2, c3570);
    wire[0:0] s6630, in6630_1, in6630_2;
    wire c6630;
    assign in6630_1 = {c3574};
    assign in6630_2 = {c3575};
    Full_Adder FA_6630(s6630, c6630, in6630_1, in6630_2, c3573);
    wire[0:0] s6631, in6631_1, in6631_2;
    wire c6631;
    assign in6631_1 = {c3577};
    assign in6631_2 = {c3578};
    Full_Adder FA_6631(s6631, c6631, in6631_1, in6631_2, c3576);
    wire[0:0] s6632, in6632_1, in6632_2;
    wire c6632;
    assign in6632_1 = {c3580};
    assign in6632_2 = {c3581};
    Full_Adder FA_6632(s6632, c6632, in6632_1, in6632_2, c3579);
    wire[0:0] s6633, in6633_1, in6633_2;
    wire c6633;
    assign in6633_1 = {c3583};
    assign in6633_2 = {c3584};
    Full_Adder FA_6633(s6633, c6633, in6633_1, in6633_2, c3582);
    wire[0:0] s6634, in6634_1, in6634_2;
    wire c6634;
    assign in6634_1 = {s3586[0]};
    assign in6634_2 = {s3587[0]};
    Full_Adder FA_6634(s6634, c6634, in6634_1, in6634_2, s3585[0]);
    wire[0:0] s6635, in6635_1, in6635_2;
    wire c6635;
    assign in6635_1 = {s3589[0]};
    assign in6635_2 = {s3590[0]};
    Full_Adder FA_6635(s6635, c6635, in6635_1, in6635_2, s3588[0]);
    wire[0:0] s6636, in6636_1, in6636_2;
    wire c6636;
    assign in6636_1 = {s3592[0]};
    assign in6636_2 = {s3593[0]};
    Full_Adder FA_6636(s6636, c6636, in6636_1, in6636_2, s3591[0]);
    wire[0:0] s6637, in6637_1, in6637_2;
    wire c6637;
    assign in6637_1 = {s3595[0]};
    assign in6637_2 = {s3596[0]};
    Full_Adder FA_6637(s6637, c6637, in6637_1, in6637_2, s3594[0]);
    wire[0:0] s6638, in6638_1, in6638_2;
    wire c6638;
    assign in6638_1 = {s3598[0]};
    assign in6638_2 = {s3599[0]};
    Full_Adder FA_6638(s6638, c6638, in6638_1, in6638_2, s3597[0]);
    wire[0:0] s6639, in6639_1, in6639_2;
    wire c6639;
    assign in6639_1 = {s3601[0]};
    assign in6639_2 = {s3602[0]};
    Full_Adder FA_6639(s6639, c6639, in6639_1, in6639_2, s3600[0]);
    wire[0:0] s6640, in6640_1, in6640_2;
    wire c6640;
    assign in6640_1 = {s3604[0]};
    assign in6640_2 = {s3605[0]};
    Full_Adder FA_6640(s6640, c6640, in6640_1, in6640_2, s3603[0]);
    wire[0:0] s6641, in6641_1, in6641_2;
    wire c6641;
    assign in6641_1 = {s3607[0]};
    assign in6641_2 = {s3608[0]};
    Full_Adder FA_6641(s6641, c6641, in6641_1, in6641_2, s3606[0]);
    wire[0:0] s6642, in6642_1, in6642_2;
    wire c6642;
    assign in6642_1 = {s3610[0]};
    assign in6642_2 = {s3611[0]};
    Full_Adder FA_6642(s6642, c6642, in6642_1, in6642_2, s3609[0]);
    wire[0:0] s6643, in6643_1, in6643_2;
    wire c6643;
    assign in6643_1 = {s1245[0]};
    assign in6643_2 = {c3585};
    Full_Adder FA_6643(s6643, c6643, in6643_1, in6643_2, s1244[0]);
    wire[0:0] s6644, in6644_1, in6644_2;
    wire c6644;
    assign in6644_1 = {c3587};
    assign in6644_2 = {c3588};
    Full_Adder FA_6644(s6644, c6644, in6644_1, in6644_2, c3586);
    wire[0:0] s6645, in6645_1, in6645_2;
    wire c6645;
    assign in6645_1 = {c3590};
    assign in6645_2 = {c3591};
    Full_Adder FA_6645(s6645, c6645, in6645_1, in6645_2, c3589);
    wire[0:0] s6646, in6646_1, in6646_2;
    wire c6646;
    assign in6646_1 = {c3593};
    assign in6646_2 = {c3594};
    Full_Adder FA_6646(s6646, c6646, in6646_1, in6646_2, c3592);
    wire[0:0] s6647, in6647_1, in6647_2;
    wire c6647;
    assign in6647_1 = {c3596};
    assign in6647_2 = {c3597};
    Full_Adder FA_6647(s6647, c6647, in6647_1, in6647_2, c3595);
    wire[0:0] s6648, in6648_1, in6648_2;
    wire c6648;
    assign in6648_1 = {c3599};
    assign in6648_2 = {c3600};
    Full_Adder FA_6648(s6648, c6648, in6648_1, in6648_2, c3598);
    wire[0:0] s6649, in6649_1, in6649_2;
    wire c6649;
    assign in6649_1 = {c3602};
    assign in6649_2 = {c3603};
    Full_Adder FA_6649(s6649, c6649, in6649_1, in6649_2, c3601);
    wire[0:0] s6650, in6650_1, in6650_2;
    wire c6650;
    assign in6650_1 = {c3605};
    assign in6650_2 = {c3606};
    Full_Adder FA_6650(s6650, c6650, in6650_1, in6650_2, c3604);
    wire[0:0] s6651, in6651_1, in6651_2;
    wire c6651;
    assign in6651_1 = {c3608};
    assign in6651_2 = {c3609};
    Full_Adder FA_6651(s6651, c6651, in6651_1, in6651_2, c3607);
    wire[0:0] s6652, in6652_1, in6652_2;
    wire c6652;
    assign in6652_1 = {c3611};
    assign in6652_2 = {c3612};
    Full_Adder FA_6652(s6652, c6652, in6652_1, in6652_2, c3610);
    wire[0:0] s6653, in6653_1, in6653_2;
    wire c6653;
    assign in6653_1 = {s3614[0]};
    assign in6653_2 = {s3615[0]};
    Full_Adder FA_6653(s6653, c6653, in6653_1, in6653_2, s3613[0]);
    wire[0:0] s6654, in6654_1, in6654_2;
    wire c6654;
    assign in6654_1 = {s3617[0]};
    assign in6654_2 = {s3618[0]};
    Full_Adder FA_6654(s6654, c6654, in6654_1, in6654_2, s3616[0]);
    wire[0:0] s6655, in6655_1, in6655_2;
    wire c6655;
    assign in6655_1 = {s3620[0]};
    assign in6655_2 = {s3621[0]};
    Full_Adder FA_6655(s6655, c6655, in6655_1, in6655_2, s3619[0]);
    wire[0:0] s6656, in6656_1, in6656_2;
    wire c6656;
    assign in6656_1 = {s3623[0]};
    assign in6656_2 = {s3624[0]};
    Full_Adder FA_6656(s6656, c6656, in6656_1, in6656_2, s3622[0]);
    wire[0:0] s6657, in6657_1, in6657_2;
    wire c6657;
    assign in6657_1 = {s3626[0]};
    assign in6657_2 = {s3627[0]};
    Full_Adder FA_6657(s6657, c6657, in6657_1, in6657_2, s3625[0]);
    wire[0:0] s6658, in6658_1, in6658_2;
    wire c6658;
    assign in6658_1 = {s3629[0]};
    assign in6658_2 = {s3630[0]};
    Full_Adder FA_6658(s6658, c6658, in6658_1, in6658_2, s3628[0]);
    wire[0:0] s6659, in6659_1, in6659_2;
    wire c6659;
    assign in6659_1 = {s3632[0]};
    assign in6659_2 = {s3633[0]};
    Full_Adder FA_6659(s6659, c6659, in6659_1, in6659_2, s3631[0]);
    wire[0:0] s6660, in6660_1, in6660_2;
    wire c6660;
    assign in6660_1 = {s3635[0]};
    assign in6660_2 = {s3636[0]};
    Full_Adder FA_6660(s6660, c6660, in6660_1, in6660_2, s3634[0]);
    wire[0:0] s6661, in6661_1, in6661_2;
    wire c6661;
    assign in6661_1 = {s3638[0]};
    assign in6661_2 = {s3639[0]};
    Full_Adder FA_6661(s6661, c6661, in6661_1, in6661_2, s3637[0]);
    wire[0:0] s6662, in6662_1, in6662_2;
    wire c6662;
    assign in6662_1 = {s1278[0]};
    assign in6662_2 = {c3613};
    Full_Adder FA_6662(s6662, c6662, in6662_1, in6662_2, s1277[0]);
    wire[0:0] s6663, in6663_1, in6663_2;
    wire c6663;
    assign in6663_1 = {c3615};
    assign in6663_2 = {c3616};
    Full_Adder FA_6663(s6663, c6663, in6663_1, in6663_2, c3614);
    wire[0:0] s6664, in6664_1, in6664_2;
    wire c6664;
    assign in6664_1 = {c3618};
    assign in6664_2 = {c3619};
    Full_Adder FA_6664(s6664, c6664, in6664_1, in6664_2, c3617);
    wire[0:0] s6665, in6665_1, in6665_2;
    wire c6665;
    assign in6665_1 = {c3621};
    assign in6665_2 = {c3622};
    Full_Adder FA_6665(s6665, c6665, in6665_1, in6665_2, c3620);
    wire[0:0] s6666, in6666_1, in6666_2;
    wire c6666;
    assign in6666_1 = {c3624};
    assign in6666_2 = {c3625};
    Full_Adder FA_6666(s6666, c6666, in6666_1, in6666_2, c3623);
    wire[0:0] s6667, in6667_1, in6667_2;
    wire c6667;
    assign in6667_1 = {c3627};
    assign in6667_2 = {c3628};
    Full_Adder FA_6667(s6667, c6667, in6667_1, in6667_2, c3626);
    wire[0:0] s6668, in6668_1, in6668_2;
    wire c6668;
    assign in6668_1 = {c3630};
    assign in6668_2 = {c3631};
    Full_Adder FA_6668(s6668, c6668, in6668_1, in6668_2, c3629);
    wire[0:0] s6669, in6669_1, in6669_2;
    wire c6669;
    assign in6669_1 = {c3633};
    assign in6669_2 = {c3634};
    Full_Adder FA_6669(s6669, c6669, in6669_1, in6669_2, c3632);
    wire[0:0] s6670, in6670_1, in6670_2;
    wire c6670;
    assign in6670_1 = {c3636};
    assign in6670_2 = {c3637};
    Full_Adder FA_6670(s6670, c6670, in6670_1, in6670_2, c3635);
    wire[0:0] s6671, in6671_1, in6671_2;
    wire c6671;
    assign in6671_1 = {c3639};
    assign in6671_2 = {c3640};
    Full_Adder FA_6671(s6671, c6671, in6671_1, in6671_2, c3638);
    wire[0:0] s6672, in6672_1, in6672_2;
    wire c6672;
    assign in6672_1 = {s3642[0]};
    assign in6672_2 = {s3643[0]};
    Full_Adder FA_6672(s6672, c6672, in6672_1, in6672_2, s3641[0]);
    wire[0:0] s6673, in6673_1, in6673_2;
    wire c6673;
    assign in6673_1 = {s3645[0]};
    assign in6673_2 = {s3646[0]};
    Full_Adder FA_6673(s6673, c6673, in6673_1, in6673_2, s3644[0]);
    wire[0:0] s6674, in6674_1, in6674_2;
    wire c6674;
    assign in6674_1 = {s3648[0]};
    assign in6674_2 = {s3649[0]};
    Full_Adder FA_6674(s6674, c6674, in6674_1, in6674_2, s3647[0]);
    wire[0:0] s6675, in6675_1, in6675_2;
    wire c6675;
    assign in6675_1 = {s3651[0]};
    assign in6675_2 = {s3652[0]};
    Full_Adder FA_6675(s6675, c6675, in6675_1, in6675_2, s3650[0]);
    wire[0:0] s6676, in6676_1, in6676_2;
    wire c6676;
    assign in6676_1 = {s3654[0]};
    assign in6676_2 = {s3655[0]};
    Full_Adder FA_6676(s6676, c6676, in6676_1, in6676_2, s3653[0]);
    wire[0:0] s6677, in6677_1, in6677_2;
    wire c6677;
    assign in6677_1 = {s3657[0]};
    assign in6677_2 = {s3658[0]};
    Full_Adder FA_6677(s6677, c6677, in6677_1, in6677_2, s3656[0]);
    wire[0:0] s6678, in6678_1, in6678_2;
    wire c6678;
    assign in6678_1 = {s3660[0]};
    assign in6678_2 = {s3661[0]};
    Full_Adder FA_6678(s6678, c6678, in6678_1, in6678_2, s3659[0]);
    wire[0:0] s6679, in6679_1, in6679_2;
    wire c6679;
    assign in6679_1 = {s3663[0]};
    assign in6679_2 = {s3664[0]};
    Full_Adder FA_6679(s6679, c6679, in6679_1, in6679_2, s3662[0]);
    wire[0:0] s6680, in6680_1, in6680_2;
    wire c6680;
    assign in6680_1 = {s3666[0]};
    assign in6680_2 = {s3667[0]};
    Full_Adder FA_6680(s6680, c6680, in6680_1, in6680_2, s3665[0]);
    wire[0:0] s6681, in6681_1, in6681_2;
    wire c6681;
    assign in6681_1 = {s1310[0]};
    assign in6681_2 = {c3641};
    Full_Adder FA_6681(s6681, c6681, in6681_1, in6681_2, s1309[0]);
    wire[0:0] s6682, in6682_1, in6682_2;
    wire c6682;
    assign in6682_1 = {c3643};
    assign in6682_2 = {c3644};
    Full_Adder FA_6682(s6682, c6682, in6682_1, in6682_2, c3642);
    wire[0:0] s6683, in6683_1, in6683_2;
    wire c6683;
    assign in6683_1 = {c3646};
    assign in6683_2 = {c3647};
    Full_Adder FA_6683(s6683, c6683, in6683_1, in6683_2, c3645);
    wire[0:0] s6684, in6684_1, in6684_2;
    wire c6684;
    assign in6684_1 = {c3649};
    assign in6684_2 = {c3650};
    Full_Adder FA_6684(s6684, c6684, in6684_1, in6684_2, c3648);
    wire[0:0] s6685, in6685_1, in6685_2;
    wire c6685;
    assign in6685_1 = {c3652};
    assign in6685_2 = {c3653};
    Full_Adder FA_6685(s6685, c6685, in6685_1, in6685_2, c3651);
    wire[0:0] s6686, in6686_1, in6686_2;
    wire c6686;
    assign in6686_1 = {c3655};
    assign in6686_2 = {c3656};
    Full_Adder FA_6686(s6686, c6686, in6686_1, in6686_2, c3654);
    wire[0:0] s6687, in6687_1, in6687_2;
    wire c6687;
    assign in6687_1 = {c3658};
    assign in6687_2 = {c3659};
    Full_Adder FA_6687(s6687, c6687, in6687_1, in6687_2, c3657);
    wire[0:0] s6688, in6688_1, in6688_2;
    wire c6688;
    assign in6688_1 = {c3661};
    assign in6688_2 = {c3662};
    Full_Adder FA_6688(s6688, c6688, in6688_1, in6688_2, c3660);
    wire[0:0] s6689, in6689_1, in6689_2;
    wire c6689;
    assign in6689_1 = {c3664};
    assign in6689_2 = {c3665};
    Full_Adder FA_6689(s6689, c6689, in6689_1, in6689_2, c3663);
    wire[0:0] s6690, in6690_1, in6690_2;
    wire c6690;
    assign in6690_1 = {c3667};
    assign in6690_2 = {c3668};
    Full_Adder FA_6690(s6690, c6690, in6690_1, in6690_2, c3666);
    wire[0:0] s6691, in6691_1, in6691_2;
    wire c6691;
    assign in6691_1 = {s3670[0]};
    assign in6691_2 = {s3671[0]};
    Full_Adder FA_6691(s6691, c6691, in6691_1, in6691_2, s3669[0]);
    wire[0:0] s6692, in6692_1, in6692_2;
    wire c6692;
    assign in6692_1 = {s3673[0]};
    assign in6692_2 = {s3674[0]};
    Full_Adder FA_6692(s6692, c6692, in6692_1, in6692_2, s3672[0]);
    wire[0:0] s6693, in6693_1, in6693_2;
    wire c6693;
    assign in6693_1 = {s3676[0]};
    assign in6693_2 = {s3677[0]};
    Full_Adder FA_6693(s6693, c6693, in6693_1, in6693_2, s3675[0]);
    wire[0:0] s6694, in6694_1, in6694_2;
    wire c6694;
    assign in6694_1 = {s3679[0]};
    assign in6694_2 = {s3680[0]};
    Full_Adder FA_6694(s6694, c6694, in6694_1, in6694_2, s3678[0]);
    wire[0:0] s6695, in6695_1, in6695_2;
    wire c6695;
    assign in6695_1 = {s3682[0]};
    assign in6695_2 = {s3683[0]};
    Full_Adder FA_6695(s6695, c6695, in6695_1, in6695_2, s3681[0]);
    wire[0:0] s6696, in6696_1, in6696_2;
    wire c6696;
    assign in6696_1 = {s3685[0]};
    assign in6696_2 = {s3686[0]};
    Full_Adder FA_6696(s6696, c6696, in6696_1, in6696_2, s3684[0]);
    wire[0:0] s6697, in6697_1, in6697_2;
    wire c6697;
    assign in6697_1 = {s3688[0]};
    assign in6697_2 = {s3689[0]};
    Full_Adder FA_6697(s6697, c6697, in6697_1, in6697_2, s3687[0]);
    wire[0:0] s6698, in6698_1, in6698_2;
    wire c6698;
    assign in6698_1 = {s3691[0]};
    assign in6698_2 = {s3692[0]};
    Full_Adder FA_6698(s6698, c6698, in6698_1, in6698_2, s3690[0]);
    wire[0:0] s6699, in6699_1, in6699_2;
    wire c6699;
    assign in6699_1 = {s3694[0]};
    assign in6699_2 = {s3695[0]};
    Full_Adder FA_6699(s6699, c6699, in6699_1, in6699_2, s3693[0]);
    wire[0:0] s6700, in6700_1, in6700_2;
    wire c6700;
    assign in6700_1 = {s1341[0]};
    assign in6700_2 = {c3669};
    Full_Adder FA_6700(s6700, c6700, in6700_1, in6700_2, s1340[0]);
    wire[0:0] s6701, in6701_1, in6701_2;
    wire c6701;
    assign in6701_1 = {c3671};
    assign in6701_2 = {c3672};
    Full_Adder FA_6701(s6701, c6701, in6701_1, in6701_2, c3670);
    wire[0:0] s6702, in6702_1, in6702_2;
    wire c6702;
    assign in6702_1 = {c3674};
    assign in6702_2 = {c3675};
    Full_Adder FA_6702(s6702, c6702, in6702_1, in6702_2, c3673);
    wire[0:0] s6703, in6703_1, in6703_2;
    wire c6703;
    assign in6703_1 = {c3677};
    assign in6703_2 = {c3678};
    Full_Adder FA_6703(s6703, c6703, in6703_1, in6703_2, c3676);
    wire[0:0] s6704, in6704_1, in6704_2;
    wire c6704;
    assign in6704_1 = {c3680};
    assign in6704_2 = {c3681};
    Full_Adder FA_6704(s6704, c6704, in6704_1, in6704_2, c3679);
    wire[0:0] s6705, in6705_1, in6705_2;
    wire c6705;
    assign in6705_1 = {c3683};
    assign in6705_2 = {c3684};
    Full_Adder FA_6705(s6705, c6705, in6705_1, in6705_2, c3682);
    wire[0:0] s6706, in6706_1, in6706_2;
    wire c6706;
    assign in6706_1 = {c3686};
    assign in6706_2 = {c3687};
    Full_Adder FA_6706(s6706, c6706, in6706_1, in6706_2, c3685);
    wire[0:0] s6707, in6707_1, in6707_2;
    wire c6707;
    assign in6707_1 = {c3689};
    assign in6707_2 = {c3690};
    Full_Adder FA_6707(s6707, c6707, in6707_1, in6707_2, c3688);
    wire[0:0] s6708, in6708_1, in6708_2;
    wire c6708;
    assign in6708_1 = {c3692};
    assign in6708_2 = {c3693};
    Full_Adder FA_6708(s6708, c6708, in6708_1, in6708_2, c3691);
    wire[0:0] s6709, in6709_1, in6709_2;
    wire c6709;
    assign in6709_1 = {c3695};
    assign in6709_2 = {c3696};
    Full_Adder FA_6709(s6709, c6709, in6709_1, in6709_2, c3694);
    wire[0:0] s6710, in6710_1, in6710_2;
    wire c6710;
    assign in6710_1 = {s3698[0]};
    assign in6710_2 = {s3699[0]};
    Full_Adder FA_6710(s6710, c6710, in6710_1, in6710_2, s3697[0]);
    wire[0:0] s6711, in6711_1, in6711_2;
    wire c6711;
    assign in6711_1 = {s3701[0]};
    assign in6711_2 = {s3702[0]};
    Full_Adder FA_6711(s6711, c6711, in6711_1, in6711_2, s3700[0]);
    wire[0:0] s6712, in6712_1, in6712_2;
    wire c6712;
    assign in6712_1 = {s3704[0]};
    assign in6712_2 = {s3705[0]};
    Full_Adder FA_6712(s6712, c6712, in6712_1, in6712_2, s3703[0]);
    wire[0:0] s6713, in6713_1, in6713_2;
    wire c6713;
    assign in6713_1 = {s3707[0]};
    assign in6713_2 = {s3708[0]};
    Full_Adder FA_6713(s6713, c6713, in6713_1, in6713_2, s3706[0]);
    wire[0:0] s6714, in6714_1, in6714_2;
    wire c6714;
    assign in6714_1 = {s3710[0]};
    assign in6714_2 = {s3711[0]};
    Full_Adder FA_6714(s6714, c6714, in6714_1, in6714_2, s3709[0]);
    wire[0:0] s6715, in6715_1, in6715_2;
    wire c6715;
    assign in6715_1 = {s3713[0]};
    assign in6715_2 = {s3714[0]};
    Full_Adder FA_6715(s6715, c6715, in6715_1, in6715_2, s3712[0]);
    wire[0:0] s6716, in6716_1, in6716_2;
    wire c6716;
    assign in6716_1 = {s3716[0]};
    assign in6716_2 = {s3717[0]};
    Full_Adder FA_6716(s6716, c6716, in6716_1, in6716_2, s3715[0]);
    wire[0:0] s6717, in6717_1, in6717_2;
    wire c6717;
    assign in6717_1 = {s3719[0]};
    assign in6717_2 = {s3720[0]};
    Full_Adder FA_6717(s6717, c6717, in6717_1, in6717_2, s3718[0]);
    wire[0:0] s6718, in6718_1, in6718_2;
    wire c6718;
    assign in6718_1 = {s3722[0]};
    assign in6718_2 = {s3723[0]};
    Full_Adder FA_6718(s6718, c6718, in6718_1, in6718_2, s3721[0]);
    wire[0:0] s6719, in6719_1, in6719_2;
    wire c6719;
    assign in6719_1 = {s1371[0]};
    assign in6719_2 = {c3697};
    Full_Adder FA_6719(s6719, c6719, in6719_1, in6719_2, s1370[0]);
    wire[0:0] s6720, in6720_1, in6720_2;
    wire c6720;
    assign in6720_1 = {c3699};
    assign in6720_2 = {c3700};
    Full_Adder FA_6720(s6720, c6720, in6720_1, in6720_2, c3698);
    wire[0:0] s6721, in6721_1, in6721_2;
    wire c6721;
    assign in6721_1 = {c3702};
    assign in6721_2 = {c3703};
    Full_Adder FA_6721(s6721, c6721, in6721_1, in6721_2, c3701);
    wire[0:0] s6722, in6722_1, in6722_2;
    wire c6722;
    assign in6722_1 = {c3705};
    assign in6722_2 = {c3706};
    Full_Adder FA_6722(s6722, c6722, in6722_1, in6722_2, c3704);
    wire[0:0] s6723, in6723_1, in6723_2;
    wire c6723;
    assign in6723_1 = {c3708};
    assign in6723_2 = {c3709};
    Full_Adder FA_6723(s6723, c6723, in6723_1, in6723_2, c3707);
    wire[0:0] s6724, in6724_1, in6724_2;
    wire c6724;
    assign in6724_1 = {c3711};
    assign in6724_2 = {c3712};
    Full_Adder FA_6724(s6724, c6724, in6724_1, in6724_2, c3710);
    wire[0:0] s6725, in6725_1, in6725_2;
    wire c6725;
    assign in6725_1 = {c3714};
    assign in6725_2 = {c3715};
    Full_Adder FA_6725(s6725, c6725, in6725_1, in6725_2, c3713);
    wire[0:0] s6726, in6726_1, in6726_2;
    wire c6726;
    assign in6726_1 = {c3717};
    assign in6726_2 = {c3718};
    Full_Adder FA_6726(s6726, c6726, in6726_1, in6726_2, c3716);
    wire[0:0] s6727, in6727_1, in6727_2;
    wire c6727;
    assign in6727_1 = {c3720};
    assign in6727_2 = {c3721};
    Full_Adder FA_6727(s6727, c6727, in6727_1, in6727_2, c3719);
    wire[0:0] s6728, in6728_1, in6728_2;
    wire c6728;
    assign in6728_1 = {c3723};
    assign in6728_2 = {c3724};
    Full_Adder FA_6728(s6728, c6728, in6728_1, in6728_2, c3722);
    wire[0:0] s6729, in6729_1, in6729_2;
    wire c6729;
    assign in6729_1 = {s3726[0]};
    assign in6729_2 = {s3727[0]};
    Full_Adder FA_6729(s6729, c6729, in6729_1, in6729_2, s3725[0]);
    wire[0:0] s6730, in6730_1, in6730_2;
    wire c6730;
    assign in6730_1 = {s3729[0]};
    assign in6730_2 = {s3730[0]};
    Full_Adder FA_6730(s6730, c6730, in6730_1, in6730_2, s3728[0]);
    wire[0:0] s6731, in6731_1, in6731_2;
    wire c6731;
    assign in6731_1 = {s3732[0]};
    assign in6731_2 = {s3733[0]};
    Full_Adder FA_6731(s6731, c6731, in6731_1, in6731_2, s3731[0]);
    wire[0:0] s6732, in6732_1, in6732_2;
    wire c6732;
    assign in6732_1 = {s3735[0]};
    assign in6732_2 = {s3736[0]};
    Full_Adder FA_6732(s6732, c6732, in6732_1, in6732_2, s3734[0]);
    wire[0:0] s6733, in6733_1, in6733_2;
    wire c6733;
    assign in6733_1 = {s3738[0]};
    assign in6733_2 = {s3739[0]};
    Full_Adder FA_6733(s6733, c6733, in6733_1, in6733_2, s3737[0]);
    wire[0:0] s6734, in6734_1, in6734_2;
    wire c6734;
    assign in6734_1 = {s3741[0]};
    assign in6734_2 = {s3742[0]};
    Full_Adder FA_6734(s6734, c6734, in6734_1, in6734_2, s3740[0]);
    wire[0:0] s6735, in6735_1, in6735_2;
    wire c6735;
    assign in6735_1 = {s3744[0]};
    assign in6735_2 = {s3745[0]};
    Full_Adder FA_6735(s6735, c6735, in6735_1, in6735_2, s3743[0]);
    wire[0:0] s6736, in6736_1, in6736_2;
    wire c6736;
    assign in6736_1 = {s3747[0]};
    assign in6736_2 = {s3748[0]};
    Full_Adder FA_6736(s6736, c6736, in6736_1, in6736_2, s3746[0]);
    wire[0:0] s6737, in6737_1, in6737_2;
    wire c6737;
    assign in6737_1 = {s3750[0]};
    assign in6737_2 = {s3751[0]};
    Full_Adder FA_6737(s6737, c6737, in6737_1, in6737_2, s3749[0]);
    wire[0:0] s6738, in6738_1, in6738_2;
    wire c6738;
    assign in6738_1 = {s1400[0]};
    assign in6738_2 = {c3725};
    Full_Adder FA_6738(s6738, c6738, in6738_1, in6738_2, s1399[0]);
    wire[0:0] s6739, in6739_1, in6739_2;
    wire c6739;
    assign in6739_1 = {c3727};
    assign in6739_2 = {c3728};
    Full_Adder FA_6739(s6739, c6739, in6739_1, in6739_2, c3726);
    wire[0:0] s6740, in6740_1, in6740_2;
    wire c6740;
    assign in6740_1 = {c3730};
    assign in6740_2 = {c3731};
    Full_Adder FA_6740(s6740, c6740, in6740_1, in6740_2, c3729);
    wire[0:0] s6741, in6741_1, in6741_2;
    wire c6741;
    assign in6741_1 = {c3733};
    assign in6741_2 = {c3734};
    Full_Adder FA_6741(s6741, c6741, in6741_1, in6741_2, c3732);
    wire[0:0] s6742, in6742_1, in6742_2;
    wire c6742;
    assign in6742_1 = {c3736};
    assign in6742_2 = {c3737};
    Full_Adder FA_6742(s6742, c6742, in6742_1, in6742_2, c3735);
    wire[0:0] s6743, in6743_1, in6743_2;
    wire c6743;
    assign in6743_1 = {c3739};
    assign in6743_2 = {c3740};
    Full_Adder FA_6743(s6743, c6743, in6743_1, in6743_2, c3738);
    wire[0:0] s6744, in6744_1, in6744_2;
    wire c6744;
    assign in6744_1 = {c3742};
    assign in6744_2 = {c3743};
    Full_Adder FA_6744(s6744, c6744, in6744_1, in6744_2, c3741);
    wire[0:0] s6745, in6745_1, in6745_2;
    wire c6745;
    assign in6745_1 = {c3745};
    assign in6745_2 = {c3746};
    Full_Adder FA_6745(s6745, c6745, in6745_1, in6745_2, c3744);
    wire[0:0] s6746, in6746_1, in6746_2;
    wire c6746;
    assign in6746_1 = {c3748};
    assign in6746_2 = {c3749};
    Full_Adder FA_6746(s6746, c6746, in6746_1, in6746_2, c3747);
    wire[0:0] s6747, in6747_1, in6747_2;
    wire c6747;
    assign in6747_1 = {c3751};
    assign in6747_2 = {c3752};
    Full_Adder FA_6747(s6747, c6747, in6747_1, in6747_2, c3750);
    wire[0:0] s6748, in6748_1, in6748_2;
    wire c6748;
    assign in6748_1 = {s3754[0]};
    assign in6748_2 = {s3755[0]};
    Full_Adder FA_6748(s6748, c6748, in6748_1, in6748_2, s3753[0]);
    wire[0:0] s6749, in6749_1, in6749_2;
    wire c6749;
    assign in6749_1 = {s3757[0]};
    assign in6749_2 = {s3758[0]};
    Full_Adder FA_6749(s6749, c6749, in6749_1, in6749_2, s3756[0]);
    wire[0:0] s6750, in6750_1, in6750_2;
    wire c6750;
    assign in6750_1 = {s3760[0]};
    assign in6750_2 = {s3761[0]};
    Full_Adder FA_6750(s6750, c6750, in6750_1, in6750_2, s3759[0]);
    wire[0:0] s6751, in6751_1, in6751_2;
    wire c6751;
    assign in6751_1 = {s3763[0]};
    assign in6751_2 = {s3764[0]};
    Full_Adder FA_6751(s6751, c6751, in6751_1, in6751_2, s3762[0]);
    wire[0:0] s6752, in6752_1, in6752_2;
    wire c6752;
    assign in6752_1 = {s3766[0]};
    assign in6752_2 = {s3767[0]};
    Full_Adder FA_6752(s6752, c6752, in6752_1, in6752_2, s3765[0]);
    wire[0:0] s6753, in6753_1, in6753_2;
    wire c6753;
    assign in6753_1 = {s3769[0]};
    assign in6753_2 = {s3770[0]};
    Full_Adder FA_6753(s6753, c6753, in6753_1, in6753_2, s3768[0]);
    wire[0:0] s6754, in6754_1, in6754_2;
    wire c6754;
    assign in6754_1 = {s3772[0]};
    assign in6754_2 = {s3773[0]};
    Full_Adder FA_6754(s6754, c6754, in6754_1, in6754_2, s3771[0]);
    wire[0:0] s6755, in6755_1, in6755_2;
    wire c6755;
    assign in6755_1 = {s3775[0]};
    assign in6755_2 = {s3776[0]};
    Full_Adder FA_6755(s6755, c6755, in6755_1, in6755_2, s3774[0]);
    wire[0:0] s6756, in6756_1, in6756_2;
    wire c6756;
    assign in6756_1 = {s3778[0]};
    assign in6756_2 = {s3779[0]};
    Full_Adder FA_6756(s6756, c6756, in6756_1, in6756_2, s3777[0]);
    wire[0:0] s6757, in6757_1, in6757_2;
    wire c6757;
    assign in6757_1 = {s1428[0]};
    assign in6757_2 = {c3753};
    Full_Adder FA_6757(s6757, c6757, in6757_1, in6757_2, s1427[0]);
    wire[0:0] s6758, in6758_1, in6758_2;
    wire c6758;
    assign in6758_1 = {c3755};
    assign in6758_2 = {c3756};
    Full_Adder FA_6758(s6758, c6758, in6758_1, in6758_2, c3754);
    wire[0:0] s6759, in6759_1, in6759_2;
    wire c6759;
    assign in6759_1 = {c3758};
    assign in6759_2 = {c3759};
    Full_Adder FA_6759(s6759, c6759, in6759_1, in6759_2, c3757);
    wire[0:0] s6760, in6760_1, in6760_2;
    wire c6760;
    assign in6760_1 = {c3761};
    assign in6760_2 = {c3762};
    Full_Adder FA_6760(s6760, c6760, in6760_1, in6760_2, c3760);
    wire[0:0] s6761, in6761_1, in6761_2;
    wire c6761;
    assign in6761_1 = {c3764};
    assign in6761_2 = {c3765};
    Full_Adder FA_6761(s6761, c6761, in6761_1, in6761_2, c3763);
    wire[0:0] s6762, in6762_1, in6762_2;
    wire c6762;
    assign in6762_1 = {c3767};
    assign in6762_2 = {c3768};
    Full_Adder FA_6762(s6762, c6762, in6762_1, in6762_2, c3766);
    wire[0:0] s6763, in6763_1, in6763_2;
    wire c6763;
    assign in6763_1 = {c3770};
    assign in6763_2 = {c3771};
    Full_Adder FA_6763(s6763, c6763, in6763_1, in6763_2, c3769);
    wire[0:0] s6764, in6764_1, in6764_2;
    wire c6764;
    assign in6764_1 = {c3773};
    assign in6764_2 = {c3774};
    Full_Adder FA_6764(s6764, c6764, in6764_1, in6764_2, c3772);
    wire[0:0] s6765, in6765_1, in6765_2;
    wire c6765;
    assign in6765_1 = {c3776};
    assign in6765_2 = {c3777};
    Full_Adder FA_6765(s6765, c6765, in6765_1, in6765_2, c3775);
    wire[0:0] s6766, in6766_1, in6766_2;
    wire c6766;
    assign in6766_1 = {c3779};
    assign in6766_2 = {c3780};
    Full_Adder FA_6766(s6766, c6766, in6766_1, in6766_2, c3778);
    wire[0:0] s6767, in6767_1, in6767_2;
    wire c6767;
    assign in6767_1 = {s3782[0]};
    assign in6767_2 = {s3783[0]};
    Full_Adder FA_6767(s6767, c6767, in6767_1, in6767_2, s3781[0]);
    wire[0:0] s6768, in6768_1, in6768_2;
    wire c6768;
    assign in6768_1 = {s3785[0]};
    assign in6768_2 = {s3786[0]};
    Full_Adder FA_6768(s6768, c6768, in6768_1, in6768_2, s3784[0]);
    wire[0:0] s6769, in6769_1, in6769_2;
    wire c6769;
    assign in6769_1 = {s3788[0]};
    assign in6769_2 = {s3789[0]};
    Full_Adder FA_6769(s6769, c6769, in6769_1, in6769_2, s3787[0]);
    wire[0:0] s6770, in6770_1, in6770_2;
    wire c6770;
    assign in6770_1 = {s3791[0]};
    assign in6770_2 = {s3792[0]};
    Full_Adder FA_6770(s6770, c6770, in6770_1, in6770_2, s3790[0]);
    wire[0:0] s6771, in6771_1, in6771_2;
    wire c6771;
    assign in6771_1 = {s3794[0]};
    assign in6771_2 = {s3795[0]};
    Full_Adder FA_6771(s6771, c6771, in6771_1, in6771_2, s3793[0]);
    wire[0:0] s6772, in6772_1, in6772_2;
    wire c6772;
    assign in6772_1 = {s3797[0]};
    assign in6772_2 = {s3798[0]};
    Full_Adder FA_6772(s6772, c6772, in6772_1, in6772_2, s3796[0]);
    wire[0:0] s6773, in6773_1, in6773_2;
    wire c6773;
    assign in6773_1 = {s3800[0]};
    assign in6773_2 = {s3801[0]};
    Full_Adder FA_6773(s6773, c6773, in6773_1, in6773_2, s3799[0]);
    wire[0:0] s6774, in6774_1, in6774_2;
    wire c6774;
    assign in6774_1 = {s3803[0]};
    assign in6774_2 = {s3804[0]};
    Full_Adder FA_6774(s6774, c6774, in6774_1, in6774_2, s3802[0]);
    wire[0:0] s6775, in6775_1, in6775_2;
    wire c6775;
    assign in6775_1 = {s3806[0]};
    assign in6775_2 = {s3807[0]};
    Full_Adder FA_6775(s6775, c6775, in6775_1, in6775_2, s3805[0]);
    wire[0:0] s6776, in6776_1, in6776_2;
    wire c6776;
    assign in6776_1 = {s1455[0]};
    assign in6776_2 = {c3781};
    Full_Adder FA_6776(s6776, c6776, in6776_1, in6776_2, s1454[0]);
    wire[0:0] s6777, in6777_1, in6777_2;
    wire c6777;
    assign in6777_1 = {c3783};
    assign in6777_2 = {c3784};
    Full_Adder FA_6777(s6777, c6777, in6777_1, in6777_2, c3782);
    wire[0:0] s6778, in6778_1, in6778_2;
    wire c6778;
    assign in6778_1 = {c3786};
    assign in6778_2 = {c3787};
    Full_Adder FA_6778(s6778, c6778, in6778_1, in6778_2, c3785);
    wire[0:0] s6779, in6779_1, in6779_2;
    wire c6779;
    assign in6779_1 = {c3789};
    assign in6779_2 = {c3790};
    Full_Adder FA_6779(s6779, c6779, in6779_1, in6779_2, c3788);
    wire[0:0] s6780, in6780_1, in6780_2;
    wire c6780;
    assign in6780_1 = {c3792};
    assign in6780_2 = {c3793};
    Full_Adder FA_6780(s6780, c6780, in6780_1, in6780_2, c3791);
    wire[0:0] s6781, in6781_1, in6781_2;
    wire c6781;
    assign in6781_1 = {c3795};
    assign in6781_2 = {c3796};
    Full_Adder FA_6781(s6781, c6781, in6781_1, in6781_2, c3794);
    wire[0:0] s6782, in6782_1, in6782_2;
    wire c6782;
    assign in6782_1 = {c3798};
    assign in6782_2 = {c3799};
    Full_Adder FA_6782(s6782, c6782, in6782_1, in6782_2, c3797);
    wire[0:0] s6783, in6783_1, in6783_2;
    wire c6783;
    assign in6783_1 = {c3801};
    assign in6783_2 = {c3802};
    Full_Adder FA_6783(s6783, c6783, in6783_1, in6783_2, c3800);
    wire[0:0] s6784, in6784_1, in6784_2;
    wire c6784;
    assign in6784_1 = {c3804};
    assign in6784_2 = {c3805};
    Full_Adder FA_6784(s6784, c6784, in6784_1, in6784_2, c3803);
    wire[0:0] s6785, in6785_1, in6785_2;
    wire c6785;
    assign in6785_1 = {c3807};
    assign in6785_2 = {c3808};
    Full_Adder FA_6785(s6785, c6785, in6785_1, in6785_2, c3806);
    wire[0:0] s6786, in6786_1, in6786_2;
    wire c6786;
    assign in6786_1 = {s3810[0]};
    assign in6786_2 = {s3811[0]};
    Full_Adder FA_6786(s6786, c6786, in6786_1, in6786_2, s3809[0]);
    wire[0:0] s6787, in6787_1, in6787_2;
    wire c6787;
    assign in6787_1 = {s3813[0]};
    assign in6787_2 = {s3814[0]};
    Full_Adder FA_6787(s6787, c6787, in6787_1, in6787_2, s3812[0]);
    wire[0:0] s6788, in6788_1, in6788_2;
    wire c6788;
    assign in6788_1 = {s3816[0]};
    assign in6788_2 = {s3817[0]};
    Full_Adder FA_6788(s6788, c6788, in6788_1, in6788_2, s3815[0]);
    wire[0:0] s6789, in6789_1, in6789_2;
    wire c6789;
    assign in6789_1 = {s3819[0]};
    assign in6789_2 = {s3820[0]};
    Full_Adder FA_6789(s6789, c6789, in6789_1, in6789_2, s3818[0]);
    wire[0:0] s6790, in6790_1, in6790_2;
    wire c6790;
    assign in6790_1 = {s3822[0]};
    assign in6790_2 = {s3823[0]};
    Full_Adder FA_6790(s6790, c6790, in6790_1, in6790_2, s3821[0]);
    wire[0:0] s6791, in6791_1, in6791_2;
    wire c6791;
    assign in6791_1 = {s3825[0]};
    assign in6791_2 = {s3826[0]};
    Full_Adder FA_6791(s6791, c6791, in6791_1, in6791_2, s3824[0]);
    wire[0:0] s6792, in6792_1, in6792_2;
    wire c6792;
    assign in6792_1 = {s3828[0]};
    assign in6792_2 = {s3829[0]};
    Full_Adder FA_6792(s6792, c6792, in6792_1, in6792_2, s3827[0]);
    wire[0:0] s6793, in6793_1, in6793_2;
    wire c6793;
    assign in6793_1 = {s3831[0]};
    assign in6793_2 = {s3832[0]};
    Full_Adder FA_6793(s6793, c6793, in6793_1, in6793_2, s3830[0]);
    wire[0:0] s6794, in6794_1, in6794_2;
    wire c6794;
    assign in6794_1 = {s3834[0]};
    assign in6794_2 = {s3835[0]};
    Full_Adder FA_6794(s6794, c6794, in6794_1, in6794_2, s3833[0]);
    wire[0:0] s6795, in6795_1, in6795_2;
    wire c6795;
    assign in6795_1 = {s1481[0]};
    assign in6795_2 = {c3809};
    Full_Adder FA_6795(s6795, c6795, in6795_1, in6795_2, s1480[0]);
    wire[0:0] s6796, in6796_1, in6796_2;
    wire c6796;
    assign in6796_1 = {c3811};
    assign in6796_2 = {c3812};
    Full_Adder FA_6796(s6796, c6796, in6796_1, in6796_2, c3810);
    wire[0:0] s6797, in6797_1, in6797_2;
    wire c6797;
    assign in6797_1 = {c3814};
    assign in6797_2 = {c3815};
    Full_Adder FA_6797(s6797, c6797, in6797_1, in6797_2, c3813);
    wire[0:0] s6798, in6798_1, in6798_2;
    wire c6798;
    assign in6798_1 = {c3817};
    assign in6798_2 = {c3818};
    Full_Adder FA_6798(s6798, c6798, in6798_1, in6798_2, c3816);
    wire[0:0] s6799, in6799_1, in6799_2;
    wire c6799;
    assign in6799_1 = {c3820};
    assign in6799_2 = {c3821};
    Full_Adder FA_6799(s6799, c6799, in6799_1, in6799_2, c3819);
    wire[0:0] s6800, in6800_1, in6800_2;
    wire c6800;
    assign in6800_1 = {c3823};
    assign in6800_2 = {c3824};
    Full_Adder FA_6800(s6800, c6800, in6800_1, in6800_2, c3822);
    wire[0:0] s6801, in6801_1, in6801_2;
    wire c6801;
    assign in6801_1 = {c3826};
    assign in6801_2 = {c3827};
    Full_Adder FA_6801(s6801, c6801, in6801_1, in6801_2, c3825);
    wire[0:0] s6802, in6802_1, in6802_2;
    wire c6802;
    assign in6802_1 = {c3829};
    assign in6802_2 = {c3830};
    Full_Adder FA_6802(s6802, c6802, in6802_1, in6802_2, c3828);
    wire[0:0] s6803, in6803_1, in6803_2;
    wire c6803;
    assign in6803_1 = {c3832};
    assign in6803_2 = {c3833};
    Full_Adder FA_6803(s6803, c6803, in6803_1, in6803_2, c3831);
    wire[0:0] s6804, in6804_1, in6804_2;
    wire c6804;
    assign in6804_1 = {c3835};
    assign in6804_2 = {c3836};
    Full_Adder FA_6804(s6804, c6804, in6804_1, in6804_2, c3834);
    wire[0:0] s6805, in6805_1, in6805_2;
    wire c6805;
    assign in6805_1 = {s3838[0]};
    assign in6805_2 = {s3839[0]};
    Full_Adder FA_6805(s6805, c6805, in6805_1, in6805_2, s3837[0]);
    wire[0:0] s6806, in6806_1, in6806_2;
    wire c6806;
    assign in6806_1 = {s3841[0]};
    assign in6806_2 = {s3842[0]};
    Full_Adder FA_6806(s6806, c6806, in6806_1, in6806_2, s3840[0]);
    wire[0:0] s6807, in6807_1, in6807_2;
    wire c6807;
    assign in6807_1 = {s3844[0]};
    assign in6807_2 = {s3845[0]};
    Full_Adder FA_6807(s6807, c6807, in6807_1, in6807_2, s3843[0]);
    wire[0:0] s6808, in6808_1, in6808_2;
    wire c6808;
    assign in6808_1 = {s3847[0]};
    assign in6808_2 = {s3848[0]};
    Full_Adder FA_6808(s6808, c6808, in6808_1, in6808_2, s3846[0]);
    wire[0:0] s6809, in6809_1, in6809_2;
    wire c6809;
    assign in6809_1 = {s3850[0]};
    assign in6809_2 = {s3851[0]};
    Full_Adder FA_6809(s6809, c6809, in6809_1, in6809_2, s3849[0]);
    wire[0:0] s6810, in6810_1, in6810_2;
    wire c6810;
    assign in6810_1 = {s3853[0]};
    assign in6810_2 = {s3854[0]};
    Full_Adder FA_6810(s6810, c6810, in6810_1, in6810_2, s3852[0]);
    wire[0:0] s6811, in6811_1, in6811_2;
    wire c6811;
    assign in6811_1 = {s3856[0]};
    assign in6811_2 = {s3857[0]};
    Full_Adder FA_6811(s6811, c6811, in6811_1, in6811_2, s3855[0]);
    wire[0:0] s6812, in6812_1, in6812_2;
    wire c6812;
    assign in6812_1 = {s3859[0]};
    assign in6812_2 = {s3860[0]};
    Full_Adder FA_6812(s6812, c6812, in6812_1, in6812_2, s3858[0]);
    wire[0:0] s6813, in6813_1, in6813_2;
    wire c6813;
    assign in6813_1 = {s3862[0]};
    assign in6813_2 = {s3863[0]};
    Full_Adder FA_6813(s6813, c6813, in6813_1, in6813_2, s3861[0]);
    wire[0:0] s6814, in6814_1, in6814_2;
    wire c6814;
    assign in6814_1 = {s1506[0]};
    assign in6814_2 = {c3837};
    Full_Adder FA_6814(s6814, c6814, in6814_1, in6814_2, s1505[0]);
    wire[0:0] s6815, in6815_1, in6815_2;
    wire c6815;
    assign in6815_1 = {c3839};
    assign in6815_2 = {c3840};
    Full_Adder FA_6815(s6815, c6815, in6815_1, in6815_2, c3838);
    wire[0:0] s6816, in6816_1, in6816_2;
    wire c6816;
    assign in6816_1 = {c3842};
    assign in6816_2 = {c3843};
    Full_Adder FA_6816(s6816, c6816, in6816_1, in6816_2, c3841);
    wire[0:0] s6817, in6817_1, in6817_2;
    wire c6817;
    assign in6817_1 = {c3845};
    assign in6817_2 = {c3846};
    Full_Adder FA_6817(s6817, c6817, in6817_1, in6817_2, c3844);
    wire[0:0] s6818, in6818_1, in6818_2;
    wire c6818;
    assign in6818_1 = {c3848};
    assign in6818_2 = {c3849};
    Full_Adder FA_6818(s6818, c6818, in6818_1, in6818_2, c3847);
    wire[0:0] s6819, in6819_1, in6819_2;
    wire c6819;
    assign in6819_1 = {c3851};
    assign in6819_2 = {c3852};
    Full_Adder FA_6819(s6819, c6819, in6819_1, in6819_2, c3850);
    wire[0:0] s6820, in6820_1, in6820_2;
    wire c6820;
    assign in6820_1 = {c3854};
    assign in6820_2 = {c3855};
    Full_Adder FA_6820(s6820, c6820, in6820_1, in6820_2, c3853);
    wire[0:0] s6821, in6821_1, in6821_2;
    wire c6821;
    assign in6821_1 = {c3857};
    assign in6821_2 = {c3858};
    Full_Adder FA_6821(s6821, c6821, in6821_1, in6821_2, c3856);
    wire[0:0] s6822, in6822_1, in6822_2;
    wire c6822;
    assign in6822_1 = {c3860};
    assign in6822_2 = {c3861};
    Full_Adder FA_6822(s6822, c6822, in6822_1, in6822_2, c3859);
    wire[0:0] s6823, in6823_1, in6823_2;
    wire c6823;
    assign in6823_1 = {c3863};
    assign in6823_2 = {c3864};
    Full_Adder FA_6823(s6823, c6823, in6823_1, in6823_2, c3862);
    wire[0:0] s6824, in6824_1, in6824_2;
    wire c6824;
    assign in6824_1 = {s3866[0]};
    assign in6824_2 = {s3867[0]};
    Full_Adder FA_6824(s6824, c6824, in6824_1, in6824_2, s3865[0]);
    wire[0:0] s6825, in6825_1, in6825_2;
    wire c6825;
    assign in6825_1 = {s3869[0]};
    assign in6825_2 = {s3870[0]};
    Full_Adder FA_6825(s6825, c6825, in6825_1, in6825_2, s3868[0]);
    wire[0:0] s6826, in6826_1, in6826_2;
    wire c6826;
    assign in6826_1 = {s3872[0]};
    assign in6826_2 = {s3873[0]};
    Full_Adder FA_6826(s6826, c6826, in6826_1, in6826_2, s3871[0]);
    wire[0:0] s6827, in6827_1, in6827_2;
    wire c6827;
    assign in6827_1 = {s3875[0]};
    assign in6827_2 = {s3876[0]};
    Full_Adder FA_6827(s6827, c6827, in6827_1, in6827_2, s3874[0]);
    wire[0:0] s6828, in6828_1, in6828_2;
    wire c6828;
    assign in6828_1 = {s3878[0]};
    assign in6828_2 = {s3879[0]};
    Full_Adder FA_6828(s6828, c6828, in6828_1, in6828_2, s3877[0]);
    wire[0:0] s6829, in6829_1, in6829_2;
    wire c6829;
    assign in6829_1 = {s3881[0]};
    assign in6829_2 = {s3882[0]};
    Full_Adder FA_6829(s6829, c6829, in6829_1, in6829_2, s3880[0]);
    wire[0:0] s6830, in6830_1, in6830_2;
    wire c6830;
    assign in6830_1 = {s3884[0]};
    assign in6830_2 = {s3885[0]};
    Full_Adder FA_6830(s6830, c6830, in6830_1, in6830_2, s3883[0]);
    wire[0:0] s6831, in6831_1, in6831_2;
    wire c6831;
    assign in6831_1 = {s3887[0]};
    assign in6831_2 = {s3888[0]};
    Full_Adder FA_6831(s6831, c6831, in6831_1, in6831_2, s3886[0]);
    wire[0:0] s6832, in6832_1, in6832_2;
    wire c6832;
    assign in6832_1 = {s3890[0]};
    assign in6832_2 = {s3891[0]};
    Full_Adder FA_6832(s6832, c6832, in6832_1, in6832_2, s3889[0]);
    wire[0:0] s6833, in6833_1, in6833_2;
    wire c6833;
    assign in6833_1 = {s1530[0]};
    assign in6833_2 = {c3865};
    Full_Adder FA_6833(s6833, c6833, in6833_1, in6833_2, s1529[0]);
    wire[0:0] s6834, in6834_1, in6834_2;
    wire c6834;
    assign in6834_1 = {c3867};
    assign in6834_2 = {c3868};
    Full_Adder FA_6834(s6834, c6834, in6834_1, in6834_2, c3866);
    wire[0:0] s6835, in6835_1, in6835_2;
    wire c6835;
    assign in6835_1 = {c3870};
    assign in6835_2 = {c3871};
    Full_Adder FA_6835(s6835, c6835, in6835_1, in6835_2, c3869);
    wire[0:0] s6836, in6836_1, in6836_2;
    wire c6836;
    assign in6836_1 = {c3873};
    assign in6836_2 = {c3874};
    Full_Adder FA_6836(s6836, c6836, in6836_1, in6836_2, c3872);
    wire[0:0] s6837, in6837_1, in6837_2;
    wire c6837;
    assign in6837_1 = {c3876};
    assign in6837_2 = {c3877};
    Full_Adder FA_6837(s6837, c6837, in6837_1, in6837_2, c3875);
    wire[0:0] s6838, in6838_1, in6838_2;
    wire c6838;
    assign in6838_1 = {c3879};
    assign in6838_2 = {c3880};
    Full_Adder FA_6838(s6838, c6838, in6838_1, in6838_2, c3878);
    wire[0:0] s6839, in6839_1, in6839_2;
    wire c6839;
    assign in6839_1 = {c3882};
    assign in6839_2 = {c3883};
    Full_Adder FA_6839(s6839, c6839, in6839_1, in6839_2, c3881);
    wire[0:0] s6840, in6840_1, in6840_2;
    wire c6840;
    assign in6840_1 = {c3885};
    assign in6840_2 = {c3886};
    Full_Adder FA_6840(s6840, c6840, in6840_1, in6840_2, c3884);
    wire[0:0] s6841, in6841_1, in6841_2;
    wire c6841;
    assign in6841_1 = {c3888};
    assign in6841_2 = {c3889};
    Full_Adder FA_6841(s6841, c6841, in6841_1, in6841_2, c3887);
    wire[0:0] s6842, in6842_1, in6842_2;
    wire c6842;
    assign in6842_1 = {c3891};
    assign in6842_2 = {c3892};
    Full_Adder FA_6842(s6842, c6842, in6842_1, in6842_2, c3890);
    wire[0:0] s6843, in6843_1, in6843_2;
    wire c6843;
    assign in6843_1 = {s3894[0]};
    assign in6843_2 = {s3895[0]};
    Full_Adder FA_6843(s6843, c6843, in6843_1, in6843_2, s3893[0]);
    wire[0:0] s6844, in6844_1, in6844_2;
    wire c6844;
    assign in6844_1 = {s3897[0]};
    assign in6844_2 = {s3898[0]};
    Full_Adder FA_6844(s6844, c6844, in6844_1, in6844_2, s3896[0]);
    wire[0:0] s6845, in6845_1, in6845_2;
    wire c6845;
    assign in6845_1 = {s3900[0]};
    assign in6845_2 = {s3901[0]};
    Full_Adder FA_6845(s6845, c6845, in6845_1, in6845_2, s3899[0]);
    wire[0:0] s6846, in6846_1, in6846_2;
    wire c6846;
    assign in6846_1 = {s3903[0]};
    assign in6846_2 = {s3904[0]};
    Full_Adder FA_6846(s6846, c6846, in6846_1, in6846_2, s3902[0]);
    wire[0:0] s6847, in6847_1, in6847_2;
    wire c6847;
    assign in6847_1 = {s3906[0]};
    assign in6847_2 = {s3907[0]};
    Full_Adder FA_6847(s6847, c6847, in6847_1, in6847_2, s3905[0]);
    wire[0:0] s6848, in6848_1, in6848_2;
    wire c6848;
    assign in6848_1 = {s3909[0]};
    assign in6848_2 = {s3910[0]};
    Full_Adder FA_6848(s6848, c6848, in6848_1, in6848_2, s3908[0]);
    wire[0:0] s6849, in6849_1, in6849_2;
    wire c6849;
    assign in6849_1 = {s3912[0]};
    assign in6849_2 = {s3913[0]};
    Full_Adder FA_6849(s6849, c6849, in6849_1, in6849_2, s3911[0]);
    wire[0:0] s6850, in6850_1, in6850_2;
    wire c6850;
    assign in6850_1 = {s3915[0]};
    assign in6850_2 = {s3916[0]};
    Full_Adder FA_6850(s6850, c6850, in6850_1, in6850_2, s3914[0]);
    wire[0:0] s6851, in6851_1, in6851_2;
    wire c6851;
    assign in6851_1 = {s3918[0]};
    assign in6851_2 = {s3919[0]};
    Full_Adder FA_6851(s6851, c6851, in6851_1, in6851_2, s3917[0]);
    wire[0:0] s6852, in6852_1, in6852_2;
    wire c6852;
    assign in6852_1 = {s1553[0]};
    assign in6852_2 = {c3893};
    Full_Adder FA_6852(s6852, c6852, in6852_1, in6852_2, s1552[0]);
    wire[0:0] s6853, in6853_1, in6853_2;
    wire c6853;
    assign in6853_1 = {c3895};
    assign in6853_2 = {c3896};
    Full_Adder FA_6853(s6853, c6853, in6853_1, in6853_2, c3894);
    wire[0:0] s6854, in6854_1, in6854_2;
    wire c6854;
    assign in6854_1 = {c3898};
    assign in6854_2 = {c3899};
    Full_Adder FA_6854(s6854, c6854, in6854_1, in6854_2, c3897);
    wire[0:0] s6855, in6855_1, in6855_2;
    wire c6855;
    assign in6855_1 = {c3901};
    assign in6855_2 = {c3902};
    Full_Adder FA_6855(s6855, c6855, in6855_1, in6855_2, c3900);
    wire[0:0] s6856, in6856_1, in6856_2;
    wire c6856;
    assign in6856_1 = {c3904};
    assign in6856_2 = {c3905};
    Full_Adder FA_6856(s6856, c6856, in6856_1, in6856_2, c3903);
    wire[0:0] s6857, in6857_1, in6857_2;
    wire c6857;
    assign in6857_1 = {c3907};
    assign in6857_2 = {c3908};
    Full_Adder FA_6857(s6857, c6857, in6857_1, in6857_2, c3906);
    wire[0:0] s6858, in6858_1, in6858_2;
    wire c6858;
    assign in6858_1 = {c3910};
    assign in6858_2 = {c3911};
    Full_Adder FA_6858(s6858, c6858, in6858_1, in6858_2, c3909);
    wire[0:0] s6859, in6859_1, in6859_2;
    wire c6859;
    assign in6859_1 = {c3913};
    assign in6859_2 = {c3914};
    Full_Adder FA_6859(s6859, c6859, in6859_1, in6859_2, c3912);
    wire[0:0] s6860, in6860_1, in6860_2;
    wire c6860;
    assign in6860_1 = {c3916};
    assign in6860_2 = {c3917};
    Full_Adder FA_6860(s6860, c6860, in6860_1, in6860_2, c3915);
    wire[0:0] s6861, in6861_1, in6861_2;
    wire c6861;
    assign in6861_1 = {c3919};
    assign in6861_2 = {c3920};
    Full_Adder FA_6861(s6861, c6861, in6861_1, in6861_2, c3918);
    wire[0:0] s6862, in6862_1, in6862_2;
    wire c6862;
    assign in6862_1 = {s3922[0]};
    assign in6862_2 = {s3923[0]};
    Full_Adder FA_6862(s6862, c6862, in6862_1, in6862_2, s3921[0]);
    wire[0:0] s6863, in6863_1, in6863_2;
    wire c6863;
    assign in6863_1 = {s3925[0]};
    assign in6863_2 = {s3926[0]};
    Full_Adder FA_6863(s6863, c6863, in6863_1, in6863_2, s3924[0]);
    wire[0:0] s6864, in6864_1, in6864_2;
    wire c6864;
    assign in6864_1 = {s3928[0]};
    assign in6864_2 = {s3929[0]};
    Full_Adder FA_6864(s6864, c6864, in6864_1, in6864_2, s3927[0]);
    wire[0:0] s6865, in6865_1, in6865_2;
    wire c6865;
    assign in6865_1 = {s3931[0]};
    assign in6865_2 = {s3932[0]};
    Full_Adder FA_6865(s6865, c6865, in6865_1, in6865_2, s3930[0]);
    wire[0:0] s6866, in6866_1, in6866_2;
    wire c6866;
    assign in6866_1 = {s3934[0]};
    assign in6866_2 = {s3935[0]};
    Full_Adder FA_6866(s6866, c6866, in6866_1, in6866_2, s3933[0]);
    wire[0:0] s6867, in6867_1, in6867_2;
    wire c6867;
    assign in6867_1 = {s3937[0]};
    assign in6867_2 = {s3938[0]};
    Full_Adder FA_6867(s6867, c6867, in6867_1, in6867_2, s3936[0]);
    wire[0:0] s6868, in6868_1, in6868_2;
    wire c6868;
    assign in6868_1 = {s3940[0]};
    assign in6868_2 = {s3941[0]};
    Full_Adder FA_6868(s6868, c6868, in6868_1, in6868_2, s3939[0]);
    wire[0:0] s6869, in6869_1, in6869_2;
    wire c6869;
    assign in6869_1 = {s3943[0]};
    assign in6869_2 = {s3944[0]};
    Full_Adder FA_6869(s6869, c6869, in6869_1, in6869_2, s3942[0]);
    wire[0:0] s6870, in6870_1, in6870_2;
    wire c6870;
    assign in6870_1 = {s3946[0]};
    assign in6870_2 = {s3947[0]};
    Full_Adder FA_6870(s6870, c6870, in6870_1, in6870_2, s3945[0]);
    wire[0:0] s6871, in6871_1, in6871_2;
    wire c6871;
    assign in6871_1 = {s1575[0]};
    assign in6871_2 = {c3921};
    Full_Adder FA_6871(s6871, c6871, in6871_1, in6871_2, s1574[0]);
    wire[0:0] s6872, in6872_1, in6872_2;
    wire c6872;
    assign in6872_1 = {c3923};
    assign in6872_2 = {c3924};
    Full_Adder FA_6872(s6872, c6872, in6872_1, in6872_2, c3922);
    wire[0:0] s6873, in6873_1, in6873_2;
    wire c6873;
    assign in6873_1 = {c3926};
    assign in6873_2 = {c3927};
    Full_Adder FA_6873(s6873, c6873, in6873_1, in6873_2, c3925);
    wire[0:0] s6874, in6874_1, in6874_2;
    wire c6874;
    assign in6874_1 = {c3929};
    assign in6874_2 = {c3930};
    Full_Adder FA_6874(s6874, c6874, in6874_1, in6874_2, c3928);
    wire[0:0] s6875, in6875_1, in6875_2;
    wire c6875;
    assign in6875_1 = {c3932};
    assign in6875_2 = {c3933};
    Full_Adder FA_6875(s6875, c6875, in6875_1, in6875_2, c3931);
    wire[0:0] s6876, in6876_1, in6876_2;
    wire c6876;
    assign in6876_1 = {c3935};
    assign in6876_2 = {c3936};
    Full_Adder FA_6876(s6876, c6876, in6876_1, in6876_2, c3934);
    wire[0:0] s6877, in6877_1, in6877_2;
    wire c6877;
    assign in6877_1 = {c3938};
    assign in6877_2 = {c3939};
    Full_Adder FA_6877(s6877, c6877, in6877_1, in6877_2, c3937);
    wire[0:0] s6878, in6878_1, in6878_2;
    wire c6878;
    assign in6878_1 = {c3941};
    assign in6878_2 = {c3942};
    Full_Adder FA_6878(s6878, c6878, in6878_1, in6878_2, c3940);
    wire[0:0] s6879, in6879_1, in6879_2;
    wire c6879;
    assign in6879_1 = {c3944};
    assign in6879_2 = {c3945};
    Full_Adder FA_6879(s6879, c6879, in6879_1, in6879_2, c3943);
    wire[0:0] s6880, in6880_1, in6880_2;
    wire c6880;
    assign in6880_1 = {c3947};
    assign in6880_2 = {c3948};
    Full_Adder FA_6880(s6880, c6880, in6880_1, in6880_2, c3946);
    wire[0:0] s6881, in6881_1, in6881_2;
    wire c6881;
    assign in6881_1 = {s3950[0]};
    assign in6881_2 = {s3951[0]};
    Full_Adder FA_6881(s6881, c6881, in6881_1, in6881_2, s3949[0]);
    wire[0:0] s6882, in6882_1, in6882_2;
    wire c6882;
    assign in6882_1 = {s3953[0]};
    assign in6882_2 = {s3954[0]};
    Full_Adder FA_6882(s6882, c6882, in6882_1, in6882_2, s3952[0]);
    wire[0:0] s6883, in6883_1, in6883_2;
    wire c6883;
    assign in6883_1 = {s3956[0]};
    assign in6883_2 = {s3957[0]};
    Full_Adder FA_6883(s6883, c6883, in6883_1, in6883_2, s3955[0]);
    wire[0:0] s6884, in6884_1, in6884_2;
    wire c6884;
    assign in6884_1 = {s3959[0]};
    assign in6884_2 = {s3960[0]};
    Full_Adder FA_6884(s6884, c6884, in6884_1, in6884_2, s3958[0]);
    wire[0:0] s6885, in6885_1, in6885_2;
    wire c6885;
    assign in6885_1 = {s3962[0]};
    assign in6885_2 = {s3963[0]};
    Full_Adder FA_6885(s6885, c6885, in6885_1, in6885_2, s3961[0]);
    wire[0:0] s6886, in6886_1, in6886_2;
    wire c6886;
    assign in6886_1 = {s3965[0]};
    assign in6886_2 = {s3966[0]};
    Full_Adder FA_6886(s6886, c6886, in6886_1, in6886_2, s3964[0]);
    wire[0:0] s6887, in6887_1, in6887_2;
    wire c6887;
    assign in6887_1 = {s3968[0]};
    assign in6887_2 = {s3969[0]};
    Full_Adder FA_6887(s6887, c6887, in6887_1, in6887_2, s3967[0]);
    wire[0:0] s6888, in6888_1, in6888_2;
    wire c6888;
    assign in6888_1 = {s3971[0]};
    assign in6888_2 = {s3972[0]};
    Full_Adder FA_6888(s6888, c6888, in6888_1, in6888_2, s3970[0]);
    wire[0:0] s6889, in6889_1, in6889_2;
    wire c6889;
    assign in6889_1 = {s3974[0]};
    assign in6889_2 = {s3975[0]};
    Full_Adder FA_6889(s6889, c6889, in6889_1, in6889_2, s3973[0]);
    wire[0:0] s6890, in6890_1, in6890_2;
    wire c6890;
    assign in6890_1 = {s1596[0]};
    assign in6890_2 = {c3949};
    Full_Adder FA_6890(s6890, c6890, in6890_1, in6890_2, s1595[0]);
    wire[0:0] s6891, in6891_1, in6891_2;
    wire c6891;
    assign in6891_1 = {c3951};
    assign in6891_2 = {c3952};
    Full_Adder FA_6891(s6891, c6891, in6891_1, in6891_2, c3950);
    wire[0:0] s6892, in6892_1, in6892_2;
    wire c6892;
    assign in6892_1 = {c3954};
    assign in6892_2 = {c3955};
    Full_Adder FA_6892(s6892, c6892, in6892_1, in6892_2, c3953);
    wire[0:0] s6893, in6893_1, in6893_2;
    wire c6893;
    assign in6893_1 = {c3957};
    assign in6893_2 = {c3958};
    Full_Adder FA_6893(s6893, c6893, in6893_1, in6893_2, c3956);
    wire[0:0] s6894, in6894_1, in6894_2;
    wire c6894;
    assign in6894_1 = {c3960};
    assign in6894_2 = {c3961};
    Full_Adder FA_6894(s6894, c6894, in6894_1, in6894_2, c3959);
    wire[0:0] s6895, in6895_1, in6895_2;
    wire c6895;
    assign in6895_1 = {c3963};
    assign in6895_2 = {c3964};
    Full_Adder FA_6895(s6895, c6895, in6895_1, in6895_2, c3962);
    wire[0:0] s6896, in6896_1, in6896_2;
    wire c6896;
    assign in6896_1 = {c3966};
    assign in6896_2 = {c3967};
    Full_Adder FA_6896(s6896, c6896, in6896_1, in6896_2, c3965);
    wire[0:0] s6897, in6897_1, in6897_2;
    wire c6897;
    assign in6897_1 = {c3969};
    assign in6897_2 = {c3970};
    Full_Adder FA_6897(s6897, c6897, in6897_1, in6897_2, c3968);
    wire[0:0] s6898, in6898_1, in6898_2;
    wire c6898;
    assign in6898_1 = {c3972};
    assign in6898_2 = {c3973};
    Full_Adder FA_6898(s6898, c6898, in6898_1, in6898_2, c3971);
    wire[0:0] s6899, in6899_1, in6899_2;
    wire c6899;
    assign in6899_1 = {c3975};
    assign in6899_2 = {c3976};
    Full_Adder FA_6899(s6899, c6899, in6899_1, in6899_2, c3974);
    wire[0:0] s6900, in6900_1, in6900_2;
    wire c6900;
    assign in6900_1 = {s3978[0]};
    assign in6900_2 = {s3979[0]};
    Full_Adder FA_6900(s6900, c6900, in6900_1, in6900_2, s3977[0]);
    wire[0:0] s6901, in6901_1, in6901_2;
    wire c6901;
    assign in6901_1 = {s3981[0]};
    assign in6901_2 = {s3982[0]};
    Full_Adder FA_6901(s6901, c6901, in6901_1, in6901_2, s3980[0]);
    wire[0:0] s6902, in6902_1, in6902_2;
    wire c6902;
    assign in6902_1 = {s3984[0]};
    assign in6902_2 = {s3985[0]};
    Full_Adder FA_6902(s6902, c6902, in6902_1, in6902_2, s3983[0]);
    wire[0:0] s6903, in6903_1, in6903_2;
    wire c6903;
    assign in6903_1 = {s3987[0]};
    assign in6903_2 = {s3988[0]};
    Full_Adder FA_6903(s6903, c6903, in6903_1, in6903_2, s3986[0]);
    wire[0:0] s6904, in6904_1, in6904_2;
    wire c6904;
    assign in6904_1 = {s3990[0]};
    assign in6904_2 = {s3991[0]};
    Full_Adder FA_6904(s6904, c6904, in6904_1, in6904_2, s3989[0]);
    wire[0:0] s6905, in6905_1, in6905_2;
    wire c6905;
    assign in6905_1 = {s3993[0]};
    assign in6905_2 = {s3994[0]};
    Full_Adder FA_6905(s6905, c6905, in6905_1, in6905_2, s3992[0]);
    wire[0:0] s6906, in6906_1, in6906_2;
    wire c6906;
    assign in6906_1 = {s3996[0]};
    assign in6906_2 = {s3997[0]};
    Full_Adder FA_6906(s6906, c6906, in6906_1, in6906_2, s3995[0]);
    wire[0:0] s6907, in6907_1, in6907_2;
    wire c6907;
    assign in6907_1 = {s3999[0]};
    assign in6907_2 = {s4000[0]};
    Full_Adder FA_6907(s6907, c6907, in6907_1, in6907_2, s3998[0]);
    wire[0:0] s6908, in6908_1, in6908_2;
    wire c6908;
    assign in6908_1 = {s4002[0]};
    assign in6908_2 = {s4003[0]};
    Full_Adder FA_6908(s6908, c6908, in6908_1, in6908_2, s4001[0]);
    wire[0:0] s6909, in6909_1, in6909_2;
    wire c6909;
    assign in6909_1 = {s1616[0]};
    assign in6909_2 = {c3977};
    Full_Adder FA_6909(s6909, c6909, in6909_1, in6909_2, s1615[0]);
    wire[0:0] s6910, in6910_1, in6910_2;
    wire c6910;
    assign in6910_1 = {c3979};
    assign in6910_2 = {c3980};
    Full_Adder FA_6910(s6910, c6910, in6910_1, in6910_2, c3978);
    wire[0:0] s6911, in6911_1, in6911_2;
    wire c6911;
    assign in6911_1 = {c3982};
    assign in6911_2 = {c3983};
    Full_Adder FA_6911(s6911, c6911, in6911_1, in6911_2, c3981);
    wire[0:0] s6912, in6912_1, in6912_2;
    wire c6912;
    assign in6912_1 = {c3985};
    assign in6912_2 = {c3986};
    Full_Adder FA_6912(s6912, c6912, in6912_1, in6912_2, c3984);
    wire[0:0] s6913, in6913_1, in6913_2;
    wire c6913;
    assign in6913_1 = {c3988};
    assign in6913_2 = {c3989};
    Full_Adder FA_6913(s6913, c6913, in6913_1, in6913_2, c3987);
    wire[0:0] s6914, in6914_1, in6914_2;
    wire c6914;
    assign in6914_1 = {c3991};
    assign in6914_2 = {c3992};
    Full_Adder FA_6914(s6914, c6914, in6914_1, in6914_2, c3990);
    wire[0:0] s6915, in6915_1, in6915_2;
    wire c6915;
    assign in6915_1 = {c3994};
    assign in6915_2 = {c3995};
    Full_Adder FA_6915(s6915, c6915, in6915_1, in6915_2, c3993);
    wire[0:0] s6916, in6916_1, in6916_2;
    wire c6916;
    assign in6916_1 = {c3997};
    assign in6916_2 = {c3998};
    Full_Adder FA_6916(s6916, c6916, in6916_1, in6916_2, c3996);
    wire[0:0] s6917, in6917_1, in6917_2;
    wire c6917;
    assign in6917_1 = {c4000};
    assign in6917_2 = {c4001};
    Full_Adder FA_6917(s6917, c6917, in6917_1, in6917_2, c3999);
    wire[0:0] s6918, in6918_1, in6918_2;
    wire c6918;
    assign in6918_1 = {c4003};
    assign in6918_2 = {c4004};
    Full_Adder FA_6918(s6918, c6918, in6918_1, in6918_2, c4002);
    wire[0:0] s6919, in6919_1, in6919_2;
    wire c6919;
    assign in6919_1 = {s4006[0]};
    assign in6919_2 = {s4007[0]};
    Full_Adder FA_6919(s6919, c6919, in6919_1, in6919_2, s4005[0]);
    wire[0:0] s6920, in6920_1, in6920_2;
    wire c6920;
    assign in6920_1 = {s4009[0]};
    assign in6920_2 = {s4010[0]};
    Full_Adder FA_6920(s6920, c6920, in6920_1, in6920_2, s4008[0]);
    wire[0:0] s6921, in6921_1, in6921_2;
    wire c6921;
    assign in6921_1 = {s4012[0]};
    assign in6921_2 = {s4013[0]};
    Full_Adder FA_6921(s6921, c6921, in6921_1, in6921_2, s4011[0]);
    wire[0:0] s6922, in6922_1, in6922_2;
    wire c6922;
    assign in6922_1 = {s4015[0]};
    assign in6922_2 = {s4016[0]};
    Full_Adder FA_6922(s6922, c6922, in6922_1, in6922_2, s4014[0]);
    wire[0:0] s6923, in6923_1, in6923_2;
    wire c6923;
    assign in6923_1 = {s4018[0]};
    assign in6923_2 = {s4019[0]};
    Full_Adder FA_6923(s6923, c6923, in6923_1, in6923_2, s4017[0]);
    wire[0:0] s6924, in6924_1, in6924_2;
    wire c6924;
    assign in6924_1 = {s4021[0]};
    assign in6924_2 = {s4022[0]};
    Full_Adder FA_6924(s6924, c6924, in6924_1, in6924_2, s4020[0]);
    wire[0:0] s6925, in6925_1, in6925_2;
    wire c6925;
    assign in6925_1 = {s4024[0]};
    assign in6925_2 = {s4025[0]};
    Full_Adder FA_6925(s6925, c6925, in6925_1, in6925_2, s4023[0]);
    wire[0:0] s6926, in6926_1, in6926_2;
    wire c6926;
    assign in6926_1 = {s4027[0]};
    assign in6926_2 = {s4028[0]};
    Full_Adder FA_6926(s6926, c6926, in6926_1, in6926_2, s4026[0]);
    wire[0:0] s6927, in6927_1, in6927_2;
    wire c6927;
    assign in6927_1 = {s4030[0]};
    assign in6927_2 = {s4031[0]};
    Full_Adder FA_6927(s6927, c6927, in6927_1, in6927_2, s4029[0]);
    wire[0:0] s6928, in6928_1, in6928_2;
    wire c6928;
    assign in6928_1 = {s1635[0]};
    assign in6928_2 = {c4005};
    Full_Adder FA_6928(s6928, c6928, in6928_1, in6928_2, s1634[0]);
    wire[0:0] s6929, in6929_1, in6929_2;
    wire c6929;
    assign in6929_1 = {c4007};
    assign in6929_2 = {c4008};
    Full_Adder FA_6929(s6929, c6929, in6929_1, in6929_2, c4006);
    wire[0:0] s6930, in6930_1, in6930_2;
    wire c6930;
    assign in6930_1 = {c4010};
    assign in6930_2 = {c4011};
    Full_Adder FA_6930(s6930, c6930, in6930_1, in6930_2, c4009);
    wire[0:0] s6931, in6931_1, in6931_2;
    wire c6931;
    assign in6931_1 = {c4013};
    assign in6931_2 = {c4014};
    Full_Adder FA_6931(s6931, c6931, in6931_1, in6931_2, c4012);
    wire[0:0] s6932, in6932_1, in6932_2;
    wire c6932;
    assign in6932_1 = {c4016};
    assign in6932_2 = {c4017};
    Full_Adder FA_6932(s6932, c6932, in6932_1, in6932_2, c4015);
    wire[0:0] s6933, in6933_1, in6933_2;
    wire c6933;
    assign in6933_1 = {c4019};
    assign in6933_2 = {c4020};
    Full_Adder FA_6933(s6933, c6933, in6933_1, in6933_2, c4018);
    wire[0:0] s6934, in6934_1, in6934_2;
    wire c6934;
    assign in6934_1 = {c4022};
    assign in6934_2 = {c4023};
    Full_Adder FA_6934(s6934, c6934, in6934_1, in6934_2, c4021);
    wire[0:0] s6935, in6935_1, in6935_2;
    wire c6935;
    assign in6935_1 = {c4025};
    assign in6935_2 = {c4026};
    Full_Adder FA_6935(s6935, c6935, in6935_1, in6935_2, c4024);
    wire[0:0] s6936, in6936_1, in6936_2;
    wire c6936;
    assign in6936_1 = {c4028};
    assign in6936_2 = {c4029};
    Full_Adder FA_6936(s6936, c6936, in6936_1, in6936_2, c4027);
    wire[0:0] s6937, in6937_1, in6937_2;
    wire c6937;
    assign in6937_1 = {c4031};
    assign in6937_2 = {c4032};
    Full_Adder FA_6937(s6937, c6937, in6937_1, in6937_2, c4030);
    wire[0:0] s6938, in6938_1, in6938_2;
    wire c6938;
    assign in6938_1 = {s4034[0]};
    assign in6938_2 = {s4035[0]};
    Full_Adder FA_6938(s6938, c6938, in6938_1, in6938_2, s4033[0]);
    wire[0:0] s6939, in6939_1, in6939_2;
    wire c6939;
    assign in6939_1 = {s4037[0]};
    assign in6939_2 = {s4038[0]};
    Full_Adder FA_6939(s6939, c6939, in6939_1, in6939_2, s4036[0]);
    wire[0:0] s6940, in6940_1, in6940_2;
    wire c6940;
    assign in6940_1 = {s4040[0]};
    assign in6940_2 = {s4041[0]};
    Full_Adder FA_6940(s6940, c6940, in6940_1, in6940_2, s4039[0]);
    wire[0:0] s6941, in6941_1, in6941_2;
    wire c6941;
    assign in6941_1 = {s4043[0]};
    assign in6941_2 = {s4044[0]};
    Full_Adder FA_6941(s6941, c6941, in6941_1, in6941_2, s4042[0]);
    wire[0:0] s6942, in6942_1, in6942_2;
    wire c6942;
    assign in6942_1 = {s4046[0]};
    assign in6942_2 = {s4047[0]};
    Full_Adder FA_6942(s6942, c6942, in6942_1, in6942_2, s4045[0]);
    wire[0:0] s6943, in6943_1, in6943_2;
    wire c6943;
    assign in6943_1 = {s4049[0]};
    assign in6943_2 = {s4050[0]};
    Full_Adder FA_6943(s6943, c6943, in6943_1, in6943_2, s4048[0]);
    wire[0:0] s6944, in6944_1, in6944_2;
    wire c6944;
    assign in6944_1 = {s4052[0]};
    assign in6944_2 = {s4053[0]};
    Full_Adder FA_6944(s6944, c6944, in6944_1, in6944_2, s4051[0]);
    wire[0:0] s6945, in6945_1, in6945_2;
    wire c6945;
    assign in6945_1 = {s4055[0]};
    assign in6945_2 = {s4056[0]};
    Full_Adder FA_6945(s6945, c6945, in6945_1, in6945_2, s4054[0]);
    wire[0:0] s6946, in6946_1, in6946_2;
    wire c6946;
    assign in6946_1 = {s4058[0]};
    assign in6946_2 = {s4059[0]};
    Full_Adder FA_6946(s6946, c6946, in6946_1, in6946_2, s4057[0]);
    wire[0:0] s6947, in6947_1, in6947_2;
    wire c6947;
    assign in6947_1 = {s1653[0]};
    assign in6947_2 = {c4033};
    Full_Adder FA_6947(s6947, c6947, in6947_1, in6947_2, s1652[0]);
    wire[0:0] s6948, in6948_1, in6948_2;
    wire c6948;
    assign in6948_1 = {c4035};
    assign in6948_2 = {c4036};
    Full_Adder FA_6948(s6948, c6948, in6948_1, in6948_2, c4034);
    wire[0:0] s6949, in6949_1, in6949_2;
    wire c6949;
    assign in6949_1 = {c4038};
    assign in6949_2 = {c4039};
    Full_Adder FA_6949(s6949, c6949, in6949_1, in6949_2, c4037);
    wire[0:0] s6950, in6950_1, in6950_2;
    wire c6950;
    assign in6950_1 = {c4041};
    assign in6950_2 = {c4042};
    Full_Adder FA_6950(s6950, c6950, in6950_1, in6950_2, c4040);
    wire[0:0] s6951, in6951_1, in6951_2;
    wire c6951;
    assign in6951_1 = {c4044};
    assign in6951_2 = {c4045};
    Full_Adder FA_6951(s6951, c6951, in6951_1, in6951_2, c4043);
    wire[0:0] s6952, in6952_1, in6952_2;
    wire c6952;
    assign in6952_1 = {c4047};
    assign in6952_2 = {c4048};
    Full_Adder FA_6952(s6952, c6952, in6952_1, in6952_2, c4046);
    wire[0:0] s6953, in6953_1, in6953_2;
    wire c6953;
    assign in6953_1 = {c4050};
    assign in6953_2 = {c4051};
    Full_Adder FA_6953(s6953, c6953, in6953_1, in6953_2, c4049);
    wire[0:0] s6954, in6954_1, in6954_2;
    wire c6954;
    assign in6954_1 = {c4053};
    assign in6954_2 = {c4054};
    Full_Adder FA_6954(s6954, c6954, in6954_1, in6954_2, c4052);
    wire[0:0] s6955, in6955_1, in6955_2;
    wire c6955;
    assign in6955_1 = {c4056};
    assign in6955_2 = {c4057};
    Full_Adder FA_6955(s6955, c6955, in6955_1, in6955_2, c4055);
    wire[0:0] s6956, in6956_1, in6956_2;
    wire c6956;
    assign in6956_1 = {c4059};
    assign in6956_2 = {c4060};
    Full_Adder FA_6956(s6956, c6956, in6956_1, in6956_2, c4058);
    wire[0:0] s6957, in6957_1, in6957_2;
    wire c6957;
    assign in6957_1 = {s4062[0]};
    assign in6957_2 = {s4063[0]};
    Full_Adder FA_6957(s6957, c6957, in6957_1, in6957_2, s4061[0]);
    wire[0:0] s6958, in6958_1, in6958_2;
    wire c6958;
    assign in6958_1 = {s4065[0]};
    assign in6958_2 = {s4066[0]};
    Full_Adder FA_6958(s6958, c6958, in6958_1, in6958_2, s4064[0]);
    wire[0:0] s6959, in6959_1, in6959_2;
    wire c6959;
    assign in6959_1 = {s4068[0]};
    assign in6959_2 = {s4069[0]};
    Full_Adder FA_6959(s6959, c6959, in6959_1, in6959_2, s4067[0]);
    wire[0:0] s6960, in6960_1, in6960_2;
    wire c6960;
    assign in6960_1 = {s4071[0]};
    assign in6960_2 = {s4072[0]};
    Full_Adder FA_6960(s6960, c6960, in6960_1, in6960_2, s4070[0]);
    wire[0:0] s6961, in6961_1, in6961_2;
    wire c6961;
    assign in6961_1 = {s4074[0]};
    assign in6961_2 = {s4075[0]};
    Full_Adder FA_6961(s6961, c6961, in6961_1, in6961_2, s4073[0]);
    wire[0:0] s6962, in6962_1, in6962_2;
    wire c6962;
    assign in6962_1 = {s4077[0]};
    assign in6962_2 = {s4078[0]};
    Full_Adder FA_6962(s6962, c6962, in6962_1, in6962_2, s4076[0]);
    wire[0:0] s6963, in6963_1, in6963_2;
    wire c6963;
    assign in6963_1 = {s4080[0]};
    assign in6963_2 = {s4081[0]};
    Full_Adder FA_6963(s6963, c6963, in6963_1, in6963_2, s4079[0]);
    wire[0:0] s6964, in6964_1, in6964_2;
    wire c6964;
    assign in6964_1 = {s4083[0]};
    assign in6964_2 = {s4084[0]};
    Full_Adder FA_6964(s6964, c6964, in6964_1, in6964_2, s4082[0]);
    wire[0:0] s6965, in6965_1, in6965_2;
    wire c6965;
    assign in6965_1 = {s4086[0]};
    assign in6965_2 = {s4087[0]};
    Full_Adder FA_6965(s6965, c6965, in6965_1, in6965_2, s4085[0]);
    wire[0:0] s6966, in6966_1, in6966_2;
    wire c6966;
    assign in6966_1 = {s1670[0]};
    assign in6966_2 = {c4061};
    Full_Adder FA_6966(s6966, c6966, in6966_1, in6966_2, s1669[0]);
    wire[0:0] s6967, in6967_1, in6967_2;
    wire c6967;
    assign in6967_1 = {c4063};
    assign in6967_2 = {c4064};
    Full_Adder FA_6967(s6967, c6967, in6967_1, in6967_2, c4062);
    wire[0:0] s6968, in6968_1, in6968_2;
    wire c6968;
    assign in6968_1 = {c4066};
    assign in6968_2 = {c4067};
    Full_Adder FA_6968(s6968, c6968, in6968_1, in6968_2, c4065);
    wire[0:0] s6969, in6969_1, in6969_2;
    wire c6969;
    assign in6969_1 = {c4069};
    assign in6969_2 = {c4070};
    Full_Adder FA_6969(s6969, c6969, in6969_1, in6969_2, c4068);
    wire[0:0] s6970, in6970_1, in6970_2;
    wire c6970;
    assign in6970_1 = {c4072};
    assign in6970_2 = {c4073};
    Full_Adder FA_6970(s6970, c6970, in6970_1, in6970_2, c4071);
    wire[0:0] s6971, in6971_1, in6971_2;
    wire c6971;
    assign in6971_1 = {c4075};
    assign in6971_2 = {c4076};
    Full_Adder FA_6971(s6971, c6971, in6971_1, in6971_2, c4074);
    wire[0:0] s6972, in6972_1, in6972_2;
    wire c6972;
    assign in6972_1 = {c4078};
    assign in6972_2 = {c4079};
    Full_Adder FA_6972(s6972, c6972, in6972_1, in6972_2, c4077);
    wire[0:0] s6973, in6973_1, in6973_2;
    wire c6973;
    assign in6973_1 = {c4081};
    assign in6973_2 = {c4082};
    Full_Adder FA_6973(s6973, c6973, in6973_1, in6973_2, c4080);
    wire[0:0] s6974, in6974_1, in6974_2;
    wire c6974;
    assign in6974_1 = {c4084};
    assign in6974_2 = {c4085};
    Full_Adder FA_6974(s6974, c6974, in6974_1, in6974_2, c4083);
    wire[0:0] s6975, in6975_1, in6975_2;
    wire c6975;
    assign in6975_1 = {c4087};
    assign in6975_2 = {c4088};
    Full_Adder FA_6975(s6975, c6975, in6975_1, in6975_2, c4086);
    wire[0:0] s6976, in6976_1, in6976_2;
    wire c6976;
    assign in6976_1 = {s4090[0]};
    assign in6976_2 = {s4091[0]};
    Full_Adder FA_6976(s6976, c6976, in6976_1, in6976_2, s4089[0]);
    wire[0:0] s6977, in6977_1, in6977_2;
    wire c6977;
    assign in6977_1 = {s4093[0]};
    assign in6977_2 = {s4094[0]};
    Full_Adder FA_6977(s6977, c6977, in6977_1, in6977_2, s4092[0]);
    wire[0:0] s6978, in6978_1, in6978_2;
    wire c6978;
    assign in6978_1 = {s4096[0]};
    assign in6978_2 = {s4097[0]};
    Full_Adder FA_6978(s6978, c6978, in6978_1, in6978_2, s4095[0]);
    wire[0:0] s6979, in6979_1, in6979_2;
    wire c6979;
    assign in6979_1 = {s4099[0]};
    assign in6979_2 = {s4100[0]};
    Full_Adder FA_6979(s6979, c6979, in6979_1, in6979_2, s4098[0]);
    wire[0:0] s6980, in6980_1, in6980_2;
    wire c6980;
    assign in6980_1 = {s4102[0]};
    assign in6980_2 = {s4103[0]};
    Full_Adder FA_6980(s6980, c6980, in6980_1, in6980_2, s4101[0]);
    wire[0:0] s6981, in6981_1, in6981_2;
    wire c6981;
    assign in6981_1 = {s4105[0]};
    assign in6981_2 = {s4106[0]};
    Full_Adder FA_6981(s6981, c6981, in6981_1, in6981_2, s4104[0]);
    wire[0:0] s6982, in6982_1, in6982_2;
    wire c6982;
    assign in6982_1 = {s4108[0]};
    assign in6982_2 = {s4109[0]};
    Full_Adder FA_6982(s6982, c6982, in6982_1, in6982_2, s4107[0]);
    wire[0:0] s6983, in6983_1, in6983_2;
    wire c6983;
    assign in6983_1 = {s4111[0]};
    assign in6983_2 = {s4112[0]};
    Full_Adder FA_6983(s6983, c6983, in6983_1, in6983_2, s4110[0]);
    wire[0:0] s6984, in6984_1, in6984_2;
    wire c6984;
    assign in6984_1 = {s4114[0]};
    assign in6984_2 = {s4115[0]};
    Full_Adder FA_6984(s6984, c6984, in6984_1, in6984_2, s4113[0]);
    wire[0:0] s6985, in6985_1, in6985_2;
    wire c6985;
    assign in6985_1 = {s1686[0]};
    assign in6985_2 = {c4089};
    Full_Adder FA_6985(s6985, c6985, in6985_1, in6985_2, s1685[0]);
    wire[0:0] s6986, in6986_1, in6986_2;
    wire c6986;
    assign in6986_1 = {c4091};
    assign in6986_2 = {c4092};
    Full_Adder FA_6986(s6986, c6986, in6986_1, in6986_2, c4090);
    wire[0:0] s6987, in6987_1, in6987_2;
    wire c6987;
    assign in6987_1 = {c4094};
    assign in6987_2 = {c4095};
    Full_Adder FA_6987(s6987, c6987, in6987_1, in6987_2, c4093);
    wire[0:0] s6988, in6988_1, in6988_2;
    wire c6988;
    assign in6988_1 = {c4097};
    assign in6988_2 = {c4098};
    Full_Adder FA_6988(s6988, c6988, in6988_1, in6988_2, c4096);
    wire[0:0] s6989, in6989_1, in6989_2;
    wire c6989;
    assign in6989_1 = {c4100};
    assign in6989_2 = {c4101};
    Full_Adder FA_6989(s6989, c6989, in6989_1, in6989_2, c4099);
    wire[0:0] s6990, in6990_1, in6990_2;
    wire c6990;
    assign in6990_1 = {c4103};
    assign in6990_2 = {c4104};
    Full_Adder FA_6990(s6990, c6990, in6990_1, in6990_2, c4102);
    wire[0:0] s6991, in6991_1, in6991_2;
    wire c6991;
    assign in6991_1 = {c4106};
    assign in6991_2 = {c4107};
    Full_Adder FA_6991(s6991, c6991, in6991_1, in6991_2, c4105);
    wire[0:0] s6992, in6992_1, in6992_2;
    wire c6992;
    assign in6992_1 = {c4109};
    assign in6992_2 = {c4110};
    Full_Adder FA_6992(s6992, c6992, in6992_1, in6992_2, c4108);
    wire[0:0] s6993, in6993_1, in6993_2;
    wire c6993;
    assign in6993_1 = {c4112};
    assign in6993_2 = {c4113};
    Full_Adder FA_6993(s6993, c6993, in6993_1, in6993_2, c4111);
    wire[0:0] s6994, in6994_1, in6994_2;
    wire c6994;
    assign in6994_1 = {c4115};
    assign in6994_2 = {c4116};
    Full_Adder FA_6994(s6994, c6994, in6994_1, in6994_2, c4114);
    wire[0:0] s6995, in6995_1, in6995_2;
    wire c6995;
    assign in6995_1 = {s4118[0]};
    assign in6995_2 = {s4119[0]};
    Full_Adder FA_6995(s6995, c6995, in6995_1, in6995_2, s4117[0]);
    wire[0:0] s6996, in6996_1, in6996_2;
    wire c6996;
    assign in6996_1 = {s4121[0]};
    assign in6996_2 = {s4122[0]};
    Full_Adder FA_6996(s6996, c6996, in6996_1, in6996_2, s4120[0]);
    wire[0:0] s6997, in6997_1, in6997_2;
    wire c6997;
    assign in6997_1 = {s4124[0]};
    assign in6997_2 = {s4125[0]};
    Full_Adder FA_6997(s6997, c6997, in6997_1, in6997_2, s4123[0]);
    wire[0:0] s6998, in6998_1, in6998_2;
    wire c6998;
    assign in6998_1 = {s4127[0]};
    assign in6998_2 = {s4128[0]};
    Full_Adder FA_6998(s6998, c6998, in6998_1, in6998_2, s4126[0]);
    wire[0:0] s6999, in6999_1, in6999_2;
    wire c6999;
    assign in6999_1 = {s4130[0]};
    assign in6999_2 = {s4131[0]};
    Full_Adder FA_6999(s6999, c6999, in6999_1, in6999_2, s4129[0]);
    wire[0:0] s7000, in7000_1, in7000_2;
    wire c7000;
    assign in7000_1 = {s4133[0]};
    assign in7000_2 = {s4134[0]};
    Full_Adder FA_7000(s7000, c7000, in7000_1, in7000_2, s4132[0]);
    wire[0:0] s7001, in7001_1, in7001_2;
    wire c7001;
    assign in7001_1 = {s4136[0]};
    assign in7001_2 = {s4137[0]};
    Full_Adder FA_7001(s7001, c7001, in7001_1, in7001_2, s4135[0]);
    wire[0:0] s7002, in7002_1, in7002_2;
    wire c7002;
    assign in7002_1 = {s4139[0]};
    assign in7002_2 = {s4140[0]};
    Full_Adder FA_7002(s7002, c7002, in7002_1, in7002_2, s4138[0]);
    wire[0:0] s7003, in7003_1, in7003_2;
    wire c7003;
    assign in7003_1 = {s4142[0]};
    assign in7003_2 = {s4143[0]};
    Full_Adder FA_7003(s7003, c7003, in7003_1, in7003_2, s4141[0]);
    wire[0:0] s7004, in7004_1, in7004_2;
    wire c7004;
    assign in7004_1 = {s1701[0]};
    assign in7004_2 = {c4117};
    Full_Adder FA_7004(s7004, c7004, in7004_1, in7004_2, s1700[0]);
    wire[0:0] s7005, in7005_1, in7005_2;
    wire c7005;
    assign in7005_1 = {c4119};
    assign in7005_2 = {c4120};
    Full_Adder FA_7005(s7005, c7005, in7005_1, in7005_2, c4118);
    wire[0:0] s7006, in7006_1, in7006_2;
    wire c7006;
    assign in7006_1 = {c4122};
    assign in7006_2 = {c4123};
    Full_Adder FA_7006(s7006, c7006, in7006_1, in7006_2, c4121);
    wire[0:0] s7007, in7007_1, in7007_2;
    wire c7007;
    assign in7007_1 = {c4125};
    assign in7007_2 = {c4126};
    Full_Adder FA_7007(s7007, c7007, in7007_1, in7007_2, c4124);
    wire[0:0] s7008, in7008_1, in7008_2;
    wire c7008;
    assign in7008_1 = {c4128};
    assign in7008_2 = {c4129};
    Full_Adder FA_7008(s7008, c7008, in7008_1, in7008_2, c4127);
    wire[0:0] s7009, in7009_1, in7009_2;
    wire c7009;
    assign in7009_1 = {c4131};
    assign in7009_2 = {c4132};
    Full_Adder FA_7009(s7009, c7009, in7009_1, in7009_2, c4130);
    wire[0:0] s7010, in7010_1, in7010_2;
    wire c7010;
    assign in7010_1 = {c4134};
    assign in7010_2 = {c4135};
    Full_Adder FA_7010(s7010, c7010, in7010_1, in7010_2, c4133);
    wire[0:0] s7011, in7011_1, in7011_2;
    wire c7011;
    assign in7011_1 = {c4137};
    assign in7011_2 = {c4138};
    Full_Adder FA_7011(s7011, c7011, in7011_1, in7011_2, c4136);
    wire[0:0] s7012, in7012_1, in7012_2;
    wire c7012;
    assign in7012_1 = {c4140};
    assign in7012_2 = {c4141};
    Full_Adder FA_7012(s7012, c7012, in7012_1, in7012_2, c4139);
    wire[0:0] s7013, in7013_1, in7013_2;
    wire c7013;
    assign in7013_1 = {c4143};
    assign in7013_2 = {c4144};
    Full_Adder FA_7013(s7013, c7013, in7013_1, in7013_2, c4142);
    wire[0:0] s7014, in7014_1, in7014_2;
    wire c7014;
    assign in7014_1 = {s4146[0]};
    assign in7014_2 = {s4147[0]};
    Full_Adder FA_7014(s7014, c7014, in7014_1, in7014_2, s4145[0]);
    wire[0:0] s7015, in7015_1, in7015_2;
    wire c7015;
    assign in7015_1 = {s4149[0]};
    assign in7015_2 = {s4150[0]};
    Full_Adder FA_7015(s7015, c7015, in7015_1, in7015_2, s4148[0]);
    wire[0:0] s7016, in7016_1, in7016_2;
    wire c7016;
    assign in7016_1 = {s4152[0]};
    assign in7016_2 = {s4153[0]};
    Full_Adder FA_7016(s7016, c7016, in7016_1, in7016_2, s4151[0]);
    wire[0:0] s7017, in7017_1, in7017_2;
    wire c7017;
    assign in7017_1 = {s4155[0]};
    assign in7017_2 = {s4156[0]};
    Full_Adder FA_7017(s7017, c7017, in7017_1, in7017_2, s4154[0]);
    wire[0:0] s7018, in7018_1, in7018_2;
    wire c7018;
    assign in7018_1 = {s4158[0]};
    assign in7018_2 = {s4159[0]};
    Full_Adder FA_7018(s7018, c7018, in7018_1, in7018_2, s4157[0]);
    wire[0:0] s7019, in7019_1, in7019_2;
    wire c7019;
    assign in7019_1 = {s4161[0]};
    assign in7019_2 = {s4162[0]};
    Full_Adder FA_7019(s7019, c7019, in7019_1, in7019_2, s4160[0]);
    wire[0:0] s7020, in7020_1, in7020_2;
    wire c7020;
    assign in7020_1 = {s4164[0]};
    assign in7020_2 = {s4165[0]};
    Full_Adder FA_7020(s7020, c7020, in7020_1, in7020_2, s4163[0]);
    wire[0:0] s7021, in7021_1, in7021_2;
    wire c7021;
    assign in7021_1 = {s4167[0]};
    assign in7021_2 = {s4168[0]};
    Full_Adder FA_7021(s7021, c7021, in7021_1, in7021_2, s4166[0]);
    wire[0:0] s7022, in7022_1, in7022_2;
    wire c7022;
    assign in7022_1 = {s4170[0]};
    assign in7022_2 = {s4171[0]};
    Full_Adder FA_7022(s7022, c7022, in7022_1, in7022_2, s4169[0]);
    wire[0:0] s7023, in7023_1, in7023_2;
    wire c7023;
    assign in7023_1 = {s1715[0]};
    assign in7023_2 = {c4145};
    Full_Adder FA_7023(s7023, c7023, in7023_1, in7023_2, s1714[0]);
    wire[0:0] s7024, in7024_1, in7024_2;
    wire c7024;
    assign in7024_1 = {c4147};
    assign in7024_2 = {c4148};
    Full_Adder FA_7024(s7024, c7024, in7024_1, in7024_2, c4146);
    wire[0:0] s7025, in7025_1, in7025_2;
    wire c7025;
    assign in7025_1 = {c4150};
    assign in7025_2 = {c4151};
    Full_Adder FA_7025(s7025, c7025, in7025_1, in7025_2, c4149);
    wire[0:0] s7026, in7026_1, in7026_2;
    wire c7026;
    assign in7026_1 = {c4153};
    assign in7026_2 = {c4154};
    Full_Adder FA_7026(s7026, c7026, in7026_1, in7026_2, c4152);
    wire[0:0] s7027, in7027_1, in7027_2;
    wire c7027;
    assign in7027_1 = {c4156};
    assign in7027_2 = {c4157};
    Full_Adder FA_7027(s7027, c7027, in7027_1, in7027_2, c4155);
    wire[0:0] s7028, in7028_1, in7028_2;
    wire c7028;
    assign in7028_1 = {c4159};
    assign in7028_2 = {c4160};
    Full_Adder FA_7028(s7028, c7028, in7028_1, in7028_2, c4158);
    wire[0:0] s7029, in7029_1, in7029_2;
    wire c7029;
    assign in7029_1 = {c4162};
    assign in7029_2 = {c4163};
    Full_Adder FA_7029(s7029, c7029, in7029_1, in7029_2, c4161);
    wire[0:0] s7030, in7030_1, in7030_2;
    wire c7030;
    assign in7030_1 = {c4165};
    assign in7030_2 = {c4166};
    Full_Adder FA_7030(s7030, c7030, in7030_1, in7030_2, c4164);
    wire[0:0] s7031, in7031_1, in7031_2;
    wire c7031;
    assign in7031_1 = {c4168};
    assign in7031_2 = {c4169};
    Full_Adder FA_7031(s7031, c7031, in7031_1, in7031_2, c4167);
    wire[0:0] s7032, in7032_1, in7032_2;
    wire c7032;
    assign in7032_1 = {c4171};
    assign in7032_2 = {c4172};
    Full_Adder FA_7032(s7032, c7032, in7032_1, in7032_2, c4170);
    wire[0:0] s7033, in7033_1, in7033_2;
    wire c7033;
    assign in7033_1 = {s4174[0]};
    assign in7033_2 = {s4175[0]};
    Full_Adder FA_7033(s7033, c7033, in7033_1, in7033_2, s4173[0]);
    wire[0:0] s7034, in7034_1, in7034_2;
    wire c7034;
    assign in7034_1 = {s4177[0]};
    assign in7034_2 = {s4178[0]};
    Full_Adder FA_7034(s7034, c7034, in7034_1, in7034_2, s4176[0]);
    wire[0:0] s7035, in7035_1, in7035_2;
    wire c7035;
    assign in7035_1 = {s4180[0]};
    assign in7035_2 = {s4181[0]};
    Full_Adder FA_7035(s7035, c7035, in7035_1, in7035_2, s4179[0]);
    wire[0:0] s7036, in7036_1, in7036_2;
    wire c7036;
    assign in7036_1 = {s4183[0]};
    assign in7036_2 = {s4184[0]};
    Full_Adder FA_7036(s7036, c7036, in7036_1, in7036_2, s4182[0]);
    wire[0:0] s7037, in7037_1, in7037_2;
    wire c7037;
    assign in7037_1 = {s4186[0]};
    assign in7037_2 = {s4187[0]};
    Full_Adder FA_7037(s7037, c7037, in7037_1, in7037_2, s4185[0]);
    wire[0:0] s7038, in7038_1, in7038_2;
    wire c7038;
    assign in7038_1 = {s4189[0]};
    assign in7038_2 = {s4190[0]};
    Full_Adder FA_7038(s7038, c7038, in7038_1, in7038_2, s4188[0]);
    wire[0:0] s7039, in7039_1, in7039_2;
    wire c7039;
    assign in7039_1 = {s4192[0]};
    assign in7039_2 = {s4193[0]};
    Full_Adder FA_7039(s7039, c7039, in7039_1, in7039_2, s4191[0]);
    wire[0:0] s7040, in7040_1, in7040_2;
    wire c7040;
    assign in7040_1 = {s4195[0]};
    assign in7040_2 = {s4196[0]};
    Full_Adder FA_7040(s7040, c7040, in7040_1, in7040_2, s4194[0]);
    wire[0:0] s7041, in7041_1, in7041_2;
    wire c7041;
    assign in7041_1 = {s4198[0]};
    assign in7041_2 = {s4199[0]};
    Full_Adder FA_7041(s7041, c7041, in7041_1, in7041_2, s4197[0]);
    wire[0:0] s7042, in7042_1, in7042_2;
    wire c7042;
    assign in7042_1 = {s1728[0]};
    assign in7042_2 = {c4173};
    Full_Adder FA_7042(s7042, c7042, in7042_1, in7042_2, s1727[0]);
    wire[0:0] s7043, in7043_1, in7043_2;
    wire c7043;
    assign in7043_1 = {c4175};
    assign in7043_2 = {c4176};
    Full_Adder FA_7043(s7043, c7043, in7043_1, in7043_2, c4174);
    wire[0:0] s7044, in7044_1, in7044_2;
    wire c7044;
    assign in7044_1 = {c4178};
    assign in7044_2 = {c4179};
    Full_Adder FA_7044(s7044, c7044, in7044_1, in7044_2, c4177);
    wire[0:0] s7045, in7045_1, in7045_2;
    wire c7045;
    assign in7045_1 = {c4181};
    assign in7045_2 = {c4182};
    Full_Adder FA_7045(s7045, c7045, in7045_1, in7045_2, c4180);
    wire[0:0] s7046, in7046_1, in7046_2;
    wire c7046;
    assign in7046_1 = {c4184};
    assign in7046_2 = {c4185};
    Full_Adder FA_7046(s7046, c7046, in7046_1, in7046_2, c4183);
    wire[0:0] s7047, in7047_1, in7047_2;
    wire c7047;
    assign in7047_1 = {c4187};
    assign in7047_2 = {c4188};
    Full_Adder FA_7047(s7047, c7047, in7047_1, in7047_2, c4186);
    wire[0:0] s7048, in7048_1, in7048_2;
    wire c7048;
    assign in7048_1 = {c4190};
    assign in7048_2 = {c4191};
    Full_Adder FA_7048(s7048, c7048, in7048_1, in7048_2, c4189);
    wire[0:0] s7049, in7049_1, in7049_2;
    wire c7049;
    assign in7049_1 = {c4193};
    assign in7049_2 = {c4194};
    Full_Adder FA_7049(s7049, c7049, in7049_1, in7049_2, c4192);
    wire[0:0] s7050, in7050_1, in7050_2;
    wire c7050;
    assign in7050_1 = {c4196};
    assign in7050_2 = {c4197};
    Full_Adder FA_7050(s7050, c7050, in7050_1, in7050_2, c4195);
    wire[0:0] s7051, in7051_1, in7051_2;
    wire c7051;
    assign in7051_1 = {c4199};
    assign in7051_2 = {c4200};
    Full_Adder FA_7051(s7051, c7051, in7051_1, in7051_2, c4198);
    wire[0:0] s7052, in7052_1, in7052_2;
    wire c7052;
    assign in7052_1 = {s4202[0]};
    assign in7052_2 = {s4203[0]};
    Full_Adder FA_7052(s7052, c7052, in7052_1, in7052_2, s4201[0]);
    wire[0:0] s7053, in7053_1, in7053_2;
    wire c7053;
    assign in7053_1 = {s4205[0]};
    assign in7053_2 = {s4206[0]};
    Full_Adder FA_7053(s7053, c7053, in7053_1, in7053_2, s4204[0]);
    wire[0:0] s7054, in7054_1, in7054_2;
    wire c7054;
    assign in7054_1 = {s4208[0]};
    assign in7054_2 = {s4209[0]};
    Full_Adder FA_7054(s7054, c7054, in7054_1, in7054_2, s4207[0]);
    wire[0:0] s7055, in7055_1, in7055_2;
    wire c7055;
    assign in7055_1 = {s4211[0]};
    assign in7055_2 = {s4212[0]};
    Full_Adder FA_7055(s7055, c7055, in7055_1, in7055_2, s4210[0]);
    wire[0:0] s7056, in7056_1, in7056_2;
    wire c7056;
    assign in7056_1 = {s4214[0]};
    assign in7056_2 = {s4215[0]};
    Full_Adder FA_7056(s7056, c7056, in7056_1, in7056_2, s4213[0]);
    wire[0:0] s7057, in7057_1, in7057_2;
    wire c7057;
    assign in7057_1 = {s4217[0]};
    assign in7057_2 = {s4218[0]};
    Full_Adder FA_7057(s7057, c7057, in7057_1, in7057_2, s4216[0]);
    wire[0:0] s7058, in7058_1, in7058_2;
    wire c7058;
    assign in7058_1 = {s4220[0]};
    assign in7058_2 = {s4221[0]};
    Full_Adder FA_7058(s7058, c7058, in7058_1, in7058_2, s4219[0]);
    wire[0:0] s7059, in7059_1, in7059_2;
    wire c7059;
    assign in7059_1 = {s4223[0]};
    assign in7059_2 = {s4224[0]};
    Full_Adder FA_7059(s7059, c7059, in7059_1, in7059_2, s4222[0]);
    wire[0:0] s7060, in7060_1, in7060_2;
    wire c7060;
    assign in7060_1 = {s4226[0]};
    assign in7060_2 = {s4227[0]};
    Full_Adder FA_7060(s7060, c7060, in7060_1, in7060_2, s4225[0]);
    wire[0:0] s7061, in7061_1, in7061_2;
    wire c7061;
    assign in7061_1 = {s1740[0]};
    assign in7061_2 = {c4201};
    Full_Adder FA_7061(s7061, c7061, in7061_1, in7061_2, s1739[0]);
    wire[0:0] s7062, in7062_1, in7062_2;
    wire c7062;
    assign in7062_1 = {c4203};
    assign in7062_2 = {c4204};
    Full_Adder FA_7062(s7062, c7062, in7062_1, in7062_2, c4202);
    wire[0:0] s7063, in7063_1, in7063_2;
    wire c7063;
    assign in7063_1 = {c4206};
    assign in7063_2 = {c4207};
    Full_Adder FA_7063(s7063, c7063, in7063_1, in7063_2, c4205);
    wire[0:0] s7064, in7064_1, in7064_2;
    wire c7064;
    assign in7064_1 = {c4209};
    assign in7064_2 = {c4210};
    Full_Adder FA_7064(s7064, c7064, in7064_1, in7064_2, c4208);
    wire[0:0] s7065, in7065_1, in7065_2;
    wire c7065;
    assign in7065_1 = {c4212};
    assign in7065_2 = {c4213};
    Full_Adder FA_7065(s7065, c7065, in7065_1, in7065_2, c4211);
    wire[0:0] s7066, in7066_1, in7066_2;
    wire c7066;
    assign in7066_1 = {c4215};
    assign in7066_2 = {c4216};
    Full_Adder FA_7066(s7066, c7066, in7066_1, in7066_2, c4214);
    wire[0:0] s7067, in7067_1, in7067_2;
    wire c7067;
    assign in7067_1 = {c4218};
    assign in7067_2 = {c4219};
    Full_Adder FA_7067(s7067, c7067, in7067_1, in7067_2, c4217);
    wire[0:0] s7068, in7068_1, in7068_2;
    wire c7068;
    assign in7068_1 = {c4221};
    assign in7068_2 = {c4222};
    Full_Adder FA_7068(s7068, c7068, in7068_1, in7068_2, c4220);
    wire[0:0] s7069, in7069_1, in7069_2;
    wire c7069;
    assign in7069_1 = {c4224};
    assign in7069_2 = {c4225};
    Full_Adder FA_7069(s7069, c7069, in7069_1, in7069_2, c4223);
    wire[0:0] s7070, in7070_1, in7070_2;
    wire c7070;
    assign in7070_1 = {c4227};
    assign in7070_2 = {c4228};
    Full_Adder FA_7070(s7070, c7070, in7070_1, in7070_2, c4226);
    wire[0:0] s7071, in7071_1, in7071_2;
    wire c7071;
    assign in7071_1 = {s4230[0]};
    assign in7071_2 = {s4231[0]};
    Full_Adder FA_7071(s7071, c7071, in7071_1, in7071_2, s4229[0]);
    wire[0:0] s7072, in7072_1, in7072_2;
    wire c7072;
    assign in7072_1 = {s4233[0]};
    assign in7072_2 = {s4234[0]};
    Full_Adder FA_7072(s7072, c7072, in7072_1, in7072_2, s4232[0]);
    wire[0:0] s7073, in7073_1, in7073_2;
    wire c7073;
    assign in7073_1 = {s4236[0]};
    assign in7073_2 = {s4237[0]};
    Full_Adder FA_7073(s7073, c7073, in7073_1, in7073_2, s4235[0]);
    wire[0:0] s7074, in7074_1, in7074_2;
    wire c7074;
    assign in7074_1 = {s4239[0]};
    assign in7074_2 = {s4240[0]};
    Full_Adder FA_7074(s7074, c7074, in7074_1, in7074_2, s4238[0]);
    wire[0:0] s7075, in7075_1, in7075_2;
    wire c7075;
    assign in7075_1 = {s4242[0]};
    assign in7075_2 = {s4243[0]};
    Full_Adder FA_7075(s7075, c7075, in7075_1, in7075_2, s4241[0]);
    wire[0:0] s7076, in7076_1, in7076_2;
    wire c7076;
    assign in7076_1 = {s4245[0]};
    assign in7076_2 = {s4246[0]};
    Full_Adder FA_7076(s7076, c7076, in7076_1, in7076_2, s4244[0]);
    wire[0:0] s7077, in7077_1, in7077_2;
    wire c7077;
    assign in7077_1 = {s4248[0]};
    assign in7077_2 = {s4249[0]};
    Full_Adder FA_7077(s7077, c7077, in7077_1, in7077_2, s4247[0]);
    wire[0:0] s7078, in7078_1, in7078_2;
    wire c7078;
    assign in7078_1 = {s4251[0]};
    assign in7078_2 = {s4252[0]};
    Full_Adder FA_7078(s7078, c7078, in7078_1, in7078_2, s4250[0]);
    wire[0:0] s7079, in7079_1, in7079_2;
    wire c7079;
    assign in7079_1 = {s4254[0]};
    assign in7079_2 = {s4255[0]};
    Full_Adder FA_7079(s7079, c7079, in7079_1, in7079_2, s4253[0]);
    wire[0:0] s7080, in7080_1, in7080_2;
    wire c7080;
    assign in7080_1 = {s1751[0]};
    assign in7080_2 = {c4229};
    Full_Adder FA_7080(s7080, c7080, in7080_1, in7080_2, s1750[0]);
    wire[0:0] s7081, in7081_1, in7081_2;
    wire c7081;
    assign in7081_1 = {c4231};
    assign in7081_2 = {c4232};
    Full_Adder FA_7081(s7081, c7081, in7081_1, in7081_2, c4230);
    wire[0:0] s7082, in7082_1, in7082_2;
    wire c7082;
    assign in7082_1 = {c4234};
    assign in7082_2 = {c4235};
    Full_Adder FA_7082(s7082, c7082, in7082_1, in7082_2, c4233);
    wire[0:0] s7083, in7083_1, in7083_2;
    wire c7083;
    assign in7083_1 = {c4237};
    assign in7083_2 = {c4238};
    Full_Adder FA_7083(s7083, c7083, in7083_1, in7083_2, c4236);
    wire[0:0] s7084, in7084_1, in7084_2;
    wire c7084;
    assign in7084_1 = {c4240};
    assign in7084_2 = {c4241};
    Full_Adder FA_7084(s7084, c7084, in7084_1, in7084_2, c4239);
    wire[0:0] s7085, in7085_1, in7085_2;
    wire c7085;
    assign in7085_1 = {c4243};
    assign in7085_2 = {c4244};
    Full_Adder FA_7085(s7085, c7085, in7085_1, in7085_2, c4242);
    wire[0:0] s7086, in7086_1, in7086_2;
    wire c7086;
    assign in7086_1 = {c4246};
    assign in7086_2 = {c4247};
    Full_Adder FA_7086(s7086, c7086, in7086_1, in7086_2, c4245);
    wire[0:0] s7087, in7087_1, in7087_2;
    wire c7087;
    assign in7087_1 = {c4249};
    assign in7087_2 = {c4250};
    Full_Adder FA_7087(s7087, c7087, in7087_1, in7087_2, c4248);
    wire[0:0] s7088, in7088_1, in7088_2;
    wire c7088;
    assign in7088_1 = {c4252};
    assign in7088_2 = {c4253};
    Full_Adder FA_7088(s7088, c7088, in7088_1, in7088_2, c4251);
    wire[0:0] s7089, in7089_1, in7089_2;
    wire c7089;
    assign in7089_1 = {c4255};
    assign in7089_2 = {c4256};
    Full_Adder FA_7089(s7089, c7089, in7089_1, in7089_2, c4254);
    wire[0:0] s7090, in7090_1, in7090_2;
    wire c7090;
    assign in7090_1 = {s4258[0]};
    assign in7090_2 = {s4259[0]};
    Full_Adder FA_7090(s7090, c7090, in7090_1, in7090_2, s4257[0]);
    wire[0:0] s7091, in7091_1, in7091_2;
    wire c7091;
    assign in7091_1 = {s4261[0]};
    assign in7091_2 = {s4262[0]};
    Full_Adder FA_7091(s7091, c7091, in7091_1, in7091_2, s4260[0]);
    wire[0:0] s7092, in7092_1, in7092_2;
    wire c7092;
    assign in7092_1 = {s4264[0]};
    assign in7092_2 = {s4265[0]};
    Full_Adder FA_7092(s7092, c7092, in7092_1, in7092_2, s4263[0]);
    wire[0:0] s7093, in7093_1, in7093_2;
    wire c7093;
    assign in7093_1 = {s4267[0]};
    assign in7093_2 = {s4268[0]};
    Full_Adder FA_7093(s7093, c7093, in7093_1, in7093_2, s4266[0]);
    wire[0:0] s7094, in7094_1, in7094_2;
    wire c7094;
    assign in7094_1 = {s4270[0]};
    assign in7094_2 = {s4271[0]};
    Full_Adder FA_7094(s7094, c7094, in7094_1, in7094_2, s4269[0]);
    wire[0:0] s7095, in7095_1, in7095_2;
    wire c7095;
    assign in7095_1 = {s4273[0]};
    assign in7095_2 = {s4274[0]};
    Full_Adder FA_7095(s7095, c7095, in7095_1, in7095_2, s4272[0]);
    wire[0:0] s7096, in7096_1, in7096_2;
    wire c7096;
    assign in7096_1 = {s4276[0]};
    assign in7096_2 = {s4277[0]};
    Full_Adder FA_7096(s7096, c7096, in7096_1, in7096_2, s4275[0]);
    wire[0:0] s7097, in7097_1, in7097_2;
    wire c7097;
    assign in7097_1 = {s4279[0]};
    assign in7097_2 = {s4280[0]};
    Full_Adder FA_7097(s7097, c7097, in7097_1, in7097_2, s4278[0]);
    wire[0:0] s7098, in7098_1, in7098_2;
    wire c7098;
    assign in7098_1 = {s4282[0]};
    assign in7098_2 = {s4283[0]};
    Full_Adder FA_7098(s7098, c7098, in7098_1, in7098_2, s4281[0]);
    wire[0:0] s7099, in7099_1, in7099_2;
    wire c7099;
    assign in7099_1 = {s1761[0]};
    assign in7099_2 = {c4257};
    Full_Adder FA_7099(s7099, c7099, in7099_1, in7099_2, s1760[0]);
    wire[0:0] s7100, in7100_1, in7100_2;
    wire c7100;
    assign in7100_1 = {c4259};
    assign in7100_2 = {c4260};
    Full_Adder FA_7100(s7100, c7100, in7100_1, in7100_2, c4258);
    wire[0:0] s7101, in7101_1, in7101_2;
    wire c7101;
    assign in7101_1 = {c4262};
    assign in7101_2 = {c4263};
    Full_Adder FA_7101(s7101, c7101, in7101_1, in7101_2, c4261);
    wire[0:0] s7102, in7102_1, in7102_2;
    wire c7102;
    assign in7102_1 = {c4265};
    assign in7102_2 = {c4266};
    Full_Adder FA_7102(s7102, c7102, in7102_1, in7102_2, c4264);
    wire[0:0] s7103, in7103_1, in7103_2;
    wire c7103;
    assign in7103_1 = {c4268};
    assign in7103_2 = {c4269};
    Full_Adder FA_7103(s7103, c7103, in7103_1, in7103_2, c4267);
    wire[0:0] s7104, in7104_1, in7104_2;
    wire c7104;
    assign in7104_1 = {c4271};
    assign in7104_2 = {c4272};
    Full_Adder FA_7104(s7104, c7104, in7104_1, in7104_2, c4270);
    wire[0:0] s7105, in7105_1, in7105_2;
    wire c7105;
    assign in7105_1 = {c4274};
    assign in7105_2 = {c4275};
    Full_Adder FA_7105(s7105, c7105, in7105_1, in7105_2, c4273);
    wire[0:0] s7106, in7106_1, in7106_2;
    wire c7106;
    assign in7106_1 = {c4277};
    assign in7106_2 = {c4278};
    Full_Adder FA_7106(s7106, c7106, in7106_1, in7106_2, c4276);
    wire[0:0] s7107, in7107_1, in7107_2;
    wire c7107;
    assign in7107_1 = {c4280};
    assign in7107_2 = {c4281};
    Full_Adder FA_7107(s7107, c7107, in7107_1, in7107_2, c4279);
    wire[0:0] s7108, in7108_1, in7108_2;
    wire c7108;
    assign in7108_1 = {c4283};
    assign in7108_2 = {c4284};
    Full_Adder FA_7108(s7108, c7108, in7108_1, in7108_2, c4282);
    wire[0:0] s7109, in7109_1, in7109_2;
    wire c7109;
    assign in7109_1 = {s4286[0]};
    assign in7109_2 = {s4287[0]};
    Full_Adder FA_7109(s7109, c7109, in7109_1, in7109_2, s4285[0]);
    wire[0:0] s7110, in7110_1, in7110_2;
    wire c7110;
    assign in7110_1 = {s4289[0]};
    assign in7110_2 = {s4290[0]};
    Full_Adder FA_7110(s7110, c7110, in7110_1, in7110_2, s4288[0]);
    wire[0:0] s7111, in7111_1, in7111_2;
    wire c7111;
    assign in7111_1 = {s4292[0]};
    assign in7111_2 = {s4293[0]};
    Full_Adder FA_7111(s7111, c7111, in7111_1, in7111_2, s4291[0]);
    wire[0:0] s7112, in7112_1, in7112_2;
    wire c7112;
    assign in7112_1 = {s4295[0]};
    assign in7112_2 = {s4296[0]};
    Full_Adder FA_7112(s7112, c7112, in7112_1, in7112_2, s4294[0]);
    wire[0:0] s7113, in7113_1, in7113_2;
    wire c7113;
    assign in7113_1 = {s4298[0]};
    assign in7113_2 = {s4299[0]};
    Full_Adder FA_7113(s7113, c7113, in7113_1, in7113_2, s4297[0]);
    wire[0:0] s7114, in7114_1, in7114_2;
    wire c7114;
    assign in7114_1 = {s4301[0]};
    assign in7114_2 = {s4302[0]};
    Full_Adder FA_7114(s7114, c7114, in7114_1, in7114_2, s4300[0]);
    wire[0:0] s7115, in7115_1, in7115_2;
    wire c7115;
    assign in7115_1 = {s4304[0]};
    assign in7115_2 = {s4305[0]};
    Full_Adder FA_7115(s7115, c7115, in7115_1, in7115_2, s4303[0]);
    wire[0:0] s7116, in7116_1, in7116_2;
    wire c7116;
    assign in7116_1 = {s4307[0]};
    assign in7116_2 = {s4308[0]};
    Full_Adder FA_7116(s7116, c7116, in7116_1, in7116_2, s4306[0]);
    wire[0:0] s7117, in7117_1, in7117_2;
    wire c7117;
    assign in7117_1 = {s4310[0]};
    assign in7117_2 = {s4311[0]};
    Full_Adder FA_7117(s7117, c7117, in7117_1, in7117_2, s4309[0]);
    wire[0:0] s7118, in7118_1, in7118_2;
    wire c7118;
    assign in7118_1 = {s1770[0]};
    assign in7118_2 = {c4285};
    Full_Adder FA_7118(s7118, c7118, in7118_1, in7118_2, s1769[0]);
    wire[0:0] s7119, in7119_1, in7119_2;
    wire c7119;
    assign in7119_1 = {c4287};
    assign in7119_2 = {c4288};
    Full_Adder FA_7119(s7119, c7119, in7119_1, in7119_2, c4286);
    wire[0:0] s7120, in7120_1, in7120_2;
    wire c7120;
    assign in7120_1 = {c4290};
    assign in7120_2 = {c4291};
    Full_Adder FA_7120(s7120, c7120, in7120_1, in7120_2, c4289);
    wire[0:0] s7121, in7121_1, in7121_2;
    wire c7121;
    assign in7121_1 = {c4293};
    assign in7121_2 = {c4294};
    Full_Adder FA_7121(s7121, c7121, in7121_1, in7121_2, c4292);
    wire[0:0] s7122, in7122_1, in7122_2;
    wire c7122;
    assign in7122_1 = {c4296};
    assign in7122_2 = {c4297};
    Full_Adder FA_7122(s7122, c7122, in7122_1, in7122_2, c4295);
    wire[0:0] s7123, in7123_1, in7123_2;
    wire c7123;
    assign in7123_1 = {c4299};
    assign in7123_2 = {c4300};
    Full_Adder FA_7123(s7123, c7123, in7123_1, in7123_2, c4298);
    wire[0:0] s7124, in7124_1, in7124_2;
    wire c7124;
    assign in7124_1 = {c4302};
    assign in7124_2 = {c4303};
    Full_Adder FA_7124(s7124, c7124, in7124_1, in7124_2, c4301);
    wire[0:0] s7125, in7125_1, in7125_2;
    wire c7125;
    assign in7125_1 = {c4305};
    assign in7125_2 = {c4306};
    Full_Adder FA_7125(s7125, c7125, in7125_1, in7125_2, c4304);
    wire[0:0] s7126, in7126_1, in7126_2;
    wire c7126;
    assign in7126_1 = {c4308};
    assign in7126_2 = {c4309};
    Full_Adder FA_7126(s7126, c7126, in7126_1, in7126_2, c4307);
    wire[0:0] s7127, in7127_1, in7127_2;
    wire c7127;
    assign in7127_1 = {c4311};
    assign in7127_2 = {c4312};
    Full_Adder FA_7127(s7127, c7127, in7127_1, in7127_2, c4310);
    wire[0:0] s7128, in7128_1, in7128_2;
    wire c7128;
    assign in7128_1 = {s4314[0]};
    assign in7128_2 = {s4315[0]};
    Full_Adder FA_7128(s7128, c7128, in7128_1, in7128_2, s4313[0]);
    wire[0:0] s7129, in7129_1, in7129_2;
    wire c7129;
    assign in7129_1 = {s4317[0]};
    assign in7129_2 = {s4318[0]};
    Full_Adder FA_7129(s7129, c7129, in7129_1, in7129_2, s4316[0]);
    wire[0:0] s7130, in7130_1, in7130_2;
    wire c7130;
    assign in7130_1 = {s4320[0]};
    assign in7130_2 = {s4321[0]};
    Full_Adder FA_7130(s7130, c7130, in7130_1, in7130_2, s4319[0]);
    wire[0:0] s7131, in7131_1, in7131_2;
    wire c7131;
    assign in7131_1 = {s4323[0]};
    assign in7131_2 = {s4324[0]};
    Full_Adder FA_7131(s7131, c7131, in7131_1, in7131_2, s4322[0]);
    wire[0:0] s7132, in7132_1, in7132_2;
    wire c7132;
    assign in7132_1 = {s4326[0]};
    assign in7132_2 = {s4327[0]};
    Full_Adder FA_7132(s7132, c7132, in7132_1, in7132_2, s4325[0]);
    wire[0:0] s7133, in7133_1, in7133_2;
    wire c7133;
    assign in7133_1 = {s4329[0]};
    assign in7133_2 = {s4330[0]};
    Full_Adder FA_7133(s7133, c7133, in7133_1, in7133_2, s4328[0]);
    wire[0:0] s7134, in7134_1, in7134_2;
    wire c7134;
    assign in7134_1 = {s4332[0]};
    assign in7134_2 = {s4333[0]};
    Full_Adder FA_7134(s7134, c7134, in7134_1, in7134_2, s4331[0]);
    wire[0:0] s7135, in7135_1, in7135_2;
    wire c7135;
    assign in7135_1 = {s4335[0]};
    assign in7135_2 = {s4336[0]};
    Full_Adder FA_7135(s7135, c7135, in7135_1, in7135_2, s4334[0]);
    wire[0:0] s7136, in7136_1, in7136_2;
    wire c7136;
    assign in7136_1 = {s4338[0]};
    assign in7136_2 = {s4339[0]};
    Full_Adder FA_7136(s7136, c7136, in7136_1, in7136_2, s4337[0]);
    wire[0:0] s7137, in7137_1, in7137_2;
    wire c7137;
    assign in7137_1 = {s1778[0]};
    assign in7137_2 = {c4313};
    Full_Adder FA_7137(s7137, c7137, in7137_1, in7137_2, s1777[0]);
    wire[0:0] s7138, in7138_1, in7138_2;
    wire c7138;
    assign in7138_1 = {c4315};
    assign in7138_2 = {c4316};
    Full_Adder FA_7138(s7138, c7138, in7138_1, in7138_2, c4314);
    wire[0:0] s7139, in7139_1, in7139_2;
    wire c7139;
    assign in7139_1 = {c4318};
    assign in7139_2 = {c4319};
    Full_Adder FA_7139(s7139, c7139, in7139_1, in7139_2, c4317);
    wire[0:0] s7140, in7140_1, in7140_2;
    wire c7140;
    assign in7140_1 = {c4321};
    assign in7140_2 = {c4322};
    Full_Adder FA_7140(s7140, c7140, in7140_1, in7140_2, c4320);
    wire[0:0] s7141, in7141_1, in7141_2;
    wire c7141;
    assign in7141_1 = {c4324};
    assign in7141_2 = {c4325};
    Full_Adder FA_7141(s7141, c7141, in7141_1, in7141_2, c4323);
    wire[0:0] s7142, in7142_1, in7142_2;
    wire c7142;
    assign in7142_1 = {c4327};
    assign in7142_2 = {c4328};
    Full_Adder FA_7142(s7142, c7142, in7142_1, in7142_2, c4326);
    wire[0:0] s7143, in7143_1, in7143_2;
    wire c7143;
    assign in7143_1 = {c4330};
    assign in7143_2 = {c4331};
    Full_Adder FA_7143(s7143, c7143, in7143_1, in7143_2, c4329);
    wire[0:0] s7144, in7144_1, in7144_2;
    wire c7144;
    assign in7144_1 = {c4333};
    assign in7144_2 = {c4334};
    Full_Adder FA_7144(s7144, c7144, in7144_1, in7144_2, c4332);
    wire[0:0] s7145, in7145_1, in7145_2;
    wire c7145;
    assign in7145_1 = {c4336};
    assign in7145_2 = {c4337};
    Full_Adder FA_7145(s7145, c7145, in7145_1, in7145_2, c4335);
    wire[0:0] s7146, in7146_1, in7146_2;
    wire c7146;
    assign in7146_1 = {c4339};
    assign in7146_2 = {c4340};
    Full_Adder FA_7146(s7146, c7146, in7146_1, in7146_2, c4338);
    wire[0:0] s7147, in7147_1, in7147_2;
    wire c7147;
    assign in7147_1 = {s4342[0]};
    assign in7147_2 = {s4343[0]};
    Full_Adder FA_7147(s7147, c7147, in7147_1, in7147_2, s4341[0]);
    wire[0:0] s7148, in7148_1, in7148_2;
    wire c7148;
    assign in7148_1 = {s4345[0]};
    assign in7148_2 = {s4346[0]};
    Full_Adder FA_7148(s7148, c7148, in7148_1, in7148_2, s4344[0]);
    wire[0:0] s7149, in7149_1, in7149_2;
    wire c7149;
    assign in7149_1 = {s4348[0]};
    assign in7149_2 = {s4349[0]};
    Full_Adder FA_7149(s7149, c7149, in7149_1, in7149_2, s4347[0]);
    wire[0:0] s7150, in7150_1, in7150_2;
    wire c7150;
    assign in7150_1 = {s4351[0]};
    assign in7150_2 = {s4352[0]};
    Full_Adder FA_7150(s7150, c7150, in7150_1, in7150_2, s4350[0]);
    wire[0:0] s7151, in7151_1, in7151_2;
    wire c7151;
    assign in7151_1 = {s4354[0]};
    assign in7151_2 = {s4355[0]};
    Full_Adder FA_7151(s7151, c7151, in7151_1, in7151_2, s4353[0]);
    wire[0:0] s7152, in7152_1, in7152_2;
    wire c7152;
    assign in7152_1 = {s4357[0]};
    assign in7152_2 = {s4358[0]};
    Full_Adder FA_7152(s7152, c7152, in7152_1, in7152_2, s4356[0]);
    wire[0:0] s7153, in7153_1, in7153_2;
    wire c7153;
    assign in7153_1 = {s4360[0]};
    assign in7153_2 = {s4361[0]};
    Full_Adder FA_7153(s7153, c7153, in7153_1, in7153_2, s4359[0]);
    wire[0:0] s7154, in7154_1, in7154_2;
    wire c7154;
    assign in7154_1 = {s4363[0]};
    assign in7154_2 = {s4364[0]};
    Full_Adder FA_7154(s7154, c7154, in7154_1, in7154_2, s4362[0]);
    wire[0:0] s7155, in7155_1, in7155_2;
    wire c7155;
    assign in7155_1 = {s4366[0]};
    assign in7155_2 = {s4367[0]};
    Full_Adder FA_7155(s7155, c7155, in7155_1, in7155_2, s4365[0]);
    wire[0:0] s7156, in7156_1, in7156_2;
    wire c7156;
    assign in7156_1 = {s1785[0]};
    assign in7156_2 = {c4341};
    Full_Adder FA_7156(s7156, c7156, in7156_1, in7156_2, s1784[0]);
    wire[0:0] s7157, in7157_1, in7157_2;
    wire c7157;
    assign in7157_1 = {c4343};
    assign in7157_2 = {c4344};
    Full_Adder FA_7157(s7157, c7157, in7157_1, in7157_2, c4342);
    wire[0:0] s7158, in7158_1, in7158_2;
    wire c7158;
    assign in7158_1 = {c4346};
    assign in7158_2 = {c4347};
    Full_Adder FA_7158(s7158, c7158, in7158_1, in7158_2, c4345);
    wire[0:0] s7159, in7159_1, in7159_2;
    wire c7159;
    assign in7159_1 = {c4349};
    assign in7159_2 = {c4350};
    Full_Adder FA_7159(s7159, c7159, in7159_1, in7159_2, c4348);
    wire[0:0] s7160, in7160_1, in7160_2;
    wire c7160;
    assign in7160_1 = {c4352};
    assign in7160_2 = {c4353};
    Full_Adder FA_7160(s7160, c7160, in7160_1, in7160_2, c4351);
    wire[0:0] s7161, in7161_1, in7161_2;
    wire c7161;
    assign in7161_1 = {c4355};
    assign in7161_2 = {c4356};
    Full_Adder FA_7161(s7161, c7161, in7161_1, in7161_2, c4354);
    wire[0:0] s7162, in7162_1, in7162_2;
    wire c7162;
    assign in7162_1 = {c4358};
    assign in7162_2 = {c4359};
    Full_Adder FA_7162(s7162, c7162, in7162_1, in7162_2, c4357);
    wire[0:0] s7163, in7163_1, in7163_2;
    wire c7163;
    assign in7163_1 = {c4361};
    assign in7163_2 = {c4362};
    Full_Adder FA_7163(s7163, c7163, in7163_1, in7163_2, c4360);
    wire[0:0] s7164, in7164_1, in7164_2;
    wire c7164;
    assign in7164_1 = {c4364};
    assign in7164_2 = {c4365};
    Full_Adder FA_7164(s7164, c7164, in7164_1, in7164_2, c4363);
    wire[0:0] s7165, in7165_1, in7165_2;
    wire c7165;
    assign in7165_1 = {c4367};
    assign in7165_2 = {c4368};
    Full_Adder FA_7165(s7165, c7165, in7165_1, in7165_2, c4366);
    wire[0:0] s7166, in7166_1, in7166_2;
    wire c7166;
    assign in7166_1 = {s4370[0]};
    assign in7166_2 = {s4371[0]};
    Full_Adder FA_7166(s7166, c7166, in7166_1, in7166_2, s4369[0]);
    wire[0:0] s7167, in7167_1, in7167_2;
    wire c7167;
    assign in7167_1 = {s4373[0]};
    assign in7167_2 = {s4374[0]};
    Full_Adder FA_7167(s7167, c7167, in7167_1, in7167_2, s4372[0]);
    wire[0:0] s7168, in7168_1, in7168_2;
    wire c7168;
    assign in7168_1 = {s4376[0]};
    assign in7168_2 = {s4377[0]};
    Full_Adder FA_7168(s7168, c7168, in7168_1, in7168_2, s4375[0]);
    wire[0:0] s7169, in7169_1, in7169_2;
    wire c7169;
    assign in7169_1 = {s4379[0]};
    assign in7169_2 = {s4380[0]};
    Full_Adder FA_7169(s7169, c7169, in7169_1, in7169_2, s4378[0]);
    wire[0:0] s7170, in7170_1, in7170_2;
    wire c7170;
    assign in7170_1 = {s4382[0]};
    assign in7170_2 = {s4383[0]};
    Full_Adder FA_7170(s7170, c7170, in7170_1, in7170_2, s4381[0]);
    wire[0:0] s7171, in7171_1, in7171_2;
    wire c7171;
    assign in7171_1 = {s4385[0]};
    assign in7171_2 = {s4386[0]};
    Full_Adder FA_7171(s7171, c7171, in7171_1, in7171_2, s4384[0]);
    wire[0:0] s7172, in7172_1, in7172_2;
    wire c7172;
    assign in7172_1 = {s4388[0]};
    assign in7172_2 = {s4389[0]};
    Full_Adder FA_7172(s7172, c7172, in7172_1, in7172_2, s4387[0]);
    wire[0:0] s7173, in7173_1, in7173_2;
    wire c7173;
    assign in7173_1 = {s4391[0]};
    assign in7173_2 = {s4392[0]};
    Full_Adder FA_7173(s7173, c7173, in7173_1, in7173_2, s4390[0]);
    wire[0:0] s7174, in7174_1, in7174_2;
    wire c7174;
    assign in7174_1 = {s4394[0]};
    assign in7174_2 = {s4395[0]};
    Full_Adder FA_7174(s7174, c7174, in7174_1, in7174_2, s4393[0]);
    wire[0:0] s7175, in7175_1, in7175_2;
    wire c7175;
    assign in7175_1 = {s1791[0]};
    assign in7175_2 = {c4369};
    Full_Adder FA_7175(s7175, c7175, in7175_1, in7175_2, s1790[0]);
    wire[0:0] s7176, in7176_1, in7176_2;
    wire c7176;
    assign in7176_1 = {c4371};
    assign in7176_2 = {c4372};
    Full_Adder FA_7176(s7176, c7176, in7176_1, in7176_2, c4370);
    wire[0:0] s7177, in7177_1, in7177_2;
    wire c7177;
    assign in7177_1 = {c4374};
    assign in7177_2 = {c4375};
    Full_Adder FA_7177(s7177, c7177, in7177_1, in7177_2, c4373);
    wire[0:0] s7178, in7178_1, in7178_2;
    wire c7178;
    assign in7178_1 = {c4377};
    assign in7178_2 = {c4378};
    Full_Adder FA_7178(s7178, c7178, in7178_1, in7178_2, c4376);
    wire[0:0] s7179, in7179_1, in7179_2;
    wire c7179;
    assign in7179_1 = {c4380};
    assign in7179_2 = {c4381};
    Full_Adder FA_7179(s7179, c7179, in7179_1, in7179_2, c4379);
    wire[0:0] s7180, in7180_1, in7180_2;
    wire c7180;
    assign in7180_1 = {c4383};
    assign in7180_2 = {c4384};
    Full_Adder FA_7180(s7180, c7180, in7180_1, in7180_2, c4382);
    wire[0:0] s7181, in7181_1, in7181_2;
    wire c7181;
    assign in7181_1 = {c4386};
    assign in7181_2 = {c4387};
    Full_Adder FA_7181(s7181, c7181, in7181_1, in7181_2, c4385);
    wire[0:0] s7182, in7182_1, in7182_2;
    wire c7182;
    assign in7182_1 = {c4389};
    assign in7182_2 = {c4390};
    Full_Adder FA_7182(s7182, c7182, in7182_1, in7182_2, c4388);
    wire[0:0] s7183, in7183_1, in7183_2;
    wire c7183;
    assign in7183_1 = {c4392};
    assign in7183_2 = {c4393};
    Full_Adder FA_7183(s7183, c7183, in7183_1, in7183_2, c4391);
    wire[0:0] s7184, in7184_1, in7184_2;
    wire c7184;
    assign in7184_1 = {c4395};
    assign in7184_2 = {c4396};
    Full_Adder FA_7184(s7184, c7184, in7184_1, in7184_2, c4394);
    wire[0:0] s7185, in7185_1, in7185_2;
    wire c7185;
    assign in7185_1 = {s4398[0]};
    assign in7185_2 = {s4399[0]};
    Full_Adder FA_7185(s7185, c7185, in7185_1, in7185_2, s4397[0]);
    wire[0:0] s7186, in7186_1, in7186_2;
    wire c7186;
    assign in7186_1 = {s4401[0]};
    assign in7186_2 = {s4402[0]};
    Full_Adder FA_7186(s7186, c7186, in7186_1, in7186_2, s4400[0]);
    wire[0:0] s7187, in7187_1, in7187_2;
    wire c7187;
    assign in7187_1 = {s4404[0]};
    assign in7187_2 = {s4405[0]};
    Full_Adder FA_7187(s7187, c7187, in7187_1, in7187_2, s4403[0]);
    wire[0:0] s7188, in7188_1, in7188_2;
    wire c7188;
    assign in7188_1 = {s4407[0]};
    assign in7188_2 = {s4408[0]};
    Full_Adder FA_7188(s7188, c7188, in7188_1, in7188_2, s4406[0]);
    wire[0:0] s7189, in7189_1, in7189_2;
    wire c7189;
    assign in7189_1 = {s4410[0]};
    assign in7189_2 = {s4411[0]};
    Full_Adder FA_7189(s7189, c7189, in7189_1, in7189_2, s4409[0]);
    wire[0:0] s7190, in7190_1, in7190_2;
    wire c7190;
    assign in7190_1 = {s4413[0]};
    assign in7190_2 = {s4414[0]};
    Full_Adder FA_7190(s7190, c7190, in7190_1, in7190_2, s4412[0]);
    wire[0:0] s7191, in7191_1, in7191_2;
    wire c7191;
    assign in7191_1 = {s4416[0]};
    assign in7191_2 = {s4417[0]};
    Full_Adder FA_7191(s7191, c7191, in7191_1, in7191_2, s4415[0]);
    wire[0:0] s7192, in7192_1, in7192_2;
    wire c7192;
    assign in7192_1 = {s4419[0]};
    assign in7192_2 = {s4420[0]};
    Full_Adder FA_7192(s7192, c7192, in7192_1, in7192_2, s4418[0]);
    wire[0:0] s7193, in7193_1, in7193_2;
    wire c7193;
    assign in7193_1 = {s4422[0]};
    assign in7193_2 = {s4423[0]};
    Full_Adder FA_7193(s7193, c7193, in7193_1, in7193_2, s4421[0]);
    wire[0:0] s7194, in7194_1, in7194_2;
    wire c7194;
    assign in7194_1 = {s1796[0]};
    assign in7194_2 = {c4397};
    Full_Adder FA_7194(s7194, c7194, in7194_1, in7194_2, s1795[0]);
    wire[0:0] s7195, in7195_1, in7195_2;
    wire c7195;
    assign in7195_1 = {c4399};
    assign in7195_2 = {c4400};
    Full_Adder FA_7195(s7195, c7195, in7195_1, in7195_2, c4398);
    wire[0:0] s7196, in7196_1, in7196_2;
    wire c7196;
    assign in7196_1 = {c4402};
    assign in7196_2 = {c4403};
    Full_Adder FA_7196(s7196, c7196, in7196_1, in7196_2, c4401);
    wire[0:0] s7197, in7197_1, in7197_2;
    wire c7197;
    assign in7197_1 = {c4405};
    assign in7197_2 = {c4406};
    Full_Adder FA_7197(s7197, c7197, in7197_1, in7197_2, c4404);
    wire[0:0] s7198, in7198_1, in7198_2;
    wire c7198;
    assign in7198_1 = {c4408};
    assign in7198_2 = {c4409};
    Full_Adder FA_7198(s7198, c7198, in7198_1, in7198_2, c4407);
    wire[0:0] s7199, in7199_1, in7199_2;
    wire c7199;
    assign in7199_1 = {c4411};
    assign in7199_2 = {c4412};
    Full_Adder FA_7199(s7199, c7199, in7199_1, in7199_2, c4410);
    wire[0:0] s7200, in7200_1, in7200_2;
    wire c7200;
    assign in7200_1 = {c4414};
    assign in7200_2 = {c4415};
    Full_Adder FA_7200(s7200, c7200, in7200_1, in7200_2, c4413);
    wire[0:0] s7201, in7201_1, in7201_2;
    wire c7201;
    assign in7201_1 = {c4417};
    assign in7201_2 = {c4418};
    Full_Adder FA_7201(s7201, c7201, in7201_1, in7201_2, c4416);
    wire[0:0] s7202, in7202_1, in7202_2;
    wire c7202;
    assign in7202_1 = {c4420};
    assign in7202_2 = {c4421};
    Full_Adder FA_7202(s7202, c7202, in7202_1, in7202_2, c4419);
    wire[0:0] s7203, in7203_1, in7203_2;
    wire c7203;
    assign in7203_1 = {c4423};
    assign in7203_2 = {c4424};
    Full_Adder FA_7203(s7203, c7203, in7203_1, in7203_2, c4422);
    wire[0:0] s7204, in7204_1, in7204_2;
    wire c7204;
    assign in7204_1 = {s4426[0]};
    assign in7204_2 = {s4427[0]};
    Full_Adder FA_7204(s7204, c7204, in7204_1, in7204_2, s4425[0]);
    wire[0:0] s7205, in7205_1, in7205_2;
    wire c7205;
    assign in7205_1 = {s4429[0]};
    assign in7205_2 = {s4430[0]};
    Full_Adder FA_7205(s7205, c7205, in7205_1, in7205_2, s4428[0]);
    wire[0:0] s7206, in7206_1, in7206_2;
    wire c7206;
    assign in7206_1 = {s4432[0]};
    assign in7206_2 = {s4433[0]};
    Full_Adder FA_7206(s7206, c7206, in7206_1, in7206_2, s4431[0]);
    wire[0:0] s7207, in7207_1, in7207_2;
    wire c7207;
    assign in7207_1 = {s4435[0]};
    assign in7207_2 = {s4436[0]};
    Full_Adder FA_7207(s7207, c7207, in7207_1, in7207_2, s4434[0]);
    wire[0:0] s7208, in7208_1, in7208_2;
    wire c7208;
    assign in7208_1 = {s4438[0]};
    assign in7208_2 = {s4439[0]};
    Full_Adder FA_7208(s7208, c7208, in7208_1, in7208_2, s4437[0]);
    wire[0:0] s7209, in7209_1, in7209_2;
    wire c7209;
    assign in7209_1 = {s4441[0]};
    assign in7209_2 = {s4442[0]};
    Full_Adder FA_7209(s7209, c7209, in7209_1, in7209_2, s4440[0]);
    wire[0:0] s7210, in7210_1, in7210_2;
    wire c7210;
    assign in7210_1 = {s4444[0]};
    assign in7210_2 = {s4445[0]};
    Full_Adder FA_7210(s7210, c7210, in7210_1, in7210_2, s4443[0]);
    wire[0:0] s7211, in7211_1, in7211_2;
    wire c7211;
    assign in7211_1 = {s4447[0]};
    assign in7211_2 = {s4448[0]};
    Full_Adder FA_7211(s7211, c7211, in7211_1, in7211_2, s4446[0]);
    wire[0:0] s7212, in7212_1, in7212_2;
    wire c7212;
    assign in7212_1 = {s4450[0]};
    assign in7212_2 = {s4451[0]};
    Full_Adder FA_7212(s7212, c7212, in7212_1, in7212_2, s4449[0]);
    wire[0:0] s7213, in7213_1, in7213_2;
    wire c7213;
    assign in7213_1 = {s1800[0]};
    assign in7213_2 = {c4425};
    Full_Adder FA_7213(s7213, c7213, in7213_1, in7213_2, s1799[0]);
    wire[0:0] s7214, in7214_1, in7214_2;
    wire c7214;
    assign in7214_1 = {c4427};
    assign in7214_2 = {c4428};
    Full_Adder FA_7214(s7214, c7214, in7214_1, in7214_2, c4426);
    wire[0:0] s7215, in7215_1, in7215_2;
    wire c7215;
    assign in7215_1 = {c4430};
    assign in7215_2 = {c4431};
    Full_Adder FA_7215(s7215, c7215, in7215_1, in7215_2, c4429);
    wire[0:0] s7216, in7216_1, in7216_2;
    wire c7216;
    assign in7216_1 = {c4433};
    assign in7216_2 = {c4434};
    Full_Adder FA_7216(s7216, c7216, in7216_1, in7216_2, c4432);
    wire[0:0] s7217, in7217_1, in7217_2;
    wire c7217;
    assign in7217_1 = {c4436};
    assign in7217_2 = {c4437};
    Full_Adder FA_7217(s7217, c7217, in7217_1, in7217_2, c4435);
    wire[0:0] s7218, in7218_1, in7218_2;
    wire c7218;
    assign in7218_1 = {c4439};
    assign in7218_2 = {c4440};
    Full_Adder FA_7218(s7218, c7218, in7218_1, in7218_2, c4438);
    wire[0:0] s7219, in7219_1, in7219_2;
    wire c7219;
    assign in7219_1 = {c4442};
    assign in7219_2 = {c4443};
    Full_Adder FA_7219(s7219, c7219, in7219_1, in7219_2, c4441);
    wire[0:0] s7220, in7220_1, in7220_2;
    wire c7220;
    assign in7220_1 = {c4445};
    assign in7220_2 = {c4446};
    Full_Adder FA_7220(s7220, c7220, in7220_1, in7220_2, c4444);
    wire[0:0] s7221, in7221_1, in7221_2;
    wire c7221;
    assign in7221_1 = {c4448};
    assign in7221_2 = {c4449};
    Full_Adder FA_7221(s7221, c7221, in7221_1, in7221_2, c4447);
    wire[0:0] s7222, in7222_1, in7222_2;
    wire c7222;
    assign in7222_1 = {c4451};
    assign in7222_2 = {c4452};
    Full_Adder FA_7222(s7222, c7222, in7222_1, in7222_2, c4450);
    wire[0:0] s7223, in7223_1, in7223_2;
    wire c7223;
    assign in7223_1 = {s4454[0]};
    assign in7223_2 = {s4455[0]};
    Full_Adder FA_7223(s7223, c7223, in7223_1, in7223_2, s4453[0]);
    wire[0:0] s7224, in7224_1, in7224_2;
    wire c7224;
    assign in7224_1 = {s4457[0]};
    assign in7224_2 = {s4458[0]};
    Full_Adder FA_7224(s7224, c7224, in7224_1, in7224_2, s4456[0]);
    wire[0:0] s7225, in7225_1, in7225_2;
    wire c7225;
    assign in7225_1 = {s4460[0]};
    assign in7225_2 = {s4461[0]};
    Full_Adder FA_7225(s7225, c7225, in7225_1, in7225_2, s4459[0]);
    wire[0:0] s7226, in7226_1, in7226_2;
    wire c7226;
    assign in7226_1 = {s4463[0]};
    assign in7226_2 = {s4464[0]};
    Full_Adder FA_7226(s7226, c7226, in7226_1, in7226_2, s4462[0]);
    wire[0:0] s7227, in7227_1, in7227_2;
    wire c7227;
    assign in7227_1 = {s4466[0]};
    assign in7227_2 = {s4467[0]};
    Full_Adder FA_7227(s7227, c7227, in7227_1, in7227_2, s4465[0]);
    wire[0:0] s7228, in7228_1, in7228_2;
    wire c7228;
    assign in7228_1 = {s4469[0]};
    assign in7228_2 = {s4470[0]};
    Full_Adder FA_7228(s7228, c7228, in7228_1, in7228_2, s4468[0]);
    wire[0:0] s7229, in7229_1, in7229_2;
    wire c7229;
    assign in7229_1 = {s4472[0]};
    assign in7229_2 = {s4473[0]};
    Full_Adder FA_7229(s7229, c7229, in7229_1, in7229_2, s4471[0]);
    wire[0:0] s7230, in7230_1, in7230_2;
    wire c7230;
    assign in7230_1 = {s4475[0]};
    assign in7230_2 = {s4476[0]};
    Full_Adder FA_7230(s7230, c7230, in7230_1, in7230_2, s4474[0]);
    wire[0:0] s7231, in7231_1, in7231_2;
    wire c7231;
    assign in7231_1 = {s4478[0]};
    assign in7231_2 = {s4479[0]};
    Full_Adder FA_7231(s7231, c7231, in7231_1, in7231_2, s4477[0]);
    wire[0:0] s7232, in7232_1, in7232_2;
    wire c7232;
    assign in7232_1 = {s1803[0]};
    assign in7232_2 = {c4453};
    Full_Adder FA_7232(s7232, c7232, in7232_1, in7232_2, s1802[0]);
    wire[0:0] s7233, in7233_1, in7233_2;
    wire c7233;
    assign in7233_1 = {c4455};
    assign in7233_2 = {c4456};
    Full_Adder FA_7233(s7233, c7233, in7233_1, in7233_2, c4454);
    wire[0:0] s7234, in7234_1, in7234_2;
    wire c7234;
    assign in7234_1 = {c4458};
    assign in7234_2 = {c4459};
    Full_Adder FA_7234(s7234, c7234, in7234_1, in7234_2, c4457);
    wire[0:0] s7235, in7235_1, in7235_2;
    wire c7235;
    assign in7235_1 = {c4461};
    assign in7235_2 = {c4462};
    Full_Adder FA_7235(s7235, c7235, in7235_1, in7235_2, c4460);
    wire[0:0] s7236, in7236_1, in7236_2;
    wire c7236;
    assign in7236_1 = {c4464};
    assign in7236_2 = {c4465};
    Full_Adder FA_7236(s7236, c7236, in7236_1, in7236_2, c4463);
    wire[0:0] s7237, in7237_1, in7237_2;
    wire c7237;
    assign in7237_1 = {c4467};
    assign in7237_2 = {c4468};
    Full_Adder FA_7237(s7237, c7237, in7237_1, in7237_2, c4466);
    wire[0:0] s7238, in7238_1, in7238_2;
    wire c7238;
    assign in7238_1 = {c4470};
    assign in7238_2 = {c4471};
    Full_Adder FA_7238(s7238, c7238, in7238_1, in7238_2, c4469);
    wire[0:0] s7239, in7239_1, in7239_2;
    wire c7239;
    assign in7239_1 = {c4473};
    assign in7239_2 = {c4474};
    Full_Adder FA_7239(s7239, c7239, in7239_1, in7239_2, c4472);
    wire[0:0] s7240, in7240_1, in7240_2;
    wire c7240;
    assign in7240_1 = {c4476};
    assign in7240_2 = {c4477};
    Full_Adder FA_7240(s7240, c7240, in7240_1, in7240_2, c4475);
    wire[0:0] s7241, in7241_1, in7241_2;
    wire c7241;
    assign in7241_1 = {c4479};
    assign in7241_2 = {c4480};
    Full_Adder FA_7241(s7241, c7241, in7241_1, in7241_2, c4478);
    wire[0:0] s7242, in7242_1, in7242_2;
    wire c7242;
    assign in7242_1 = {s4482[0]};
    assign in7242_2 = {s4483[0]};
    Full_Adder FA_7242(s7242, c7242, in7242_1, in7242_2, s4481[0]);
    wire[0:0] s7243, in7243_1, in7243_2;
    wire c7243;
    assign in7243_1 = {s4485[0]};
    assign in7243_2 = {s4486[0]};
    Full_Adder FA_7243(s7243, c7243, in7243_1, in7243_2, s4484[0]);
    wire[0:0] s7244, in7244_1, in7244_2;
    wire c7244;
    assign in7244_1 = {s4488[0]};
    assign in7244_2 = {s4489[0]};
    Full_Adder FA_7244(s7244, c7244, in7244_1, in7244_2, s4487[0]);
    wire[0:0] s7245, in7245_1, in7245_2;
    wire c7245;
    assign in7245_1 = {s4491[0]};
    assign in7245_2 = {s4492[0]};
    Full_Adder FA_7245(s7245, c7245, in7245_1, in7245_2, s4490[0]);
    wire[0:0] s7246, in7246_1, in7246_2;
    wire c7246;
    assign in7246_1 = {s4494[0]};
    assign in7246_2 = {s4495[0]};
    Full_Adder FA_7246(s7246, c7246, in7246_1, in7246_2, s4493[0]);
    wire[0:0] s7247, in7247_1, in7247_2;
    wire c7247;
    assign in7247_1 = {s4497[0]};
    assign in7247_2 = {s4498[0]};
    Full_Adder FA_7247(s7247, c7247, in7247_1, in7247_2, s4496[0]);
    wire[0:0] s7248, in7248_1, in7248_2;
    wire c7248;
    assign in7248_1 = {s4500[0]};
    assign in7248_2 = {s4501[0]};
    Full_Adder FA_7248(s7248, c7248, in7248_1, in7248_2, s4499[0]);
    wire[0:0] s7249, in7249_1, in7249_2;
    wire c7249;
    assign in7249_1 = {s4503[0]};
    assign in7249_2 = {s4504[0]};
    Full_Adder FA_7249(s7249, c7249, in7249_1, in7249_2, s4502[0]);
    wire[0:0] s7250, in7250_1, in7250_2;
    wire c7250;
    assign in7250_1 = {s4506[0]};
    assign in7250_2 = {s4507[0]};
    Full_Adder FA_7250(s7250, c7250, in7250_1, in7250_2, s4505[0]);
    wire[0:0] s7251, in7251_1, in7251_2;
    wire c7251;
    assign in7251_1 = {s1805[0]};
    assign in7251_2 = {c4481};
    Full_Adder FA_7251(s7251, c7251, in7251_1, in7251_2, s1804[0]);
    wire[0:0] s7252, in7252_1, in7252_2;
    wire c7252;
    assign in7252_1 = {c4483};
    assign in7252_2 = {c4484};
    Full_Adder FA_7252(s7252, c7252, in7252_1, in7252_2, c4482);
    wire[0:0] s7253, in7253_1, in7253_2;
    wire c7253;
    assign in7253_1 = {c4486};
    assign in7253_2 = {c4487};
    Full_Adder FA_7253(s7253, c7253, in7253_1, in7253_2, c4485);
    wire[0:0] s7254, in7254_1, in7254_2;
    wire c7254;
    assign in7254_1 = {c4489};
    assign in7254_2 = {c4490};
    Full_Adder FA_7254(s7254, c7254, in7254_1, in7254_2, c4488);
    wire[0:0] s7255, in7255_1, in7255_2;
    wire c7255;
    assign in7255_1 = {c4492};
    assign in7255_2 = {c4493};
    Full_Adder FA_7255(s7255, c7255, in7255_1, in7255_2, c4491);
    wire[0:0] s7256, in7256_1, in7256_2;
    wire c7256;
    assign in7256_1 = {c4495};
    assign in7256_2 = {c4496};
    Full_Adder FA_7256(s7256, c7256, in7256_1, in7256_2, c4494);
    wire[0:0] s7257, in7257_1, in7257_2;
    wire c7257;
    assign in7257_1 = {c4498};
    assign in7257_2 = {c4499};
    Full_Adder FA_7257(s7257, c7257, in7257_1, in7257_2, c4497);
    wire[0:0] s7258, in7258_1, in7258_2;
    wire c7258;
    assign in7258_1 = {c4501};
    assign in7258_2 = {c4502};
    Full_Adder FA_7258(s7258, c7258, in7258_1, in7258_2, c4500);
    wire[0:0] s7259, in7259_1, in7259_2;
    wire c7259;
    assign in7259_1 = {c4504};
    assign in7259_2 = {c4505};
    Full_Adder FA_7259(s7259, c7259, in7259_1, in7259_2, c4503);
    wire[0:0] s7260, in7260_1, in7260_2;
    wire c7260;
    assign in7260_1 = {c4507};
    assign in7260_2 = {c4508};
    Full_Adder FA_7260(s7260, c7260, in7260_1, in7260_2, c4506);
    wire[0:0] s7261, in7261_1, in7261_2;
    wire c7261;
    assign in7261_1 = {s4510[0]};
    assign in7261_2 = {s4511[0]};
    Full_Adder FA_7261(s7261, c7261, in7261_1, in7261_2, s4509[0]);
    wire[0:0] s7262, in7262_1, in7262_2;
    wire c7262;
    assign in7262_1 = {s4513[0]};
    assign in7262_2 = {s4514[0]};
    Full_Adder FA_7262(s7262, c7262, in7262_1, in7262_2, s4512[0]);
    wire[0:0] s7263, in7263_1, in7263_2;
    wire c7263;
    assign in7263_1 = {s4516[0]};
    assign in7263_2 = {s4517[0]};
    Full_Adder FA_7263(s7263, c7263, in7263_1, in7263_2, s4515[0]);
    wire[0:0] s7264, in7264_1, in7264_2;
    wire c7264;
    assign in7264_1 = {s4519[0]};
    assign in7264_2 = {s4520[0]};
    Full_Adder FA_7264(s7264, c7264, in7264_1, in7264_2, s4518[0]);
    wire[0:0] s7265, in7265_1, in7265_2;
    wire c7265;
    assign in7265_1 = {s4522[0]};
    assign in7265_2 = {s4523[0]};
    Full_Adder FA_7265(s7265, c7265, in7265_1, in7265_2, s4521[0]);
    wire[0:0] s7266, in7266_1, in7266_2;
    wire c7266;
    assign in7266_1 = {s4525[0]};
    assign in7266_2 = {s4526[0]};
    Full_Adder FA_7266(s7266, c7266, in7266_1, in7266_2, s4524[0]);
    wire[0:0] s7267, in7267_1, in7267_2;
    wire c7267;
    assign in7267_1 = {s4528[0]};
    assign in7267_2 = {s4529[0]};
    Full_Adder FA_7267(s7267, c7267, in7267_1, in7267_2, s4527[0]);
    wire[0:0] s7268, in7268_1, in7268_2;
    wire c7268;
    assign in7268_1 = {s4531[0]};
    assign in7268_2 = {s4532[0]};
    Full_Adder FA_7268(s7268, c7268, in7268_1, in7268_2, s4530[0]);
    wire[0:0] s7269, in7269_1, in7269_2;
    wire c7269;
    assign in7269_1 = {s4534[0]};
    assign in7269_2 = {s4535[0]};
    Full_Adder FA_7269(s7269, c7269, in7269_1, in7269_2, s4533[0]);
    wire[0:0] s7270, in7270_1, in7270_2;
    wire c7270;
    assign in7270_1 = {s1806[0]};
    assign in7270_2 = {c4509};
    Full_Adder FA_7270(s7270, c7270, in7270_1, in7270_2, c1805);
    wire[0:0] s7271, in7271_1, in7271_2;
    wire c7271;
    assign in7271_1 = {c4511};
    assign in7271_2 = {c4512};
    Full_Adder FA_7271(s7271, c7271, in7271_1, in7271_2, c4510);
    wire[0:0] s7272, in7272_1, in7272_2;
    wire c7272;
    assign in7272_1 = {c4514};
    assign in7272_2 = {c4515};
    Full_Adder FA_7272(s7272, c7272, in7272_1, in7272_2, c4513);
    wire[0:0] s7273, in7273_1, in7273_2;
    wire c7273;
    assign in7273_1 = {c4517};
    assign in7273_2 = {c4518};
    Full_Adder FA_7273(s7273, c7273, in7273_1, in7273_2, c4516);
    wire[0:0] s7274, in7274_1, in7274_2;
    wire c7274;
    assign in7274_1 = {c4520};
    assign in7274_2 = {c4521};
    Full_Adder FA_7274(s7274, c7274, in7274_1, in7274_2, c4519);
    wire[0:0] s7275, in7275_1, in7275_2;
    wire c7275;
    assign in7275_1 = {c4523};
    assign in7275_2 = {c4524};
    Full_Adder FA_7275(s7275, c7275, in7275_1, in7275_2, c4522);
    wire[0:0] s7276, in7276_1, in7276_2;
    wire c7276;
    assign in7276_1 = {c4526};
    assign in7276_2 = {c4527};
    Full_Adder FA_7276(s7276, c7276, in7276_1, in7276_2, c4525);
    wire[0:0] s7277, in7277_1, in7277_2;
    wire c7277;
    assign in7277_1 = {c4529};
    assign in7277_2 = {c4530};
    Full_Adder FA_7277(s7277, c7277, in7277_1, in7277_2, c4528);
    wire[0:0] s7278, in7278_1, in7278_2;
    wire c7278;
    assign in7278_1 = {c4532};
    assign in7278_2 = {c4533};
    Full_Adder FA_7278(s7278, c7278, in7278_1, in7278_2, c4531);
    wire[0:0] s7279, in7279_1, in7279_2;
    wire c7279;
    assign in7279_1 = {c4535};
    assign in7279_2 = {c4536};
    Full_Adder FA_7279(s7279, c7279, in7279_1, in7279_2, c4534);
    wire[0:0] s7280, in7280_1, in7280_2;
    wire c7280;
    assign in7280_1 = {s4538[0]};
    assign in7280_2 = {s4539[0]};
    Full_Adder FA_7280(s7280, c7280, in7280_1, in7280_2, s4537[0]);
    wire[0:0] s7281, in7281_1, in7281_2;
    wire c7281;
    assign in7281_1 = {s4541[0]};
    assign in7281_2 = {s4542[0]};
    Full_Adder FA_7281(s7281, c7281, in7281_1, in7281_2, s4540[0]);
    wire[0:0] s7282, in7282_1, in7282_2;
    wire c7282;
    assign in7282_1 = {s4544[0]};
    assign in7282_2 = {s4545[0]};
    Full_Adder FA_7282(s7282, c7282, in7282_1, in7282_2, s4543[0]);
    wire[0:0] s7283, in7283_1, in7283_2;
    wire c7283;
    assign in7283_1 = {s4547[0]};
    assign in7283_2 = {s4548[0]};
    Full_Adder FA_7283(s7283, c7283, in7283_1, in7283_2, s4546[0]);
    wire[0:0] s7284, in7284_1, in7284_2;
    wire c7284;
    assign in7284_1 = {s4550[0]};
    assign in7284_2 = {s4551[0]};
    Full_Adder FA_7284(s7284, c7284, in7284_1, in7284_2, s4549[0]);
    wire[0:0] s7285, in7285_1, in7285_2;
    wire c7285;
    assign in7285_1 = {s4553[0]};
    assign in7285_2 = {s4554[0]};
    Full_Adder FA_7285(s7285, c7285, in7285_1, in7285_2, s4552[0]);
    wire[0:0] s7286, in7286_1, in7286_2;
    wire c7286;
    assign in7286_1 = {s4556[0]};
    assign in7286_2 = {s4557[0]};
    Full_Adder FA_7286(s7286, c7286, in7286_1, in7286_2, s4555[0]);
    wire[0:0] s7287, in7287_1, in7287_2;
    wire c7287;
    assign in7287_1 = {s4559[0]};
    assign in7287_2 = {s4560[0]};
    Full_Adder FA_7287(s7287, c7287, in7287_1, in7287_2, s4558[0]);
    wire[0:0] s7288, in7288_1, in7288_2;
    wire c7288;
    assign in7288_1 = {s4562[0]};
    assign in7288_2 = {s4563[0]};
    Full_Adder FA_7288(s7288, c7288, in7288_1, in7288_2, s4561[0]);
    wire[0:0] s7289, in7289_1, in7289_2;
    wire c7289;
    assign in7289_1 = {c1806};
    assign in7289_2 = {c4537};
    Full_Adder FA_7289(s7289, c7289, in7289_1, in7289_2, pp127[43]);
    wire[0:0] s7290, in7290_1, in7290_2;
    wire c7290;
    assign in7290_1 = {c4539};
    assign in7290_2 = {c4540};
    Full_Adder FA_7290(s7290, c7290, in7290_1, in7290_2, c4538);
    wire[0:0] s7291, in7291_1, in7291_2;
    wire c7291;
    assign in7291_1 = {c4542};
    assign in7291_2 = {c4543};
    Full_Adder FA_7291(s7291, c7291, in7291_1, in7291_2, c4541);
    wire[0:0] s7292, in7292_1, in7292_2;
    wire c7292;
    assign in7292_1 = {c4545};
    assign in7292_2 = {c4546};
    Full_Adder FA_7292(s7292, c7292, in7292_1, in7292_2, c4544);
    wire[0:0] s7293, in7293_1, in7293_2;
    wire c7293;
    assign in7293_1 = {c4548};
    assign in7293_2 = {c4549};
    Full_Adder FA_7293(s7293, c7293, in7293_1, in7293_2, c4547);
    wire[0:0] s7294, in7294_1, in7294_2;
    wire c7294;
    assign in7294_1 = {c4551};
    assign in7294_2 = {c4552};
    Full_Adder FA_7294(s7294, c7294, in7294_1, in7294_2, c4550);
    wire[0:0] s7295, in7295_1, in7295_2;
    wire c7295;
    assign in7295_1 = {c4554};
    assign in7295_2 = {c4555};
    Full_Adder FA_7295(s7295, c7295, in7295_1, in7295_2, c4553);
    wire[0:0] s7296, in7296_1, in7296_2;
    wire c7296;
    assign in7296_1 = {c4557};
    assign in7296_2 = {c4558};
    Full_Adder FA_7296(s7296, c7296, in7296_1, in7296_2, c4556);
    wire[0:0] s7297, in7297_1, in7297_2;
    wire c7297;
    assign in7297_1 = {c4560};
    assign in7297_2 = {c4561};
    Full_Adder FA_7297(s7297, c7297, in7297_1, in7297_2, c4559);
    wire[0:0] s7298, in7298_1, in7298_2;
    wire c7298;
    assign in7298_1 = {c4563};
    assign in7298_2 = {c4564};
    Full_Adder FA_7298(s7298, c7298, in7298_1, in7298_2, c4562);
    wire[0:0] s7299, in7299_1, in7299_2;
    wire c7299;
    assign in7299_1 = {s4566[0]};
    assign in7299_2 = {s4567[0]};
    Full_Adder FA_7299(s7299, c7299, in7299_1, in7299_2, s4565[0]);
    wire[0:0] s7300, in7300_1, in7300_2;
    wire c7300;
    assign in7300_1 = {s4569[0]};
    assign in7300_2 = {s4570[0]};
    Full_Adder FA_7300(s7300, c7300, in7300_1, in7300_2, s4568[0]);
    wire[0:0] s7301, in7301_1, in7301_2;
    wire c7301;
    assign in7301_1 = {s4572[0]};
    assign in7301_2 = {s4573[0]};
    Full_Adder FA_7301(s7301, c7301, in7301_1, in7301_2, s4571[0]);
    wire[0:0] s7302, in7302_1, in7302_2;
    wire c7302;
    assign in7302_1 = {s4575[0]};
    assign in7302_2 = {s4576[0]};
    Full_Adder FA_7302(s7302, c7302, in7302_1, in7302_2, s4574[0]);
    wire[0:0] s7303, in7303_1, in7303_2;
    wire c7303;
    assign in7303_1 = {s4578[0]};
    assign in7303_2 = {s4579[0]};
    Full_Adder FA_7303(s7303, c7303, in7303_1, in7303_2, s4577[0]);
    wire[0:0] s7304, in7304_1, in7304_2;
    wire c7304;
    assign in7304_1 = {s4581[0]};
    assign in7304_2 = {s4582[0]};
    Full_Adder FA_7304(s7304, c7304, in7304_1, in7304_2, s4580[0]);
    wire[0:0] s7305, in7305_1, in7305_2;
    wire c7305;
    assign in7305_1 = {s4584[0]};
    assign in7305_2 = {s4585[0]};
    Full_Adder FA_7305(s7305, c7305, in7305_1, in7305_2, s4583[0]);
    wire[0:0] s7306, in7306_1, in7306_2;
    wire c7306;
    assign in7306_1 = {s4587[0]};
    assign in7306_2 = {s4588[0]};
    Full_Adder FA_7306(s7306, c7306, in7306_1, in7306_2, s4586[0]);
    wire[0:0] s7307, in7307_1, in7307_2;
    wire c7307;
    assign in7307_1 = {s4590[0]};
    assign in7307_2 = {s4591[0]};
    Full_Adder FA_7307(s7307, c7307, in7307_1, in7307_2, s4589[0]);
    wire[0:0] s7308, in7308_1, in7308_2;
    wire c7308;
    assign in7308_1 = {pp126[45]};
    assign in7308_2 = {pp127[44]};
    Full_Adder FA_7308(s7308, c7308, in7308_1, in7308_2, pp125[46]);
    wire[0:0] s7309, in7309_1, in7309_2;
    wire c7309;
    assign in7309_1 = {c4566};
    assign in7309_2 = {c4567};
    Full_Adder FA_7309(s7309, c7309, in7309_1, in7309_2, c4565);
    wire[0:0] s7310, in7310_1, in7310_2;
    wire c7310;
    assign in7310_1 = {c4569};
    assign in7310_2 = {c4570};
    Full_Adder FA_7310(s7310, c7310, in7310_1, in7310_2, c4568);
    wire[0:0] s7311, in7311_1, in7311_2;
    wire c7311;
    assign in7311_1 = {c4572};
    assign in7311_2 = {c4573};
    Full_Adder FA_7311(s7311, c7311, in7311_1, in7311_2, c4571);
    wire[0:0] s7312, in7312_1, in7312_2;
    wire c7312;
    assign in7312_1 = {c4575};
    assign in7312_2 = {c4576};
    Full_Adder FA_7312(s7312, c7312, in7312_1, in7312_2, c4574);
    wire[0:0] s7313, in7313_1, in7313_2;
    wire c7313;
    assign in7313_1 = {c4578};
    assign in7313_2 = {c4579};
    Full_Adder FA_7313(s7313, c7313, in7313_1, in7313_2, c4577);
    wire[0:0] s7314, in7314_1, in7314_2;
    wire c7314;
    assign in7314_1 = {c4581};
    assign in7314_2 = {c4582};
    Full_Adder FA_7314(s7314, c7314, in7314_1, in7314_2, c4580);
    wire[0:0] s7315, in7315_1, in7315_2;
    wire c7315;
    assign in7315_1 = {c4584};
    assign in7315_2 = {c4585};
    Full_Adder FA_7315(s7315, c7315, in7315_1, in7315_2, c4583);
    wire[0:0] s7316, in7316_1, in7316_2;
    wire c7316;
    assign in7316_1 = {c4587};
    assign in7316_2 = {c4588};
    Full_Adder FA_7316(s7316, c7316, in7316_1, in7316_2, c4586);
    wire[0:0] s7317, in7317_1, in7317_2;
    wire c7317;
    assign in7317_1 = {c4590};
    assign in7317_2 = {c4591};
    Full_Adder FA_7317(s7317, c7317, in7317_1, in7317_2, c4589);
    wire[0:0] s7318, in7318_1, in7318_2;
    wire c7318;
    assign in7318_1 = {s4593[0]};
    assign in7318_2 = {s4594[0]};
    Full_Adder FA_7318(s7318, c7318, in7318_1, in7318_2, c4592);
    wire[0:0] s7319, in7319_1, in7319_2;
    wire c7319;
    assign in7319_1 = {s4596[0]};
    assign in7319_2 = {s4597[0]};
    Full_Adder FA_7319(s7319, c7319, in7319_1, in7319_2, s4595[0]);
    wire[0:0] s7320, in7320_1, in7320_2;
    wire c7320;
    assign in7320_1 = {s4599[0]};
    assign in7320_2 = {s4600[0]};
    Full_Adder FA_7320(s7320, c7320, in7320_1, in7320_2, s4598[0]);
    wire[0:0] s7321, in7321_1, in7321_2;
    wire c7321;
    assign in7321_1 = {s4602[0]};
    assign in7321_2 = {s4603[0]};
    Full_Adder FA_7321(s7321, c7321, in7321_1, in7321_2, s4601[0]);
    wire[0:0] s7322, in7322_1, in7322_2;
    wire c7322;
    assign in7322_1 = {s4605[0]};
    assign in7322_2 = {s4606[0]};
    Full_Adder FA_7322(s7322, c7322, in7322_1, in7322_2, s4604[0]);
    wire[0:0] s7323, in7323_1, in7323_2;
    wire c7323;
    assign in7323_1 = {s4608[0]};
    assign in7323_2 = {s4609[0]};
    Full_Adder FA_7323(s7323, c7323, in7323_1, in7323_2, s4607[0]);
    wire[0:0] s7324, in7324_1, in7324_2;
    wire c7324;
    assign in7324_1 = {s4611[0]};
    assign in7324_2 = {s4612[0]};
    Full_Adder FA_7324(s7324, c7324, in7324_1, in7324_2, s4610[0]);
    wire[0:0] s7325, in7325_1, in7325_2;
    wire c7325;
    assign in7325_1 = {s4614[0]};
    assign in7325_2 = {s4615[0]};
    Full_Adder FA_7325(s7325, c7325, in7325_1, in7325_2, s4613[0]);
    wire[0:0] s7326, in7326_1, in7326_2;
    wire c7326;
    assign in7326_1 = {s4617[0]};
    assign in7326_2 = {s4618[0]};
    Full_Adder FA_7326(s7326, c7326, in7326_1, in7326_2, s4616[0]);
    wire[0:0] s7327, in7327_1, in7327_2;
    wire c7327;
    assign in7327_1 = {pp124[48]};
    assign in7327_2 = {pp125[47]};
    Full_Adder FA_7327(s7327, c7327, in7327_1, in7327_2, pp123[49]);
    wire[0:0] s7328, in7328_1, in7328_2;
    wire c7328;
    assign in7328_1 = {pp127[45]};
    assign in7328_2 = {c4593};
    Full_Adder FA_7328(s7328, c7328, in7328_1, in7328_2, pp126[46]);
    wire[0:0] s7329, in7329_1, in7329_2;
    wire c7329;
    assign in7329_1 = {c4595};
    assign in7329_2 = {c4596};
    Full_Adder FA_7329(s7329, c7329, in7329_1, in7329_2, c4594);
    wire[0:0] s7330, in7330_1, in7330_2;
    wire c7330;
    assign in7330_1 = {c4598};
    assign in7330_2 = {c4599};
    Full_Adder FA_7330(s7330, c7330, in7330_1, in7330_2, c4597);
    wire[0:0] s7331, in7331_1, in7331_2;
    wire c7331;
    assign in7331_1 = {c4601};
    assign in7331_2 = {c4602};
    Full_Adder FA_7331(s7331, c7331, in7331_1, in7331_2, c4600);
    wire[0:0] s7332, in7332_1, in7332_2;
    wire c7332;
    assign in7332_1 = {c4604};
    assign in7332_2 = {c4605};
    Full_Adder FA_7332(s7332, c7332, in7332_1, in7332_2, c4603);
    wire[0:0] s7333, in7333_1, in7333_2;
    wire c7333;
    assign in7333_1 = {c4607};
    assign in7333_2 = {c4608};
    Full_Adder FA_7333(s7333, c7333, in7333_1, in7333_2, c4606);
    wire[0:0] s7334, in7334_1, in7334_2;
    wire c7334;
    assign in7334_1 = {c4610};
    assign in7334_2 = {c4611};
    Full_Adder FA_7334(s7334, c7334, in7334_1, in7334_2, c4609);
    wire[0:0] s7335, in7335_1, in7335_2;
    wire c7335;
    assign in7335_1 = {c4613};
    assign in7335_2 = {c4614};
    Full_Adder FA_7335(s7335, c7335, in7335_1, in7335_2, c4612);
    wire[0:0] s7336, in7336_1, in7336_2;
    wire c7336;
    assign in7336_1 = {c4616};
    assign in7336_2 = {c4617};
    Full_Adder FA_7336(s7336, c7336, in7336_1, in7336_2, c4615);
    wire[0:0] s7337, in7337_1, in7337_2;
    wire c7337;
    assign in7337_1 = {c4619};
    assign in7337_2 = {s4620[0]};
    Full_Adder FA_7337(s7337, c7337, in7337_1, in7337_2, c4618);
    wire[0:0] s7338, in7338_1, in7338_2;
    wire c7338;
    assign in7338_1 = {s4622[0]};
    assign in7338_2 = {s4623[0]};
    Full_Adder FA_7338(s7338, c7338, in7338_1, in7338_2, s4621[0]);
    wire[0:0] s7339, in7339_1, in7339_2;
    wire c7339;
    assign in7339_1 = {s4625[0]};
    assign in7339_2 = {s4626[0]};
    Full_Adder FA_7339(s7339, c7339, in7339_1, in7339_2, s4624[0]);
    wire[0:0] s7340, in7340_1, in7340_2;
    wire c7340;
    assign in7340_1 = {s4628[0]};
    assign in7340_2 = {s4629[0]};
    Full_Adder FA_7340(s7340, c7340, in7340_1, in7340_2, s4627[0]);
    wire[0:0] s7341, in7341_1, in7341_2;
    wire c7341;
    assign in7341_1 = {s4631[0]};
    assign in7341_2 = {s4632[0]};
    Full_Adder FA_7341(s7341, c7341, in7341_1, in7341_2, s4630[0]);
    wire[0:0] s7342, in7342_1, in7342_2;
    wire c7342;
    assign in7342_1 = {s4634[0]};
    assign in7342_2 = {s4635[0]};
    Full_Adder FA_7342(s7342, c7342, in7342_1, in7342_2, s4633[0]);
    wire[0:0] s7343, in7343_1, in7343_2;
    wire c7343;
    assign in7343_1 = {s4637[0]};
    assign in7343_2 = {s4638[0]};
    Full_Adder FA_7343(s7343, c7343, in7343_1, in7343_2, s4636[0]);
    wire[0:0] s7344, in7344_1, in7344_2;
    wire c7344;
    assign in7344_1 = {s4640[0]};
    assign in7344_2 = {s4641[0]};
    Full_Adder FA_7344(s7344, c7344, in7344_1, in7344_2, s4639[0]);
    wire[0:0] s7345, in7345_1, in7345_2;
    wire c7345;
    assign in7345_1 = {s4643[0]};
    assign in7345_2 = {s4644[0]};
    Full_Adder FA_7345(s7345, c7345, in7345_1, in7345_2, s4642[0]);
    wire[0:0] s7346, in7346_1, in7346_2;
    wire c7346;
    assign in7346_1 = {pp122[51]};
    assign in7346_2 = {pp123[50]};
    Full_Adder FA_7346(s7346, c7346, in7346_1, in7346_2, pp121[52]);
    wire[0:0] s7347, in7347_1, in7347_2;
    wire c7347;
    assign in7347_1 = {pp125[48]};
    assign in7347_2 = {pp126[47]};
    Full_Adder FA_7347(s7347, c7347, in7347_1, in7347_2, pp124[49]);
    wire[0:0] s7348, in7348_1, in7348_2;
    wire c7348;
    assign in7348_1 = {c4620};
    assign in7348_2 = {c4621};
    Full_Adder FA_7348(s7348, c7348, in7348_1, in7348_2, pp127[46]);
    wire[0:0] s7349, in7349_1, in7349_2;
    wire c7349;
    assign in7349_1 = {c4623};
    assign in7349_2 = {c4624};
    Full_Adder FA_7349(s7349, c7349, in7349_1, in7349_2, c4622);
    wire[0:0] s7350, in7350_1, in7350_2;
    wire c7350;
    assign in7350_1 = {c4626};
    assign in7350_2 = {c4627};
    Full_Adder FA_7350(s7350, c7350, in7350_1, in7350_2, c4625);
    wire[0:0] s7351, in7351_1, in7351_2;
    wire c7351;
    assign in7351_1 = {c4629};
    assign in7351_2 = {c4630};
    Full_Adder FA_7351(s7351, c7351, in7351_1, in7351_2, c4628);
    wire[0:0] s7352, in7352_1, in7352_2;
    wire c7352;
    assign in7352_1 = {c4632};
    assign in7352_2 = {c4633};
    Full_Adder FA_7352(s7352, c7352, in7352_1, in7352_2, c4631);
    wire[0:0] s7353, in7353_1, in7353_2;
    wire c7353;
    assign in7353_1 = {c4635};
    assign in7353_2 = {c4636};
    Full_Adder FA_7353(s7353, c7353, in7353_1, in7353_2, c4634);
    wire[0:0] s7354, in7354_1, in7354_2;
    wire c7354;
    assign in7354_1 = {c4638};
    assign in7354_2 = {c4639};
    Full_Adder FA_7354(s7354, c7354, in7354_1, in7354_2, c4637);
    wire[0:0] s7355, in7355_1, in7355_2;
    wire c7355;
    assign in7355_1 = {c4641};
    assign in7355_2 = {c4642};
    Full_Adder FA_7355(s7355, c7355, in7355_1, in7355_2, c4640);
    wire[0:0] s7356, in7356_1, in7356_2;
    wire c7356;
    assign in7356_1 = {c4644};
    assign in7356_2 = {c4645};
    Full_Adder FA_7356(s7356, c7356, in7356_1, in7356_2, c4643);
    wire[0:0] s7357, in7357_1, in7357_2;
    wire c7357;
    assign in7357_1 = {s4647[0]};
    assign in7357_2 = {s4648[0]};
    Full_Adder FA_7357(s7357, c7357, in7357_1, in7357_2, s4646[0]);
    wire[0:0] s7358, in7358_1, in7358_2;
    wire c7358;
    assign in7358_1 = {s4650[0]};
    assign in7358_2 = {s4651[0]};
    Full_Adder FA_7358(s7358, c7358, in7358_1, in7358_2, s4649[0]);
    wire[0:0] s7359, in7359_1, in7359_2;
    wire c7359;
    assign in7359_1 = {s4653[0]};
    assign in7359_2 = {s4654[0]};
    Full_Adder FA_7359(s7359, c7359, in7359_1, in7359_2, s4652[0]);
    wire[0:0] s7360, in7360_1, in7360_2;
    wire c7360;
    assign in7360_1 = {s4656[0]};
    assign in7360_2 = {s4657[0]};
    Full_Adder FA_7360(s7360, c7360, in7360_1, in7360_2, s4655[0]);
    wire[0:0] s7361, in7361_1, in7361_2;
    wire c7361;
    assign in7361_1 = {s4659[0]};
    assign in7361_2 = {s4660[0]};
    Full_Adder FA_7361(s7361, c7361, in7361_1, in7361_2, s4658[0]);
    wire[0:0] s7362, in7362_1, in7362_2;
    wire c7362;
    assign in7362_1 = {s4662[0]};
    assign in7362_2 = {s4663[0]};
    Full_Adder FA_7362(s7362, c7362, in7362_1, in7362_2, s4661[0]);
    wire[0:0] s7363, in7363_1, in7363_2;
    wire c7363;
    assign in7363_1 = {s4665[0]};
    assign in7363_2 = {s4666[0]};
    Full_Adder FA_7363(s7363, c7363, in7363_1, in7363_2, s4664[0]);
    wire[0:0] s7364, in7364_1, in7364_2;
    wire c7364;
    assign in7364_1 = {s4668[0]};
    assign in7364_2 = {s4669[0]};
    Full_Adder FA_7364(s7364, c7364, in7364_1, in7364_2, s4667[0]);
    wire[0:0] s7365, in7365_1, in7365_2;
    wire c7365;
    assign in7365_1 = {pp120[54]};
    assign in7365_2 = {pp121[53]};
    Full_Adder FA_7365(s7365, c7365, in7365_1, in7365_2, pp119[55]);
    wire[0:0] s7366, in7366_1, in7366_2;
    wire c7366;
    assign in7366_1 = {pp123[51]};
    assign in7366_2 = {pp124[50]};
    Full_Adder FA_7366(s7366, c7366, in7366_1, in7366_2, pp122[52]);
    wire[0:0] s7367, in7367_1, in7367_2;
    wire c7367;
    assign in7367_1 = {pp126[48]};
    assign in7367_2 = {pp127[47]};
    Full_Adder FA_7367(s7367, c7367, in7367_1, in7367_2, pp125[49]);
    wire[0:0] s7368, in7368_1, in7368_2;
    wire c7368;
    assign in7368_1 = {c4647};
    assign in7368_2 = {c4648};
    Full_Adder FA_7368(s7368, c7368, in7368_1, in7368_2, c4646);
    wire[0:0] s7369, in7369_1, in7369_2;
    wire c7369;
    assign in7369_1 = {c4650};
    assign in7369_2 = {c4651};
    Full_Adder FA_7369(s7369, c7369, in7369_1, in7369_2, c4649);
    wire[0:0] s7370, in7370_1, in7370_2;
    wire c7370;
    assign in7370_1 = {c4653};
    assign in7370_2 = {c4654};
    Full_Adder FA_7370(s7370, c7370, in7370_1, in7370_2, c4652);
    wire[0:0] s7371, in7371_1, in7371_2;
    wire c7371;
    assign in7371_1 = {c4656};
    assign in7371_2 = {c4657};
    Full_Adder FA_7371(s7371, c7371, in7371_1, in7371_2, c4655);
    wire[0:0] s7372, in7372_1, in7372_2;
    wire c7372;
    assign in7372_1 = {c4659};
    assign in7372_2 = {c4660};
    Full_Adder FA_7372(s7372, c7372, in7372_1, in7372_2, c4658);
    wire[0:0] s7373, in7373_1, in7373_2;
    wire c7373;
    assign in7373_1 = {c4662};
    assign in7373_2 = {c4663};
    Full_Adder FA_7373(s7373, c7373, in7373_1, in7373_2, c4661);
    wire[0:0] s7374, in7374_1, in7374_2;
    wire c7374;
    assign in7374_1 = {c4665};
    assign in7374_2 = {c4666};
    Full_Adder FA_7374(s7374, c7374, in7374_1, in7374_2, c4664);
    wire[0:0] s7375, in7375_1, in7375_2;
    wire c7375;
    assign in7375_1 = {c4668};
    assign in7375_2 = {c4669};
    Full_Adder FA_7375(s7375, c7375, in7375_1, in7375_2, c4667);
    wire[0:0] s7376, in7376_1, in7376_2;
    wire c7376;
    assign in7376_1 = {s4671[0]};
    assign in7376_2 = {s4672[0]};
    Full_Adder FA_7376(s7376, c7376, in7376_1, in7376_2, c4670);
    wire[0:0] s7377, in7377_1, in7377_2;
    wire c7377;
    assign in7377_1 = {s4674[0]};
    assign in7377_2 = {s4675[0]};
    Full_Adder FA_7377(s7377, c7377, in7377_1, in7377_2, s4673[0]);
    wire[0:0] s7378, in7378_1, in7378_2;
    wire c7378;
    assign in7378_1 = {s4677[0]};
    assign in7378_2 = {s4678[0]};
    Full_Adder FA_7378(s7378, c7378, in7378_1, in7378_2, s4676[0]);
    wire[0:0] s7379, in7379_1, in7379_2;
    wire c7379;
    assign in7379_1 = {s4680[0]};
    assign in7379_2 = {s4681[0]};
    Full_Adder FA_7379(s7379, c7379, in7379_1, in7379_2, s4679[0]);
    wire[0:0] s7380, in7380_1, in7380_2;
    wire c7380;
    assign in7380_1 = {s4683[0]};
    assign in7380_2 = {s4684[0]};
    Full_Adder FA_7380(s7380, c7380, in7380_1, in7380_2, s4682[0]);
    wire[0:0] s7381, in7381_1, in7381_2;
    wire c7381;
    assign in7381_1 = {s4686[0]};
    assign in7381_2 = {s4687[0]};
    Full_Adder FA_7381(s7381, c7381, in7381_1, in7381_2, s4685[0]);
    wire[0:0] s7382, in7382_1, in7382_2;
    wire c7382;
    assign in7382_1 = {s4689[0]};
    assign in7382_2 = {s4690[0]};
    Full_Adder FA_7382(s7382, c7382, in7382_1, in7382_2, s4688[0]);
    wire[0:0] s7383, in7383_1, in7383_2;
    wire c7383;
    assign in7383_1 = {s4692[0]};
    assign in7383_2 = {s4693[0]};
    Full_Adder FA_7383(s7383, c7383, in7383_1, in7383_2, s4691[0]);
    wire[0:0] s7384, in7384_1, in7384_2;
    wire c7384;
    assign in7384_1 = {pp118[57]};
    assign in7384_2 = {pp119[56]};
    Full_Adder FA_7384(s7384, c7384, in7384_1, in7384_2, pp117[58]);
    wire[0:0] s7385, in7385_1, in7385_2;
    wire c7385;
    assign in7385_1 = {pp121[54]};
    assign in7385_2 = {pp122[53]};
    Full_Adder FA_7385(s7385, c7385, in7385_1, in7385_2, pp120[55]);
    wire[0:0] s7386, in7386_1, in7386_2;
    wire c7386;
    assign in7386_1 = {pp124[51]};
    assign in7386_2 = {pp125[50]};
    Full_Adder FA_7386(s7386, c7386, in7386_1, in7386_2, pp123[52]);
    wire[0:0] s7387, in7387_1, in7387_2;
    wire c7387;
    assign in7387_1 = {pp127[48]};
    assign in7387_2 = {c4671};
    Full_Adder FA_7387(s7387, c7387, in7387_1, in7387_2, pp126[49]);
    wire[0:0] s7388, in7388_1, in7388_2;
    wire c7388;
    assign in7388_1 = {c4673};
    assign in7388_2 = {c4674};
    Full_Adder FA_7388(s7388, c7388, in7388_1, in7388_2, c4672);
    wire[0:0] s7389, in7389_1, in7389_2;
    wire c7389;
    assign in7389_1 = {c4676};
    assign in7389_2 = {c4677};
    Full_Adder FA_7389(s7389, c7389, in7389_1, in7389_2, c4675);
    wire[0:0] s7390, in7390_1, in7390_2;
    wire c7390;
    assign in7390_1 = {c4679};
    assign in7390_2 = {c4680};
    Full_Adder FA_7390(s7390, c7390, in7390_1, in7390_2, c4678);
    wire[0:0] s7391, in7391_1, in7391_2;
    wire c7391;
    assign in7391_1 = {c4682};
    assign in7391_2 = {c4683};
    Full_Adder FA_7391(s7391, c7391, in7391_1, in7391_2, c4681);
    wire[0:0] s7392, in7392_1, in7392_2;
    wire c7392;
    assign in7392_1 = {c4685};
    assign in7392_2 = {c4686};
    Full_Adder FA_7392(s7392, c7392, in7392_1, in7392_2, c4684);
    wire[0:0] s7393, in7393_1, in7393_2;
    wire c7393;
    assign in7393_1 = {c4688};
    assign in7393_2 = {c4689};
    Full_Adder FA_7393(s7393, c7393, in7393_1, in7393_2, c4687);
    wire[0:0] s7394, in7394_1, in7394_2;
    wire c7394;
    assign in7394_1 = {c4691};
    assign in7394_2 = {c4692};
    Full_Adder FA_7394(s7394, c7394, in7394_1, in7394_2, c4690);
    wire[0:0] s7395, in7395_1, in7395_2;
    wire c7395;
    assign in7395_1 = {c4694};
    assign in7395_2 = {s4695[0]};
    Full_Adder FA_7395(s7395, c7395, in7395_1, in7395_2, c4693);
    wire[0:0] s7396, in7396_1, in7396_2;
    wire c7396;
    assign in7396_1 = {s4697[0]};
    assign in7396_2 = {s4698[0]};
    Full_Adder FA_7396(s7396, c7396, in7396_1, in7396_2, s4696[0]);
    wire[0:0] s7397, in7397_1, in7397_2;
    wire c7397;
    assign in7397_1 = {s4700[0]};
    assign in7397_2 = {s4701[0]};
    Full_Adder FA_7397(s7397, c7397, in7397_1, in7397_2, s4699[0]);
    wire[0:0] s7398, in7398_1, in7398_2;
    wire c7398;
    assign in7398_1 = {s4703[0]};
    assign in7398_2 = {s4704[0]};
    Full_Adder FA_7398(s7398, c7398, in7398_1, in7398_2, s4702[0]);
    wire[0:0] s7399, in7399_1, in7399_2;
    wire c7399;
    assign in7399_1 = {s4706[0]};
    assign in7399_2 = {s4707[0]};
    Full_Adder FA_7399(s7399, c7399, in7399_1, in7399_2, s4705[0]);
    wire[0:0] s7400, in7400_1, in7400_2;
    wire c7400;
    assign in7400_1 = {s4709[0]};
    assign in7400_2 = {s4710[0]};
    Full_Adder FA_7400(s7400, c7400, in7400_1, in7400_2, s4708[0]);
    wire[0:0] s7401, in7401_1, in7401_2;
    wire c7401;
    assign in7401_1 = {s4712[0]};
    assign in7401_2 = {s4713[0]};
    Full_Adder FA_7401(s7401, c7401, in7401_1, in7401_2, s4711[0]);
    wire[0:0] s7402, in7402_1, in7402_2;
    wire c7402;
    assign in7402_1 = {s4715[0]};
    assign in7402_2 = {s4716[0]};
    Full_Adder FA_7402(s7402, c7402, in7402_1, in7402_2, s4714[0]);
    wire[0:0] s7403, in7403_1, in7403_2;
    wire c7403;
    assign in7403_1 = {pp116[60]};
    assign in7403_2 = {pp117[59]};
    Full_Adder FA_7403(s7403, c7403, in7403_1, in7403_2, pp115[61]);
    wire[0:0] s7404, in7404_1, in7404_2;
    wire c7404;
    assign in7404_1 = {pp119[57]};
    assign in7404_2 = {pp120[56]};
    Full_Adder FA_7404(s7404, c7404, in7404_1, in7404_2, pp118[58]);
    wire[0:0] s7405, in7405_1, in7405_2;
    wire c7405;
    assign in7405_1 = {pp122[54]};
    assign in7405_2 = {pp123[53]};
    Full_Adder FA_7405(s7405, c7405, in7405_1, in7405_2, pp121[55]);
    wire[0:0] s7406, in7406_1, in7406_2;
    wire c7406;
    assign in7406_1 = {pp125[51]};
    assign in7406_2 = {pp126[50]};
    Full_Adder FA_7406(s7406, c7406, in7406_1, in7406_2, pp124[52]);
    wire[0:0] s7407, in7407_1, in7407_2;
    wire c7407;
    assign in7407_1 = {c4695};
    assign in7407_2 = {c4696};
    Full_Adder FA_7407(s7407, c7407, in7407_1, in7407_2, pp127[49]);
    wire[0:0] s7408, in7408_1, in7408_2;
    wire c7408;
    assign in7408_1 = {c4698};
    assign in7408_2 = {c4699};
    Full_Adder FA_7408(s7408, c7408, in7408_1, in7408_2, c4697);
    wire[0:0] s7409, in7409_1, in7409_2;
    wire c7409;
    assign in7409_1 = {c4701};
    assign in7409_2 = {c4702};
    Full_Adder FA_7409(s7409, c7409, in7409_1, in7409_2, c4700);
    wire[0:0] s7410, in7410_1, in7410_2;
    wire c7410;
    assign in7410_1 = {c4704};
    assign in7410_2 = {c4705};
    Full_Adder FA_7410(s7410, c7410, in7410_1, in7410_2, c4703);
    wire[0:0] s7411, in7411_1, in7411_2;
    wire c7411;
    assign in7411_1 = {c4707};
    assign in7411_2 = {c4708};
    Full_Adder FA_7411(s7411, c7411, in7411_1, in7411_2, c4706);
    wire[0:0] s7412, in7412_1, in7412_2;
    wire c7412;
    assign in7412_1 = {c4710};
    assign in7412_2 = {c4711};
    Full_Adder FA_7412(s7412, c7412, in7412_1, in7412_2, c4709);
    wire[0:0] s7413, in7413_1, in7413_2;
    wire c7413;
    assign in7413_1 = {c4713};
    assign in7413_2 = {c4714};
    Full_Adder FA_7413(s7413, c7413, in7413_1, in7413_2, c4712);
    wire[0:0] s7414, in7414_1, in7414_2;
    wire c7414;
    assign in7414_1 = {c4716};
    assign in7414_2 = {c4717};
    Full_Adder FA_7414(s7414, c7414, in7414_1, in7414_2, c4715);
    wire[0:0] s7415, in7415_1, in7415_2;
    wire c7415;
    assign in7415_1 = {s4719[0]};
    assign in7415_2 = {s4720[0]};
    Full_Adder FA_7415(s7415, c7415, in7415_1, in7415_2, s4718[0]);
    wire[0:0] s7416, in7416_1, in7416_2;
    wire c7416;
    assign in7416_1 = {s4722[0]};
    assign in7416_2 = {s4723[0]};
    Full_Adder FA_7416(s7416, c7416, in7416_1, in7416_2, s4721[0]);
    wire[0:0] s7417, in7417_1, in7417_2;
    wire c7417;
    assign in7417_1 = {s4725[0]};
    assign in7417_2 = {s4726[0]};
    Full_Adder FA_7417(s7417, c7417, in7417_1, in7417_2, s4724[0]);
    wire[0:0] s7418, in7418_1, in7418_2;
    wire c7418;
    assign in7418_1 = {s4728[0]};
    assign in7418_2 = {s4729[0]};
    Full_Adder FA_7418(s7418, c7418, in7418_1, in7418_2, s4727[0]);
    wire[0:0] s7419, in7419_1, in7419_2;
    wire c7419;
    assign in7419_1 = {s4731[0]};
    assign in7419_2 = {s4732[0]};
    Full_Adder FA_7419(s7419, c7419, in7419_1, in7419_2, s4730[0]);
    wire[0:0] s7420, in7420_1, in7420_2;
    wire c7420;
    assign in7420_1 = {s4734[0]};
    assign in7420_2 = {s4735[0]};
    Full_Adder FA_7420(s7420, c7420, in7420_1, in7420_2, s4733[0]);
    wire[0:0] s7421, in7421_1, in7421_2;
    wire c7421;
    assign in7421_1 = {s4737[0]};
    assign in7421_2 = {s4738[0]};
    Full_Adder FA_7421(s7421, c7421, in7421_1, in7421_2, s4736[0]);
    wire[0:0] s7422, in7422_1, in7422_2;
    wire c7422;
    assign in7422_1 = {pp114[63]};
    assign in7422_2 = {pp115[62]};
    Full_Adder FA_7422(s7422, c7422, in7422_1, in7422_2, pp113[64]);
    wire[0:0] s7423, in7423_1, in7423_2;
    wire c7423;
    assign in7423_1 = {pp117[60]};
    assign in7423_2 = {pp118[59]};
    Full_Adder FA_7423(s7423, c7423, in7423_1, in7423_2, pp116[61]);
    wire[0:0] s7424, in7424_1, in7424_2;
    wire c7424;
    assign in7424_1 = {pp120[57]};
    assign in7424_2 = {pp121[56]};
    Full_Adder FA_7424(s7424, c7424, in7424_1, in7424_2, pp119[58]);
    wire[0:0] s7425, in7425_1, in7425_2;
    wire c7425;
    assign in7425_1 = {pp123[54]};
    assign in7425_2 = {pp124[53]};
    Full_Adder FA_7425(s7425, c7425, in7425_1, in7425_2, pp122[55]);
    wire[0:0] s7426, in7426_1, in7426_2;
    wire c7426;
    assign in7426_1 = {pp126[51]};
    assign in7426_2 = {pp127[50]};
    Full_Adder FA_7426(s7426, c7426, in7426_1, in7426_2, pp125[52]);
    wire[0:0] s7427, in7427_1, in7427_2;
    wire c7427;
    assign in7427_1 = {c4719};
    assign in7427_2 = {c4720};
    Full_Adder FA_7427(s7427, c7427, in7427_1, in7427_2, c4718);
    wire[0:0] s7428, in7428_1, in7428_2;
    wire c7428;
    assign in7428_1 = {c4722};
    assign in7428_2 = {c4723};
    Full_Adder FA_7428(s7428, c7428, in7428_1, in7428_2, c4721);
    wire[0:0] s7429, in7429_1, in7429_2;
    wire c7429;
    assign in7429_1 = {c4725};
    assign in7429_2 = {c4726};
    Full_Adder FA_7429(s7429, c7429, in7429_1, in7429_2, c4724);
    wire[0:0] s7430, in7430_1, in7430_2;
    wire c7430;
    assign in7430_1 = {c4728};
    assign in7430_2 = {c4729};
    Full_Adder FA_7430(s7430, c7430, in7430_1, in7430_2, c4727);
    wire[0:0] s7431, in7431_1, in7431_2;
    wire c7431;
    assign in7431_1 = {c4731};
    assign in7431_2 = {c4732};
    Full_Adder FA_7431(s7431, c7431, in7431_1, in7431_2, c4730);
    wire[0:0] s7432, in7432_1, in7432_2;
    wire c7432;
    assign in7432_1 = {c4734};
    assign in7432_2 = {c4735};
    Full_Adder FA_7432(s7432, c7432, in7432_1, in7432_2, c4733);
    wire[0:0] s7433, in7433_1, in7433_2;
    wire c7433;
    assign in7433_1 = {c4737};
    assign in7433_2 = {c4738};
    Full_Adder FA_7433(s7433, c7433, in7433_1, in7433_2, c4736);
    wire[0:0] s7434, in7434_1, in7434_2;
    wire c7434;
    assign in7434_1 = {s4740[0]};
    assign in7434_2 = {s4741[0]};
    Full_Adder FA_7434(s7434, c7434, in7434_1, in7434_2, c4739);
    wire[0:0] s7435, in7435_1, in7435_2;
    wire c7435;
    assign in7435_1 = {s4743[0]};
    assign in7435_2 = {s4744[0]};
    Full_Adder FA_7435(s7435, c7435, in7435_1, in7435_2, s4742[0]);
    wire[0:0] s7436, in7436_1, in7436_2;
    wire c7436;
    assign in7436_1 = {s4746[0]};
    assign in7436_2 = {s4747[0]};
    Full_Adder FA_7436(s7436, c7436, in7436_1, in7436_2, s4745[0]);
    wire[0:0] s7437, in7437_1, in7437_2;
    wire c7437;
    assign in7437_1 = {s4749[0]};
    assign in7437_2 = {s4750[0]};
    Full_Adder FA_7437(s7437, c7437, in7437_1, in7437_2, s4748[0]);
    wire[0:0] s7438, in7438_1, in7438_2;
    wire c7438;
    assign in7438_1 = {s4752[0]};
    assign in7438_2 = {s4753[0]};
    Full_Adder FA_7438(s7438, c7438, in7438_1, in7438_2, s4751[0]);
    wire[0:0] s7439, in7439_1, in7439_2;
    wire c7439;
    assign in7439_1 = {s4755[0]};
    assign in7439_2 = {s4756[0]};
    Full_Adder FA_7439(s7439, c7439, in7439_1, in7439_2, s4754[0]);
    wire[0:0] s7440, in7440_1, in7440_2;
    wire c7440;
    assign in7440_1 = {s4758[0]};
    assign in7440_2 = {s4759[0]};
    Full_Adder FA_7440(s7440, c7440, in7440_1, in7440_2, s4757[0]);
    wire[0:0] s7441, in7441_1, in7441_2;
    wire c7441;
    assign in7441_1 = {pp112[66]};
    assign in7441_2 = {pp113[65]};
    Full_Adder FA_7441(s7441, c7441, in7441_1, in7441_2, pp111[67]);
    wire[0:0] s7442, in7442_1, in7442_2;
    wire c7442;
    assign in7442_1 = {pp115[63]};
    assign in7442_2 = {pp116[62]};
    Full_Adder FA_7442(s7442, c7442, in7442_1, in7442_2, pp114[64]);
    wire[0:0] s7443, in7443_1, in7443_2;
    wire c7443;
    assign in7443_1 = {pp118[60]};
    assign in7443_2 = {pp119[59]};
    Full_Adder FA_7443(s7443, c7443, in7443_1, in7443_2, pp117[61]);
    wire[0:0] s7444, in7444_1, in7444_2;
    wire c7444;
    assign in7444_1 = {pp121[57]};
    assign in7444_2 = {pp122[56]};
    Full_Adder FA_7444(s7444, c7444, in7444_1, in7444_2, pp120[58]);
    wire[0:0] s7445, in7445_1, in7445_2;
    wire c7445;
    assign in7445_1 = {pp124[54]};
    assign in7445_2 = {pp125[53]};
    Full_Adder FA_7445(s7445, c7445, in7445_1, in7445_2, pp123[55]);
    wire[0:0] s7446, in7446_1, in7446_2;
    wire c7446;
    assign in7446_1 = {pp127[51]};
    assign in7446_2 = {c4740};
    Full_Adder FA_7446(s7446, c7446, in7446_1, in7446_2, pp126[52]);
    wire[0:0] s7447, in7447_1, in7447_2;
    wire c7447;
    assign in7447_1 = {c4742};
    assign in7447_2 = {c4743};
    Full_Adder FA_7447(s7447, c7447, in7447_1, in7447_2, c4741);
    wire[0:0] s7448, in7448_1, in7448_2;
    wire c7448;
    assign in7448_1 = {c4745};
    assign in7448_2 = {c4746};
    Full_Adder FA_7448(s7448, c7448, in7448_1, in7448_2, c4744);
    wire[0:0] s7449, in7449_1, in7449_2;
    wire c7449;
    assign in7449_1 = {c4748};
    assign in7449_2 = {c4749};
    Full_Adder FA_7449(s7449, c7449, in7449_1, in7449_2, c4747);
    wire[0:0] s7450, in7450_1, in7450_2;
    wire c7450;
    assign in7450_1 = {c4751};
    assign in7450_2 = {c4752};
    Full_Adder FA_7450(s7450, c7450, in7450_1, in7450_2, c4750);
    wire[0:0] s7451, in7451_1, in7451_2;
    wire c7451;
    assign in7451_1 = {c4754};
    assign in7451_2 = {c4755};
    Full_Adder FA_7451(s7451, c7451, in7451_1, in7451_2, c4753);
    wire[0:0] s7452, in7452_1, in7452_2;
    wire c7452;
    assign in7452_1 = {c4757};
    assign in7452_2 = {c4758};
    Full_Adder FA_7452(s7452, c7452, in7452_1, in7452_2, c4756);
    wire[0:0] s7453, in7453_1, in7453_2;
    wire c7453;
    assign in7453_1 = {c4760};
    assign in7453_2 = {s4761[0]};
    Full_Adder FA_7453(s7453, c7453, in7453_1, in7453_2, c4759);
    wire[0:0] s7454, in7454_1, in7454_2;
    wire c7454;
    assign in7454_1 = {s4763[0]};
    assign in7454_2 = {s4764[0]};
    Full_Adder FA_7454(s7454, c7454, in7454_1, in7454_2, s4762[0]);
    wire[0:0] s7455, in7455_1, in7455_2;
    wire c7455;
    assign in7455_1 = {s4766[0]};
    assign in7455_2 = {s4767[0]};
    Full_Adder FA_7455(s7455, c7455, in7455_1, in7455_2, s4765[0]);
    wire[0:0] s7456, in7456_1, in7456_2;
    wire c7456;
    assign in7456_1 = {s4769[0]};
    assign in7456_2 = {s4770[0]};
    Full_Adder FA_7456(s7456, c7456, in7456_1, in7456_2, s4768[0]);
    wire[0:0] s7457, in7457_1, in7457_2;
    wire c7457;
    assign in7457_1 = {s4772[0]};
    assign in7457_2 = {s4773[0]};
    Full_Adder FA_7457(s7457, c7457, in7457_1, in7457_2, s4771[0]);
    wire[0:0] s7458, in7458_1, in7458_2;
    wire c7458;
    assign in7458_1 = {s4775[0]};
    assign in7458_2 = {s4776[0]};
    Full_Adder FA_7458(s7458, c7458, in7458_1, in7458_2, s4774[0]);
    wire[0:0] s7459, in7459_1, in7459_2;
    wire c7459;
    assign in7459_1 = {s4778[0]};
    assign in7459_2 = {s4779[0]};
    Full_Adder FA_7459(s7459, c7459, in7459_1, in7459_2, s4777[0]);
    wire[0:0] s7460, in7460_1, in7460_2;
    wire c7460;
    assign in7460_1 = {pp110[69]};
    assign in7460_2 = {pp111[68]};
    Full_Adder FA_7460(s7460, c7460, in7460_1, in7460_2, pp109[70]);
    wire[0:0] s7461, in7461_1, in7461_2;
    wire c7461;
    assign in7461_1 = {pp113[66]};
    assign in7461_2 = {pp114[65]};
    Full_Adder FA_7461(s7461, c7461, in7461_1, in7461_2, pp112[67]);
    wire[0:0] s7462, in7462_1, in7462_2;
    wire c7462;
    assign in7462_1 = {pp116[63]};
    assign in7462_2 = {pp117[62]};
    Full_Adder FA_7462(s7462, c7462, in7462_1, in7462_2, pp115[64]);
    wire[0:0] s7463, in7463_1, in7463_2;
    wire c7463;
    assign in7463_1 = {pp119[60]};
    assign in7463_2 = {pp120[59]};
    Full_Adder FA_7463(s7463, c7463, in7463_1, in7463_2, pp118[61]);
    wire[0:0] s7464, in7464_1, in7464_2;
    wire c7464;
    assign in7464_1 = {pp122[57]};
    assign in7464_2 = {pp123[56]};
    Full_Adder FA_7464(s7464, c7464, in7464_1, in7464_2, pp121[58]);
    wire[0:0] s7465, in7465_1, in7465_2;
    wire c7465;
    assign in7465_1 = {pp125[54]};
    assign in7465_2 = {pp126[53]};
    Full_Adder FA_7465(s7465, c7465, in7465_1, in7465_2, pp124[55]);
    wire[0:0] s7466, in7466_1, in7466_2;
    wire c7466;
    assign in7466_1 = {c4761};
    assign in7466_2 = {c4762};
    Full_Adder FA_7466(s7466, c7466, in7466_1, in7466_2, pp127[52]);
    wire[0:0] s7467, in7467_1, in7467_2;
    wire c7467;
    assign in7467_1 = {c4764};
    assign in7467_2 = {c4765};
    Full_Adder FA_7467(s7467, c7467, in7467_1, in7467_2, c4763);
    wire[0:0] s7468, in7468_1, in7468_2;
    wire c7468;
    assign in7468_1 = {c4767};
    assign in7468_2 = {c4768};
    Full_Adder FA_7468(s7468, c7468, in7468_1, in7468_2, c4766);
    wire[0:0] s7469, in7469_1, in7469_2;
    wire c7469;
    assign in7469_1 = {c4770};
    assign in7469_2 = {c4771};
    Full_Adder FA_7469(s7469, c7469, in7469_1, in7469_2, c4769);
    wire[0:0] s7470, in7470_1, in7470_2;
    wire c7470;
    assign in7470_1 = {c4773};
    assign in7470_2 = {c4774};
    Full_Adder FA_7470(s7470, c7470, in7470_1, in7470_2, c4772);
    wire[0:0] s7471, in7471_1, in7471_2;
    wire c7471;
    assign in7471_1 = {c4776};
    assign in7471_2 = {c4777};
    Full_Adder FA_7471(s7471, c7471, in7471_1, in7471_2, c4775);
    wire[0:0] s7472, in7472_1, in7472_2;
    wire c7472;
    assign in7472_1 = {c4779};
    assign in7472_2 = {c4780};
    Full_Adder FA_7472(s7472, c7472, in7472_1, in7472_2, c4778);
    wire[0:0] s7473, in7473_1, in7473_2;
    wire c7473;
    assign in7473_1 = {s4782[0]};
    assign in7473_2 = {s4783[0]};
    Full_Adder FA_7473(s7473, c7473, in7473_1, in7473_2, s4781[0]);
    wire[0:0] s7474, in7474_1, in7474_2;
    wire c7474;
    assign in7474_1 = {s4785[0]};
    assign in7474_2 = {s4786[0]};
    Full_Adder FA_7474(s7474, c7474, in7474_1, in7474_2, s4784[0]);
    wire[0:0] s7475, in7475_1, in7475_2;
    wire c7475;
    assign in7475_1 = {s4788[0]};
    assign in7475_2 = {s4789[0]};
    Full_Adder FA_7475(s7475, c7475, in7475_1, in7475_2, s4787[0]);
    wire[0:0] s7476, in7476_1, in7476_2;
    wire c7476;
    assign in7476_1 = {s4791[0]};
    assign in7476_2 = {s4792[0]};
    Full_Adder FA_7476(s7476, c7476, in7476_1, in7476_2, s4790[0]);
    wire[0:0] s7477, in7477_1, in7477_2;
    wire c7477;
    assign in7477_1 = {s4794[0]};
    assign in7477_2 = {s4795[0]};
    Full_Adder FA_7477(s7477, c7477, in7477_1, in7477_2, s4793[0]);
    wire[0:0] s7478, in7478_1, in7478_2;
    wire c7478;
    assign in7478_1 = {s4797[0]};
    assign in7478_2 = {s4798[0]};
    Full_Adder FA_7478(s7478, c7478, in7478_1, in7478_2, s4796[0]);
    wire[0:0] s7479, in7479_1, in7479_2;
    wire c7479;
    assign in7479_1 = {pp108[72]};
    assign in7479_2 = {pp109[71]};
    Full_Adder FA_7479(s7479, c7479, in7479_1, in7479_2, pp107[73]);
    wire[0:0] s7480, in7480_1, in7480_2;
    wire c7480;
    assign in7480_1 = {pp111[69]};
    assign in7480_2 = {pp112[68]};
    Full_Adder FA_7480(s7480, c7480, in7480_1, in7480_2, pp110[70]);
    wire[0:0] s7481, in7481_1, in7481_2;
    wire c7481;
    assign in7481_1 = {pp114[66]};
    assign in7481_2 = {pp115[65]};
    Full_Adder FA_7481(s7481, c7481, in7481_1, in7481_2, pp113[67]);
    wire[0:0] s7482, in7482_1, in7482_2;
    wire c7482;
    assign in7482_1 = {pp117[63]};
    assign in7482_2 = {pp118[62]};
    Full_Adder FA_7482(s7482, c7482, in7482_1, in7482_2, pp116[64]);
    wire[0:0] s7483, in7483_1, in7483_2;
    wire c7483;
    assign in7483_1 = {pp120[60]};
    assign in7483_2 = {pp121[59]};
    Full_Adder FA_7483(s7483, c7483, in7483_1, in7483_2, pp119[61]);
    wire[0:0] s7484, in7484_1, in7484_2;
    wire c7484;
    assign in7484_1 = {pp123[57]};
    assign in7484_2 = {pp124[56]};
    Full_Adder FA_7484(s7484, c7484, in7484_1, in7484_2, pp122[58]);
    wire[0:0] s7485, in7485_1, in7485_2;
    wire c7485;
    assign in7485_1 = {pp126[54]};
    assign in7485_2 = {pp127[53]};
    Full_Adder FA_7485(s7485, c7485, in7485_1, in7485_2, pp125[55]);
    wire[0:0] s7486, in7486_1, in7486_2;
    wire c7486;
    assign in7486_1 = {c4782};
    assign in7486_2 = {c4783};
    Full_Adder FA_7486(s7486, c7486, in7486_1, in7486_2, c4781);
    wire[0:0] s7487, in7487_1, in7487_2;
    wire c7487;
    assign in7487_1 = {c4785};
    assign in7487_2 = {c4786};
    Full_Adder FA_7487(s7487, c7487, in7487_1, in7487_2, c4784);
    wire[0:0] s7488, in7488_1, in7488_2;
    wire c7488;
    assign in7488_1 = {c4788};
    assign in7488_2 = {c4789};
    Full_Adder FA_7488(s7488, c7488, in7488_1, in7488_2, c4787);
    wire[0:0] s7489, in7489_1, in7489_2;
    wire c7489;
    assign in7489_1 = {c4791};
    assign in7489_2 = {c4792};
    Full_Adder FA_7489(s7489, c7489, in7489_1, in7489_2, c4790);
    wire[0:0] s7490, in7490_1, in7490_2;
    wire c7490;
    assign in7490_1 = {c4794};
    assign in7490_2 = {c4795};
    Full_Adder FA_7490(s7490, c7490, in7490_1, in7490_2, c4793);
    wire[0:0] s7491, in7491_1, in7491_2;
    wire c7491;
    assign in7491_1 = {c4797};
    assign in7491_2 = {c4798};
    Full_Adder FA_7491(s7491, c7491, in7491_1, in7491_2, c4796);
    wire[0:0] s7492, in7492_1, in7492_2;
    wire c7492;
    assign in7492_1 = {s4800[0]};
    assign in7492_2 = {s4801[0]};
    Full_Adder FA_7492(s7492, c7492, in7492_1, in7492_2, c4799);
    wire[0:0] s7493, in7493_1, in7493_2;
    wire c7493;
    assign in7493_1 = {s4803[0]};
    assign in7493_2 = {s4804[0]};
    Full_Adder FA_7493(s7493, c7493, in7493_1, in7493_2, s4802[0]);
    wire[0:0] s7494, in7494_1, in7494_2;
    wire c7494;
    assign in7494_1 = {s4806[0]};
    assign in7494_2 = {s4807[0]};
    Full_Adder FA_7494(s7494, c7494, in7494_1, in7494_2, s4805[0]);
    wire[0:0] s7495, in7495_1, in7495_2;
    wire c7495;
    assign in7495_1 = {s4809[0]};
    assign in7495_2 = {s4810[0]};
    Full_Adder FA_7495(s7495, c7495, in7495_1, in7495_2, s4808[0]);
    wire[0:0] s7496, in7496_1, in7496_2;
    wire c7496;
    assign in7496_1 = {s4812[0]};
    assign in7496_2 = {s4813[0]};
    Full_Adder FA_7496(s7496, c7496, in7496_1, in7496_2, s4811[0]);
    wire[0:0] s7497, in7497_1, in7497_2;
    wire c7497;
    assign in7497_1 = {s4815[0]};
    assign in7497_2 = {s4816[0]};
    Full_Adder FA_7497(s7497, c7497, in7497_1, in7497_2, s4814[0]);
    wire[0:0] s7498, in7498_1, in7498_2;
    wire c7498;
    assign in7498_1 = {pp106[75]};
    assign in7498_2 = {pp107[74]};
    Full_Adder FA_7498(s7498, c7498, in7498_1, in7498_2, pp105[76]);
    wire[0:0] s7499, in7499_1, in7499_2;
    wire c7499;
    assign in7499_1 = {pp109[72]};
    assign in7499_2 = {pp110[71]};
    Full_Adder FA_7499(s7499, c7499, in7499_1, in7499_2, pp108[73]);
    wire[0:0] s7500, in7500_1, in7500_2;
    wire c7500;
    assign in7500_1 = {pp112[69]};
    assign in7500_2 = {pp113[68]};
    Full_Adder FA_7500(s7500, c7500, in7500_1, in7500_2, pp111[70]);
    wire[0:0] s7501, in7501_1, in7501_2;
    wire c7501;
    assign in7501_1 = {pp115[66]};
    assign in7501_2 = {pp116[65]};
    Full_Adder FA_7501(s7501, c7501, in7501_1, in7501_2, pp114[67]);
    wire[0:0] s7502, in7502_1, in7502_2;
    wire c7502;
    assign in7502_1 = {pp118[63]};
    assign in7502_2 = {pp119[62]};
    Full_Adder FA_7502(s7502, c7502, in7502_1, in7502_2, pp117[64]);
    wire[0:0] s7503, in7503_1, in7503_2;
    wire c7503;
    assign in7503_1 = {pp121[60]};
    assign in7503_2 = {pp122[59]};
    Full_Adder FA_7503(s7503, c7503, in7503_1, in7503_2, pp120[61]);
    wire[0:0] s7504, in7504_1, in7504_2;
    wire c7504;
    assign in7504_1 = {pp124[57]};
    assign in7504_2 = {pp125[56]};
    Full_Adder FA_7504(s7504, c7504, in7504_1, in7504_2, pp123[58]);
    wire[0:0] s7505, in7505_1, in7505_2;
    wire c7505;
    assign in7505_1 = {pp127[54]};
    assign in7505_2 = {c4800};
    Full_Adder FA_7505(s7505, c7505, in7505_1, in7505_2, pp126[55]);
    wire[0:0] s7506, in7506_1, in7506_2;
    wire c7506;
    assign in7506_1 = {c4802};
    assign in7506_2 = {c4803};
    Full_Adder FA_7506(s7506, c7506, in7506_1, in7506_2, c4801);
    wire[0:0] s7507, in7507_1, in7507_2;
    wire c7507;
    assign in7507_1 = {c4805};
    assign in7507_2 = {c4806};
    Full_Adder FA_7507(s7507, c7507, in7507_1, in7507_2, c4804);
    wire[0:0] s7508, in7508_1, in7508_2;
    wire c7508;
    assign in7508_1 = {c4808};
    assign in7508_2 = {c4809};
    Full_Adder FA_7508(s7508, c7508, in7508_1, in7508_2, c4807);
    wire[0:0] s7509, in7509_1, in7509_2;
    wire c7509;
    assign in7509_1 = {c4811};
    assign in7509_2 = {c4812};
    Full_Adder FA_7509(s7509, c7509, in7509_1, in7509_2, c4810);
    wire[0:0] s7510, in7510_1, in7510_2;
    wire c7510;
    assign in7510_1 = {c4814};
    assign in7510_2 = {c4815};
    Full_Adder FA_7510(s7510, c7510, in7510_1, in7510_2, c4813);
    wire[0:0] s7511, in7511_1, in7511_2;
    wire c7511;
    assign in7511_1 = {c4817};
    assign in7511_2 = {s4818[0]};
    Full_Adder FA_7511(s7511, c7511, in7511_1, in7511_2, c4816);
    wire[0:0] s7512, in7512_1, in7512_2;
    wire c7512;
    assign in7512_1 = {s4820[0]};
    assign in7512_2 = {s4821[0]};
    Full_Adder FA_7512(s7512, c7512, in7512_1, in7512_2, s4819[0]);
    wire[0:0] s7513, in7513_1, in7513_2;
    wire c7513;
    assign in7513_1 = {s4823[0]};
    assign in7513_2 = {s4824[0]};
    Full_Adder FA_7513(s7513, c7513, in7513_1, in7513_2, s4822[0]);
    wire[0:0] s7514, in7514_1, in7514_2;
    wire c7514;
    assign in7514_1 = {s4826[0]};
    assign in7514_2 = {s4827[0]};
    Full_Adder FA_7514(s7514, c7514, in7514_1, in7514_2, s4825[0]);
    wire[0:0] s7515, in7515_1, in7515_2;
    wire c7515;
    assign in7515_1 = {s4829[0]};
    assign in7515_2 = {s4830[0]};
    Full_Adder FA_7515(s7515, c7515, in7515_1, in7515_2, s4828[0]);
    wire[0:0] s7516, in7516_1, in7516_2;
    wire c7516;
    assign in7516_1 = {s4832[0]};
    assign in7516_2 = {s4833[0]};
    Full_Adder FA_7516(s7516, c7516, in7516_1, in7516_2, s4831[0]);
    wire[0:0] s7517, in7517_1, in7517_2;
    wire c7517;
    assign in7517_1 = {pp104[78]};
    assign in7517_2 = {pp105[77]};
    Full_Adder FA_7517(s7517, c7517, in7517_1, in7517_2, pp103[79]);
    wire[0:0] s7518, in7518_1, in7518_2;
    wire c7518;
    assign in7518_1 = {pp107[75]};
    assign in7518_2 = {pp108[74]};
    Full_Adder FA_7518(s7518, c7518, in7518_1, in7518_2, pp106[76]);
    wire[0:0] s7519, in7519_1, in7519_2;
    wire c7519;
    assign in7519_1 = {pp110[72]};
    assign in7519_2 = {pp111[71]};
    Full_Adder FA_7519(s7519, c7519, in7519_1, in7519_2, pp109[73]);
    wire[0:0] s7520, in7520_1, in7520_2;
    wire c7520;
    assign in7520_1 = {pp113[69]};
    assign in7520_2 = {pp114[68]};
    Full_Adder FA_7520(s7520, c7520, in7520_1, in7520_2, pp112[70]);
    wire[0:0] s7521, in7521_1, in7521_2;
    wire c7521;
    assign in7521_1 = {pp116[66]};
    assign in7521_2 = {pp117[65]};
    Full_Adder FA_7521(s7521, c7521, in7521_1, in7521_2, pp115[67]);
    wire[0:0] s7522, in7522_1, in7522_2;
    wire c7522;
    assign in7522_1 = {pp119[63]};
    assign in7522_2 = {pp120[62]};
    Full_Adder FA_7522(s7522, c7522, in7522_1, in7522_2, pp118[64]);
    wire[0:0] s7523, in7523_1, in7523_2;
    wire c7523;
    assign in7523_1 = {pp122[60]};
    assign in7523_2 = {pp123[59]};
    Full_Adder FA_7523(s7523, c7523, in7523_1, in7523_2, pp121[61]);
    wire[0:0] s7524, in7524_1, in7524_2;
    wire c7524;
    assign in7524_1 = {pp125[57]};
    assign in7524_2 = {pp126[56]};
    Full_Adder FA_7524(s7524, c7524, in7524_1, in7524_2, pp124[58]);
    wire[0:0] s7525, in7525_1, in7525_2;
    wire c7525;
    assign in7525_1 = {c4818};
    assign in7525_2 = {c4819};
    Full_Adder FA_7525(s7525, c7525, in7525_1, in7525_2, pp127[55]);
    wire[0:0] s7526, in7526_1, in7526_2;
    wire c7526;
    assign in7526_1 = {c4821};
    assign in7526_2 = {c4822};
    Full_Adder FA_7526(s7526, c7526, in7526_1, in7526_2, c4820);
    wire[0:0] s7527, in7527_1, in7527_2;
    wire c7527;
    assign in7527_1 = {c4824};
    assign in7527_2 = {c4825};
    Full_Adder FA_7527(s7527, c7527, in7527_1, in7527_2, c4823);
    wire[0:0] s7528, in7528_1, in7528_2;
    wire c7528;
    assign in7528_1 = {c4827};
    assign in7528_2 = {c4828};
    Full_Adder FA_7528(s7528, c7528, in7528_1, in7528_2, c4826);
    wire[0:0] s7529, in7529_1, in7529_2;
    wire c7529;
    assign in7529_1 = {c4830};
    assign in7529_2 = {c4831};
    Full_Adder FA_7529(s7529, c7529, in7529_1, in7529_2, c4829);
    wire[0:0] s7530, in7530_1, in7530_2;
    wire c7530;
    assign in7530_1 = {c4833};
    assign in7530_2 = {c4834};
    Full_Adder FA_7530(s7530, c7530, in7530_1, in7530_2, c4832);
    wire[0:0] s7531, in7531_1, in7531_2;
    wire c7531;
    assign in7531_1 = {s4836[0]};
    assign in7531_2 = {s4837[0]};
    Full_Adder FA_7531(s7531, c7531, in7531_1, in7531_2, s4835[0]);
    wire[0:0] s7532, in7532_1, in7532_2;
    wire c7532;
    assign in7532_1 = {s4839[0]};
    assign in7532_2 = {s4840[0]};
    Full_Adder FA_7532(s7532, c7532, in7532_1, in7532_2, s4838[0]);
    wire[0:0] s7533, in7533_1, in7533_2;
    wire c7533;
    assign in7533_1 = {s4842[0]};
    assign in7533_2 = {s4843[0]};
    Full_Adder FA_7533(s7533, c7533, in7533_1, in7533_2, s4841[0]);
    wire[0:0] s7534, in7534_1, in7534_2;
    wire c7534;
    assign in7534_1 = {s4845[0]};
    assign in7534_2 = {s4846[0]};
    Full_Adder FA_7534(s7534, c7534, in7534_1, in7534_2, s4844[0]);
    wire[0:0] s7535, in7535_1, in7535_2;
    wire c7535;
    assign in7535_1 = {s4848[0]};
    assign in7535_2 = {s4849[0]};
    Full_Adder FA_7535(s7535, c7535, in7535_1, in7535_2, s4847[0]);
    wire[0:0] s7536, in7536_1, in7536_2;
    wire c7536;
    assign in7536_1 = {pp102[81]};
    assign in7536_2 = {pp103[80]};
    Full_Adder FA_7536(s7536, c7536, in7536_1, in7536_2, pp101[82]);
    wire[0:0] s7537, in7537_1, in7537_2;
    wire c7537;
    assign in7537_1 = {pp105[78]};
    assign in7537_2 = {pp106[77]};
    Full_Adder FA_7537(s7537, c7537, in7537_1, in7537_2, pp104[79]);
    wire[0:0] s7538, in7538_1, in7538_2;
    wire c7538;
    assign in7538_1 = {pp108[75]};
    assign in7538_2 = {pp109[74]};
    Full_Adder FA_7538(s7538, c7538, in7538_1, in7538_2, pp107[76]);
    wire[0:0] s7539, in7539_1, in7539_2;
    wire c7539;
    assign in7539_1 = {pp111[72]};
    assign in7539_2 = {pp112[71]};
    Full_Adder FA_7539(s7539, c7539, in7539_1, in7539_2, pp110[73]);
    wire[0:0] s7540, in7540_1, in7540_2;
    wire c7540;
    assign in7540_1 = {pp114[69]};
    assign in7540_2 = {pp115[68]};
    Full_Adder FA_7540(s7540, c7540, in7540_1, in7540_2, pp113[70]);
    wire[0:0] s7541, in7541_1, in7541_2;
    wire c7541;
    assign in7541_1 = {pp117[66]};
    assign in7541_2 = {pp118[65]};
    Full_Adder FA_7541(s7541, c7541, in7541_1, in7541_2, pp116[67]);
    wire[0:0] s7542, in7542_1, in7542_2;
    wire c7542;
    assign in7542_1 = {pp120[63]};
    assign in7542_2 = {pp121[62]};
    Full_Adder FA_7542(s7542, c7542, in7542_1, in7542_2, pp119[64]);
    wire[0:0] s7543, in7543_1, in7543_2;
    wire c7543;
    assign in7543_1 = {pp123[60]};
    assign in7543_2 = {pp124[59]};
    Full_Adder FA_7543(s7543, c7543, in7543_1, in7543_2, pp122[61]);
    wire[0:0] s7544, in7544_1, in7544_2;
    wire c7544;
    assign in7544_1 = {pp126[57]};
    assign in7544_2 = {pp127[56]};
    Full_Adder FA_7544(s7544, c7544, in7544_1, in7544_2, pp125[58]);
    wire[0:0] s7545, in7545_1, in7545_2;
    wire c7545;
    assign in7545_1 = {c4836};
    assign in7545_2 = {c4837};
    Full_Adder FA_7545(s7545, c7545, in7545_1, in7545_2, c4835);
    wire[0:0] s7546, in7546_1, in7546_2;
    wire c7546;
    assign in7546_1 = {c4839};
    assign in7546_2 = {c4840};
    Full_Adder FA_7546(s7546, c7546, in7546_1, in7546_2, c4838);
    wire[0:0] s7547, in7547_1, in7547_2;
    wire c7547;
    assign in7547_1 = {c4842};
    assign in7547_2 = {c4843};
    Full_Adder FA_7547(s7547, c7547, in7547_1, in7547_2, c4841);
    wire[0:0] s7548, in7548_1, in7548_2;
    wire c7548;
    assign in7548_1 = {c4845};
    assign in7548_2 = {c4846};
    Full_Adder FA_7548(s7548, c7548, in7548_1, in7548_2, c4844);
    wire[0:0] s7549, in7549_1, in7549_2;
    wire c7549;
    assign in7549_1 = {c4848};
    assign in7549_2 = {c4849};
    Full_Adder FA_7549(s7549, c7549, in7549_1, in7549_2, c4847);
    wire[0:0] s7550, in7550_1, in7550_2;
    wire c7550;
    assign in7550_1 = {s4851[0]};
    assign in7550_2 = {s4852[0]};
    Full_Adder FA_7550(s7550, c7550, in7550_1, in7550_2, c4850);
    wire[0:0] s7551, in7551_1, in7551_2;
    wire c7551;
    assign in7551_1 = {s4854[0]};
    assign in7551_2 = {s4855[0]};
    Full_Adder FA_7551(s7551, c7551, in7551_1, in7551_2, s4853[0]);
    wire[0:0] s7552, in7552_1, in7552_2;
    wire c7552;
    assign in7552_1 = {s4857[0]};
    assign in7552_2 = {s4858[0]};
    Full_Adder FA_7552(s7552, c7552, in7552_1, in7552_2, s4856[0]);
    wire[0:0] s7553, in7553_1, in7553_2;
    wire c7553;
    assign in7553_1 = {s4860[0]};
    assign in7553_2 = {s4861[0]};
    Full_Adder FA_7553(s7553, c7553, in7553_1, in7553_2, s4859[0]);
    wire[0:0] s7554, in7554_1, in7554_2;
    wire c7554;
    assign in7554_1 = {s4863[0]};
    assign in7554_2 = {s4864[0]};
    Full_Adder FA_7554(s7554, c7554, in7554_1, in7554_2, s4862[0]);
    wire[0:0] s7555, in7555_1, in7555_2;
    wire c7555;
    assign in7555_1 = {pp100[84]};
    assign in7555_2 = {pp101[83]};
    Full_Adder FA_7555(s7555, c7555, in7555_1, in7555_2, pp99[85]);
    wire[0:0] s7556, in7556_1, in7556_2;
    wire c7556;
    assign in7556_1 = {pp103[81]};
    assign in7556_2 = {pp104[80]};
    Full_Adder FA_7556(s7556, c7556, in7556_1, in7556_2, pp102[82]);
    wire[0:0] s7557, in7557_1, in7557_2;
    wire c7557;
    assign in7557_1 = {pp106[78]};
    assign in7557_2 = {pp107[77]};
    Full_Adder FA_7557(s7557, c7557, in7557_1, in7557_2, pp105[79]);
    wire[0:0] s7558, in7558_1, in7558_2;
    wire c7558;
    assign in7558_1 = {pp109[75]};
    assign in7558_2 = {pp110[74]};
    Full_Adder FA_7558(s7558, c7558, in7558_1, in7558_2, pp108[76]);
    wire[0:0] s7559, in7559_1, in7559_2;
    wire c7559;
    assign in7559_1 = {pp112[72]};
    assign in7559_2 = {pp113[71]};
    Full_Adder FA_7559(s7559, c7559, in7559_1, in7559_2, pp111[73]);
    wire[0:0] s7560, in7560_1, in7560_2;
    wire c7560;
    assign in7560_1 = {pp115[69]};
    assign in7560_2 = {pp116[68]};
    Full_Adder FA_7560(s7560, c7560, in7560_1, in7560_2, pp114[70]);
    wire[0:0] s7561, in7561_1, in7561_2;
    wire c7561;
    assign in7561_1 = {pp118[66]};
    assign in7561_2 = {pp119[65]};
    Full_Adder FA_7561(s7561, c7561, in7561_1, in7561_2, pp117[67]);
    wire[0:0] s7562, in7562_1, in7562_2;
    wire c7562;
    assign in7562_1 = {pp121[63]};
    assign in7562_2 = {pp122[62]};
    Full_Adder FA_7562(s7562, c7562, in7562_1, in7562_2, pp120[64]);
    wire[0:0] s7563, in7563_1, in7563_2;
    wire c7563;
    assign in7563_1 = {pp124[60]};
    assign in7563_2 = {pp125[59]};
    Full_Adder FA_7563(s7563, c7563, in7563_1, in7563_2, pp123[61]);
    wire[0:0] s7564, in7564_1, in7564_2;
    wire c7564;
    assign in7564_1 = {pp127[57]};
    assign in7564_2 = {c4851};
    Full_Adder FA_7564(s7564, c7564, in7564_1, in7564_2, pp126[58]);
    wire[0:0] s7565, in7565_1, in7565_2;
    wire c7565;
    assign in7565_1 = {c4853};
    assign in7565_2 = {c4854};
    Full_Adder FA_7565(s7565, c7565, in7565_1, in7565_2, c4852);
    wire[0:0] s7566, in7566_1, in7566_2;
    wire c7566;
    assign in7566_1 = {c4856};
    assign in7566_2 = {c4857};
    Full_Adder FA_7566(s7566, c7566, in7566_1, in7566_2, c4855);
    wire[0:0] s7567, in7567_1, in7567_2;
    wire c7567;
    assign in7567_1 = {c4859};
    assign in7567_2 = {c4860};
    Full_Adder FA_7567(s7567, c7567, in7567_1, in7567_2, c4858);
    wire[0:0] s7568, in7568_1, in7568_2;
    wire c7568;
    assign in7568_1 = {c4862};
    assign in7568_2 = {c4863};
    Full_Adder FA_7568(s7568, c7568, in7568_1, in7568_2, c4861);
    wire[0:0] s7569, in7569_1, in7569_2;
    wire c7569;
    assign in7569_1 = {c4865};
    assign in7569_2 = {s4866[0]};
    Full_Adder FA_7569(s7569, c7569, in7569_1, in7569_2, c4864);
    wire[0:0] s7570, in7570_1, in7570_2;
    wire c7570;
    assign in7570_1 = {s4868[0]};
    assign in7570_2 = {s4869[0]};
    Full_Adder FA_7570(s7570, c7570, in7570_1, in7570_2, s4867[0]);
    wire[0:0] s7571, in7571_1, in7571_2;
    wire c7571;
    assign in7571_1 = {s4871[0]};
    assign in7571_2 = {s4872[0]};
    Full_Adder FA_7571(s7571, c7571, in7571_1, in7571_2, s4870[0]);
    wire[0:0] s7572, in7572_1, in7572_2;
    wire c7572;
    assign in7572_1 = {s4874[0]};
    assign in7572_2 = {s4875[0]};
    Full_Adder FA_7572(s7572, c7572, in7572_1, in7572_2, s4873[0]);
    wire[0:0] s7573, in7573_1, in7573_2;
    wire c7573;
    assign in7573_1 = {s4877[0]};
    assign in7573_2 = {s4878[0]};
    Full_Adder FA_7573(s7573, c7573, in7573_1, in7573_2, s4876[0]);
    wire[0:0] s7574, in7574_1, in7574_2;
    wire c7574;
    assign in7574_1 = {pp98[87]};
    assign in7574_2 = {pp99[86]};
    Full_Adder FA_7574(s7574, c7574, in7574_1, in7574_2, pp97[88]);
    wire[0:0] s7575, in7575_1, in7575_2;
    wire c7575;
    assign in7575_1 = {pp101[84]};
    assign in7575_2 = {pp102[83]};
    Full_Adder FA_7575(s7575, c7575, in7575_1, in7575_2, pp100[85]);
    wire[0:0] s7576, in7576_1, in7576_2;
    wire c7576;
    assign in7576_1 = {pp104[81]};
    assign in7576_2 = {pp105[80]};
    Full_Adder FA_7576(s7576, c7576, in7576_1, in7576_2, pp103[82]);
    wire[0:0] s7577, in7577_1, in7577_2;
    wire c7577;
    assign in7577_1 = {pp107[78]};
    assign in7577_2 = {pp108[77]};
    Full_Adder FA_7577(s7577, c7577, in7577_1, in7577_2, pp106[79]);
    wire[0:0] s7578, in7578_1, in7578_2;
    wire c7578;
    assign in7578_1 = {pp110[75]};
    assign in7578_2 = {pp111[74]};
    Full_Adder FA_7578(s7578, c7578, in7578_1, in7578_2, pp109[76]);
    wire[0:0] s7579, in7579_1, in7579_2;
    wire c7579;
    assign in7579_1 = {pp113[72]};
    assign in7579_2 = {pp114[71]};
    Full_Adder FA_7579(s7579, c7579, in7579_1, in7579_2, pp112[73]);
    wire[0:0] s7580, in7580_1, in7580_2;
    wire c7580;
    assign in7580_1 = {pp116[69]};
    assign in7580_2 = {pp117[68]};
    Full_Adder FA_7580(s7580, c7580, in7580_1, in7580_2, pp115[70]);
    wire[0:0] s7581, in7581_1, in7581_2;
    wire c7581;
    assign in7581_1 = {pp119[66]};
    assign in7581_2 = {pp120[65]};
    Full_Adder FA_7581(s7581, c7581, in7581_1, in7581_2, pp118[67]);
    wire[0:0] s7582, in7582_1, in7582_2;
    wire c7582;
    assign in7582_1 = {pp122[63]};
    assign in7582_2 = {pp123[62]};
    Full_Adder FA_7582(s7582, c7582, in7582_1, in7582_2, pp121[64]);
    wire[0:0] s7583, in7583_1, in7583_2;
    wire c7583;
    assign in7583_1 = {pp125[60]};
    assign in7583_2 = {pp126[59]};
    Full_Adder FA_7583(s7583, c7583, in7583_1, in7583_2, pp124[61]);
    wire[0:0] s7584, in7584_1, in7584_2;
    wire c7584;
    assign in7584_1 = {c4866};
    assign in7584_2 = {c4867};
    Full_Adder FA_7584(s7584, c7584, in7584_1, in7584_2, pp127[58]);
    wire[0:0] s7585, in7585_1, in7585_2;
    wire c7585;
    assign in7585_1 = {c4869};
    assign in7585_2 = {c4870};
    Full_Adder FA_7585(s7585, c7585, in7585_1, in7585_2, c4868);
    wire[0:0] s7586, in7586_1, in7586_2;
    wire c7586;
    assign in7586_1 = {c4872};
    assign in7586_2 = {c4873};
    Full_Adder FA_7586(s7586, c7586, in7586_1, in7586_2, c4871);
    wire[0:0] s7587, in7587_1, in7587_2;
    wire c7587;
    assign in7587_1 = {c4875};
    assign in7587_2 = {c4876};
    Full_Adder FA_7587(s7587, c7587, in7587_1, in7587_2, c4874);
    wire[0:0] s7588, in7588_1, in7588_2;
    wire c7588;
    assign in7588_1 = {c4878};
    assign in7588_2 = {c4879};
    Full_Adder FA_7588(s7588, c7588, in7588_1, in7588_2, c4877);
    wire[0:0] s7589, in7589_1, in7589_2;
    wire c7589;
    assign in7589_1 = {s4881[0]};
    assign in7589_2 = {s4882[0]};
    Full_Adder FA_7589(s7589, c7589, in7589_1, in7589_2, s4880[0]);
    wire[0:0] s7590, in7590_1, in7590_2;
    wire c7590;
    assign in7590_1 = {s4884[0]};
    assign in7590_2 = {s4885[0]};
    Full_Adder FA_7590(s7590, c7590, in7590_1, in7590_2, s4883[0]);
    wire[0:0] s7591, in7591_1, in7591_2;
    wire c7591;
    assign in7591_1 = {s4887[0]};
    assign in7591_2 = {s4888[0]};
    Full_Adder FA_7591(s7591, c7591, in7591_1, in7591_2, s4886[0]);
    wire[0:0] s7592, in7592_1, in7592_2;
    wire c7592;
    assign in7592_1 = {s4890[0]};
    assign in7592_2 = {s4891[0]};
    Full_Adder FA_7592(s7592, c7592, in7592_1, in7592_2, s4889[0]);
    wire[0:0] s7593, in7593_1, in7593_2;
    wire c7593;
    assign in7593_1 = {pp96[90]};
    assign in7593_2 = {pp97[89]};
    Full_Adder FA_7593(s7593, c7593, in7593_1, in7593_2, pp95[91]);
    wire[0:0] s7594, in7594_1, in7594_2;
    wire c7594;
    assign in7594_1 = {pp99[87]};
    assign in7594_2 = {pp100[86]};
    Full_Adder FA_7594(s7594, c7594, in7594_1, in7594_2, pp98[88]);
    wire[0:0] s7595, in7595_1, in7595_2;
    wire c7595;
    assign in7595_1 = {pp102[84]};
    assign in7595_2 = {pp103[83]};
    Full_Adder FA_7595(s7595, c7595, in7595_1, in7595_2, pp101[85]);
    wire[0:0] s7596, in7596_1, in7596_2;
    wire c7596;
    assign in7596_1 = {pp105[81]};
    assign in7596_2 = {pp106[80]};
    Full_Adder FA_7596(s7596, c7596, in7596_1, in7596_2, pp104[82]);
    wire[0:0] s7597, in7597_1, in7597_2;
    wire c7597;
    assign in7597_1 = {pp108[78]};
    assign in7597_2 = {pp109[77]};
    Full_Adder FA_7597(s7597, c7597, in7597_1, in7597_2, pp107[79]);
    wire[0:0] s7598, in7598_1, in7598_2;
    wire c7598;
    assign in7598_1 = {pp111[75]};
    assign in7598_2 = {pp112[74]};
    Full_Adder FA_7598(s7598, c7598, in7598_1, in7598_2, pp110[76]);
    wire[0:0] s7599, in7599_1, in7599_2;
    wire c7599;
    assign in7599_1 = {pp114[72]};
    assign in7599_2 = {pp115[71]};
    Full_Adder FA_7599(s7599, c7599, in7599_1, in7599_2, pp113[73]);
    wire[0:0] s7600, in7600_1, in7600_2;
    wire c7600;
    assign in7600_1 = {pp117[69]};
    assign in7600_2 = {pp118[68]};
    Full_Adder FA_7600(s7600, c7600, in7600_1, in7600_2, pp116[70]);
    wire[0:0] s7601, in7601_1, in7601_2;
    wire c7601;
    assign in7601_1 = {pp120[66]};
    assign in7601_2 = {pp121[65]};
    Full_Adder FA_7601(s7601, c7601, in7601_1, in7601_2, pp119[67]);
    wire[0:0] s7602, in7602_1, in7602_2;
    wire c7602;
    assign in7602_1 = {pp123[63]};
    assign in7602_2 = {pp124[62]};
    Full_Adder FA_7602(s7602, c7602, in7602_1, in7602_2, pp122[64]);
    wire[0:0] s7603, in7603_1, in7603_2;
    wire c7603;
    assign in7603_1 = {pp126[60]};
    assign in7603_2 = {pp127[59]};
    Full_Adder FA_7603(s7603, c7603, in7603_1, in7603_2, pp125[61]);
    wire[0:0] s7604, in7604_1, in7604_2;
    wire c7604;
    assign in7604_1 = {c4881};
    assign in7604_2 = {c4882};
    Full_Adder FA_7604(s7604, c7604, in7604_1, in7604_2, c4880);
    wire[0:0] s7605, in7605_1, in7605_2;
    wire c7605;
    assign in7605_1 = {c4884};
    assign in7605_2 = {c4885};
    Full_Adder FA_7605(s7605, c7605, in7605_1, in7605_2, c4883);
    wire[0:0] s7606, in7606_1, in7606_2;
    wire c7606;
    assign in7606_1 = {c4887};
    assign in7606_2 = {c4888};
    Full_Adder FA_7606(s7606, c7606, in7606_1, in7606_2, c4886);
    wire[0:0] s7607, in7607_1, in7607_2;
    wire c7607;
    assign in7607_1 = {c4890};
    assign in7607_2 = {c4891};
    Full_Adder FA_7607(s7607, c7607, in7607_1, in7607_2, c4889);
    wire[0:0] s7608, in7608_1, in7608_2;
    wire c7608;
    assign in7608_1 = {s4893[0]};
    assign in7608_2 = {s4894[0]};
    Full_Adder FA_7608(s7608, c7608, in7608_1, in7608_2, c4892);
    wire[0:0] s7609, in7609_1, in7609_2;
    wire c7609;
    assign in7609_1 = {s4896[0]};
    assign in7609_2 = {s4897[0]};
    Full_Adder FA_7609(s7609, c7609, in7609_1, in7609_2, s4895[0]);
    wire[0:0] s7610, in7610_1, in7610_2;
    wire c7610;
    assign in7610_1 = {s4899[0]};
    assign in7610_2 = {s4900[0]};
    Full_Adder FA_7610(s7610, c7610, in7610_1, in7610_2, s4898[0]);
    wire[0:0] s7611, in7611_1, in7611_2;
    wire c7611;
    assign in7611_1 = {s4902[0]};
    assign in7611_2 = {s4903[0]};
    Full_Adder FA_7611(s7611, c7611, in7611_1, in7611_2, s4901[0]);
    wire[0:0] s7612, in7612_1, in7612_2;
    wire c7612;
    assign in7612_1 = {pp94[93]};
    assign in7612_2 = {pp95[92]};
    Full_Adder FA_7612(s7612, c7612, in7612_1, in7612_2, pp93[94]);
    wire[0:0] s7613, in7613_1, in7613_2;
    wire c7613;
    assign in7613_1 = {pp97[90]};
    assign in7613_2 = {pp98[89]};
    Full_Adder FA_7613(s7613, c7613, in7613_1, in7613_2, pp96[91]);
    wire[0:0] s7614, in7614_1, in7614_2;
    wire c7614;
    assign in7614_1 = {pp100[87]};
    assign in7614_2 = {pp101[86]};
    Full_Adder FA_7614(s7614, c7614, in7614_1, in7614_2, pp99[88]);
    wire[0:0] s7615, in7615_1, in7615_2;
    wire c7615;
    assign in7615_1 = {pp103[84]};
    assign in7615_2 = {pp104[83]};
    Full_Adder FA_7615(s7615, c7615, in7615_1, in7615_2, pp102[85]);
    wire[0:0] s7616, in7616_1, in7616_2;
    wire c7616;
    assign in7616_1 = {pp106[81]};
    assign in7616_2 = {pp107[80]};
    Full_Adder FA_7616(s7616, c7616, in7616_1, in7616_2, pp105[82]);
    wire[0:0] s7617, in7617_1, in7617_2;
    wire c7617;
    assign in7617_1 = {pp109[78]};
    assign in7617_2 = {pp110[77]};
    Full_Adder FA_7617(s7617, c7617, in7617_1, in7617_2, pp108[79]);
    wire[0:0] s7618, in7618_1, in7618_2;
    wire c7618;
    assign in7618_1 = {pp112[75]};
    assign in7618_2 = {pp113[74]};
    Full_Adder FA_7618(s7618, c7618, in7618_1, in7618_2, pp111[76]);
    wire[0:0] s7619, in7619_1, in7619_2;
    wire c7619;
    assign in7619_1 = {pp115[72]};
    assign in7619_2 = {pp116[71]};
    Full_Adder FA_7619(s7619, c7619, in7619_1, in7619_2, pp114[73]);
    wire[0:0] s7620, in7620_1, in7620_2;
    wire c7620;
    assign in7620_1 = {pp118[69]};
    assign in7620_2 = {pp119[68]};
    Full_Adder FA_7620(s7620, c7620, in7620_1, in7620_2, pp117[70]);
    wire[0:0] s7621, in7621_1, in7621_2;
    wire c7621;
    assign in7621_1 = {pp121[66]};
    assign in7621_2 = {pp122[65]};
    Full_Adder FA_7621(s7621, c7621, in7621_1, in7621_2, pp120[67]);
    wire[0:0] s7622, in7622_1, in7622_2;
    wire c7622;
    assign in7622_1 = {pp124[63]};
    assign in7622_2 = {pp125[62]};
    Full_Adder FA_7622(s7622, c7622, in7622_1, in7622_2, pp123[64]);
    wire[0:0] s7623, in7623_1, in7623_2;
    wire c7623;
    assign in7623_1 = {pp127[60]};
    assign in7623_2 = {c4893};
    Full_Adder FA_7623(s7623, c7623, in7623_1, in7623_2, pp126[61]);
    wire[0:0] s7624, in7624_1, in7624_2;
    wire c7624;
    assign in7624_1 = {c4895};
    assign in7624_2 = {c4896};
    Full_Adder FA_7624(s7624, c7624, in7624_1, in7624_2, c4894);
    wire[0:0] s7625, in7625_1, in7625_2;
    wire c7625;
    assign in7625_1 = {c4898};
    assign in7625_2 = {c4899};
    Full_Adder FA_7625(s7625, c7625, in7625_1, in7625_2, c4897);
    wire[0:0] s7626, in7626_1, in7626_2;
    wire c7626;
    assign in7626_1 = {c4901};
    assign in7626_2 = {c4902};
    Full_Adder FA_7626(s7626, c7626, in7626_1, in7626_2, c4900);
    wire[0:0] s7627, in7627_1, in7627_2;
    wire c7627;
    assign in7627_1 = {c4904};
    assign in7627_2 = {s4905[0]};
    Full_Adder FA_7627(s7627, c7627, in7627_1, in7627_2, c4903);
    wire[0:0] s7628, in7628_1, in7628_2;
    wire c7628;
    assign in7628_1 = {s4907[0]};
    assign in7628_2 = {s4908[0]};
    Full_Adder FA_7628(s7628, c7628, in7628_1, in7628_2, s4906[0]);
    wire[0:0] s7629, in7629_1, in7629_2;
    wire c7629;
    assign in7629_1 = {s4910[0]};
    assign in7629_2 = {s4911[0]};
    Full_Adder FA_7629(s7629, c7629, in7629_1, in7629_2, s4909[0]);
    wire[0:0] s7630, in7630_1, in7630_2;
    wire c7630;
    assign in7630_1 = {s4913[0]};
    assign in7630_2 = {s4914[0]};
    Full_Adder FA_7630(s7630, c7630, in7630_1, in7630_2, s4912[0]);
    wire[0:0] s7631, in7631_1, in7631_2;
    wire c7631;
    assign in7631_1 = {pp92[96]};
    assign in7631_2 = {pp93[95]};
    Full_Adder FA_7631(s7631, c7631, in7631_1, in7631_2, pp91[97]);
    wire[0:0] s7632, in7632_1, in7632_2;
    wire c7632;
    assign in7632_1 = {pp95[93]};
    assign in7632_2 = {pp96[92]};
    Full_Adder FA_7632(s7632, c7632, in7632_1, in7632_2, pp94[94]);
    wire[0:0] s7633, in7633_1, in7633_2;
    wire c7633;
    assign in7633_1 = {pp98[90]};
    assign in7633_2 = {pp99[89]};
    Full_Adder FA_7633(s7633, c7633, in7633_1, in7633_2, pp97[91]);
    wire[0:0] s7634, in7634_1, in7634_2;
    wire c7634;
    assign in7634_1 = {pp101[87]};
    assign in7634_2 = {pp102[86]};
    Full_Adder FA_7634(s7634, c7634, in7634_1, in7634_2, pp100[88]);
    wire[0:0] s7635, in7635_1, in7635_2;
    wire c7635;
    assign in7635_1 = {pp104[84]};
    assign in7635_2 = {pp105[83]};
    Full_Adder FA_7635(s7635, c7635, in7635_1, in7635_2, pp103[85]);
    wire[0:0] s7636, in7636_1, in7636_2;
    wire c7636;
    assign in7636_1 = {pp107[81]};
    assign in7636_2 = {pp108[80]};
    Full_Adder FA_7636(s7636, c7636, in7636_1, in7636_2, pp106[82]);
    wire[0:0] s7637, in7637_1, in7637_2;
    wire c7637;
    assign in7637_1 = {pp110[78]};
    assign in7637_2 = {pp111[77]};
    Full_Adder FA_7637(s7637, c7637, in7637_1, in7637_2, pp109[79]);
    wire[0:0] s7638, in7638_1, in7638_2;
    wire c7638;
    assign in7638_1 = {pp113[75]};
    assign in7638_2 = {pp114[74]};
    Full_Adder FA_7638(s7638, c7638, in7638_1, in7638_2, pp112[76]);
    wire[0:0] s7639, in7639_1, in7639_2;
    wire c7639;
    assign in7639_1 = {pp116[72]};
    assign in7639_2 = {pp117[71]};
    Full_Adder FA_7639(s7639, c7639, in7639_1, in7639_2, pp115[73]);
    wire[0:0] s7640, in7640_1, in7640_2;
    wire c7640;
    assign in7640_1 = {pp119[69]};
    assign in7640_2 = {pp120[68]};
    Full_Adder FA_7640(s7640, c7640, in7640_1, in7640_2, pp118[70]);
    wire[0:0] s7641, in7641_1, in7641_2;
    wire c7641;
    assign in7641_1 = {pp122[66]};
    assign in7641_2 = {pp123[65]};
    Full_Adder FA_7641(s7641, c7641, in7641_1, in7641_2, pp121[67]);
    wire[0:0] s7642, in7642_1, in7642_2;
    wire c7642;
    assign in7642_1 = {pp125[63]};
    assign in7642_2 = {pp126[62]};
    Full_Adder FA_7642(s7642, c7642, in7642_1, in7642_2, pp124[64]);
    wire[0:0] s7643, in7643_1, in7643_2;
    wire c7643;
    assign in7643_1 = {c4905};
    assign in7643_2 = {c4906};
    Full_Adder FA_7643(s7643, c7643, in7643_1, in7643_2, pp127[61]);
    wire[0:0] s7644, in7644_1, in7644_2;
    wire c7644;
    assign in7644_1 = {c4908};
    assign in7644_2 = {c4909};
    Full_Adder FA_7644(s7644, c7644, in7644_1, in7644_2, c4907);
    wire[0:0] s7645, in7645_1, in7645_2;
    wire c7645;
    assign in7645_1 = {c4911};
    assign in7645_2 = {c4912};
    Full_Adder FA_7645(s7645, c7645, in7645_1, in7645_2, c4910);
    wire[0:0] s7646, in7646_1, in7646_2;
    wire c7646;
    assign in7646_1 = {c4914};
    assign in7646_2 = {c4915};
    Full_Adder FA_7646(s7646, c7646, in7646_1, in7646_2, c4913);
    wire[0:0] s7647, in7647_1, in7647_2;
    wire c7647;
    assign in7647_1 = {s4917[0]};
    assign in7647_2 = {s4918[0]};
    Full_Adder FA_7647(s7647, c7647, in7647_1, in7647_2, s4916[0]);
    wire[0:0] s7648, in7648_1, in7648_2;
    wire c7648;
    assign in7648_1 = {s4920[0]};
    assign in7648_2 = {s4921[0]};
    Full_Adder FA_7648(s7648, c7648, in7648_1, in7648_2, s4919[0]);
    wire[0:0] s7649, in7649_1, in7649_2;
    wire c7649;
    assign in7649_1 = {s4923[0]};
    assign in7649_2 = {s4924[0]};
    Full_Adder FA_7649(s7649, c7649, in7649_1, in7649_2, s4922[0]);
    wire[0:0] s7650, in7650_1, in7650_2;
    wire c7650;
    assign in7650_1 = {pp90[99]};
    assign in7650_2 = {pp91[98]};
    Full_Adder FA_7650(s7650, c7650, in7650_1, in7650_2, pp89[100]);
    wire[0:0] s7651, in7651_1, in7651_2;
    wire c7651;
    assign in7651_1 = {pp93[96]};
    assign in7651_2 = {pp94[95]};
    Full_Adder FA_7651(s7651, c7651, in7651_1, in7651_2, pp92[97]);
    wire[0:0] s7652, in7652_1, in7652_2;
    wire c7652;
    assign in7652_1 = {pp96[93]};
    assign in7652_2 = {pp97[92]};
    Full_Adder FA_7652(s7652, c7652, in7652_1, in7652_2, pp95[94]);
    wire[0:0] s7653, in7653_1, in7653_2;
    wire c7653;
    assign in7653_1 = {pp99[90]};
    assign in7653_2 = {pp100[89]};
    Full_Adder FA_7653(s7653, c7653, in7653_1, in7653_2, pp98[91]);
    wire[0:0] s7654, in7654_1, in7654_2;
    wire c7654;
    assign in7654_1 = {pp102[87]};
    assign in7654_2 = {pp103[86]};
    Full_Adder FA_7654(s7654, c7654, in7654_1, in7654_2, pp101[88]);
    wire[0:0] s7655, in7655_1, in7655_2;
    wire c7655;
    assign in7655_1 = {pp105[84]};
    assign in7655_2 = {pp106[83]};
    Full_Adder FA_7655(s7655, c7655, in7655_1, in7655_2, pp104[85]);
    wire[0:0] s7656, in7656_1, in7656_2;
    wire c7656;
    assign in7656_1 = {pp108[81]};
    assign in7656_2 = {pp109[80]};
    Full_Adder FA_7656(s7656, c7656, in7656_1, in7656_2, pp107[82]);
    wire[0:0] s7657, in7657_1, in7657_2;
    wire c7657;
    assign in7657_1 = {pp111[78]};
    assign in7657_2 = {pp112[77]};
    Full_Adder FA_7657(s7657, c7657, in7657_1, in7657_2, pp110[79]);
    wire[0:0] s7658, in7658_1, in7658_2;
    wire c7658;
    assign in7658_1 = {pp114[75]};
    assign in7658_2 = {pp115[74]};
    Full_Adder FA_7658(s7658, c7658, in7658_1, in7658_2, pp113[76]);
    wire[0:0] s7659, in7659_1, in7659_2;
    wire c7659;
    assign in7659_1 = {pp117[72]};
    assign in7659_2 = {pp118[71]};
    Full_Adder FA_7659(s7659, c7659, in7659_1, in7659_2, pp116[73]);
    wire[0:0] s7660, in7660_1, in7660_2;
    wire c7660;
    assign in7660_1 = {pp120[69]};
    assign in7660_2 = {pp121[68]};
    Full_Adder FA_7660(s7660, c7660, in7660_1, in7660_2, pp119[70]);
    wire[0:0] s7661, in7661_1, in7661_2;
    wire c7661;
    assign in7661_1 = {pp123[66]};
    assign in7661_2 = {pp124[65]};
    Full_Adder FA_7661(s7661, c7661, in7661_1, in7661_2, pp122[67]);
    wire[0:0] s7662, in7662_1, in7662_2;
    wire c7662;
    assign in7662_1 = {pp126[63]};
    assign in7662_2 = {pp127[62]};
    Full_Adder FA_7662(s7662, c7662, in7662_1, in7662_2, pp125[64]);
    wire[0:0] s7663, in7663_1, in7663_2;
    wire c7663;
    assign in7663_1 = {c4917};
    assign in7663_2 = {c4918};
    Full_Adder FA_7663(s7663, c7663, in7663_1, in7663_2, c4916);
    wire[0:0] s7664, in7664_1, in7664_2;
    wire c7664;
    assign in7664_1 = {c4920};
    assign in7664_2 = {c4921};
    Full_Adder FA_7664(s7664, c7664, in7664_1, in7664_2, c4919);
    wire[0:0] s7665, in7665_1, in7665_2;
    wire c7665;
    assign in7665_1 = {c4923};
    assign in7665_2 = {c4924};
    Full_Adder FA_7665(s7665, c7665, in7665_1, in7665_2, c4922);
    wire[0:0] s7666, in7666_1, in7666_2;
    wire c7666;
    assign in7666_1 = {s4926[0]};
    assign in7666_2 = {s4927[0]};
    Full_Adder FA_7666(s7666, c7666, in7666_1, in7666_2, c4925);
    wire[0:0] s7667, in7667_1, in7667_2;
    wire c7667;
    assign in7667_1 = {s4929[0]};
    assign in7667_2 = {s4930[0]};
    Full_Adder FA_7667(s7667, c7667, in7667_1, in7667_2, s4928[0]);
    wire[0:0] s7668, in7668_1, in7668_2;
    wire c7668;
    assign in7668_1 = {s4932[0]};
    assign in7668_2 = {s4933[0]};
    Full_Adder FA_7668(s7668, c7668, in7668_1, in7668_2, s4931[0]);
    wire[0:0] s7669, in7669_1, in7669_2;
    wire c7669;
    assign in7669_1 = {pp88[102]};
    assign in7669_2 = {pp89[101]};
    Full_Adder FA_7669(s7669, c7669, in7669_1, in7669_2, pp87[103]);
    wire[0:0] s7670, in7670_1, in7670_2;
    wire c7670;
    assign in7670_1 = {pp91[99]};
    assign in7670_2 = {pp92[98]};
    Full_Adder FA_7670(s7670, c7670, in7670_1, in7670_2, pp90[100]);
    wire[0:0] s7671, in7671_1, in7671_2;
    wire c7671;
    assign in7671_1 = {pp94[96]};
    assign in7671_2 = {pp95[95]};
    Full_Adder FA_7671(s7671, c7671, in7671_1, in7671_2, pp93[97]);
    wire[0:0] s7672, in7672_1, in7672_2;
    wire c7672;
    assign in7672_1 = {pp97[93]};
    assign in7672_2 = {pp98[92]};
    Full_Adder FA_7672(s7672, c7672, in7672_1, in7672_2, pp96[94]);
    wire[0:0] s7673, in7673_1, in7673_2;
    wire c7673;
    assign in7673_1 = {pp100[90]};
    assign in7673_2 = {pp101[89]};
    Full_Adder FA_7673(s7673, c7673, in7673_1, in7673_2, pp99[91]);
    wire[0:0] s7674, in7674_1, in7674_2;
    wire c7674;
    assign in7674_1 = {pp103[87]};
    assign in7674_2 = {pp104[86]};
    Full_Adder FA_7674(s7674, c7674, in7674_1, in7674_2, pp102[88]);
    wire[0:0] s7675, in7675_1, in7675_2;
    wire c7675;
    assign in7675_1 = {pp106[84]};
    assign in7675_2 = {pp107[83]};
    Full_Adder FA_7675(s7675, c7675, in7675_1, in7675_2, pp105[85]);
    wire[0:0] s7676, in7676_1, in7676_2;
    wire c7676;
    assign in7676_1 = {pp109[81]};
    assign in7676_2 = {pp110[80]};
    Full_Adder FA_7676(s7676, c7676, in7676_1, in7676_2, pp108[82]);
    wire[0:0] s7677, in7677_1, in7677_2;
    wire c7677;
    assign in7677_1 = {pp112[78]};
    assign in7677_2 = {pp113[77]};
    Full_Adder FA_7677(s7677, c7677, in7677_1, in7677_2, pp111[79]);
    wire[0:0] s7678, in7678_1, in7678_2;
    wire c7678;
    assign in7678_1 = {pp115[75]};
    assign in7678_2 = {pp116[74]};
    Full_Adder FA_7678(s7678, c7678, in7678_1, in7678_2, pp114[76]);
    wire[0:0] s7679, in7679_1, in7679_2;
    wire c7679;
    assign in7679_1 = {pp118[72]};
    assign in7679_2 = {pp119[71]};
    Full_Adder FA_7679(s7679, c7679, in7679_1, in7679_2, pp117[73]);
    wire[0:0] s7680, in7680_1, in7680_2;
    wire c7680;
    assign in7680_1 = {pp121[69]};
    assign in7680_2 = {pp122[68]};
    Full_Adder FA_7680(s7680, c7680, in7680_1, in7680_2, pp120[70]);
    wire[0:0] s7681, in7681_1, in7681_2;
    wire c7681;
    assign in7681_1 = {pp124[66]};
    assign in7681_2 = {pp125[65]};
    Full_Adder FA_7681(s7681, c7681, in7681_1, in7681_2, pp123[67]);
    wire[0:0] s7682, in7682_1, in7682_2;
    wire c7682;
    assign in7682_1 = {pp127[63]};
    assign in7682_2 = {c4926};
    Full_Adder FA_7682(s7682, c7682, in7682_1, in7682_2, pp126[64]);
    wire[0:0] s7683, in7683_1, in7683_2;
    wire c7683;
    assign in7683_1 = {c4928};
    assign in7683_2 = {c4929};
    Full_Adder FA_7683(s7683, c7683, in7683_1, in7683_2, c4927);
    wire[0:0] s7684, in7684_1, in7684_2;
    wire c7684;
    assign in7684_1 = {c4931};
    assign in7684_2 = {c4932};
    Full_Adder FA_7684(s7684, c7684, in7684_1, in7684_2, c4930);
    wire[0:0] s7685, in7685_1, in7685_2;
    wire c7685;
    assign in7685_1 = {c4934};
    assign in7685_2 = {s4935[0]};
    Full_Adder FA_7685(s7685, c7685, in7685_1, in7685_2, c4933);
    wire[0:0] s7686, in7686_1, in7686_2;
    wire c7686;
    assign in7686_1 = {s4937[0]};
    assign in7686_2 = {s4938[0]};
    Full_Adder FA_7686(s7686, c7686, in7686_1, in7686_2, s4936[0]);
    wire[0:0] s7687, in7687_1, in7687_2;
    wire c7687;
    assign in7687_1 = {s4940[0]};
    assign in7687_2 = {s4941[0]};
    Full_Adder FA_7687(s7687, c7687, in7687_1, in7687_2, s4939[0]);
    wire[0:0] s7688, in7688_1, in7688_2;
    wire c7688;
    assign in7688_1 = {pp86[105]};
    assign in7688_2 = {pp87[104]};
    Full_Adder FA_7688(s7688, c7688, in7688_1, in7688_2, pp85[106]);
    wire[0:0] s7689, in7689_1, in7689_2;
    wire c7689;
    assign in7689_1 = {pp89[102]};
    assign in7689_2 = {pp90[101]};
    Full_Adder FA_7689(s7689, c7689, in7689_1, in7689_2, pp88[103]);
    wire[0:0] s7690, in7690_1, in7690_2;
    wire c7690;
    assign in7690_1 = {pp92[99]};
    assign in7690_2 = {pp93[98]};
    Full_Adder FA_7690(s7690, c7690, in7690_1, in7690_2, pp91[100]);
    wire[0:0] s7691, in7691_1, in7691_2;
    wire c7691;
    assign in7691_1 = {pp95[96]};
    assign in7691_2 = {pp96[95]};
    Full_Adder FA_7691(s7691, c7691, in7691_1, in7691_2, pp94[97]);
    wire[0:0] s7692, in7692_1, in7692_2;
    wire c7692;
    assign in7692_1 = {pp98[93]};
    assign in7692_2 = {pp99[92]};
    Full_Adder FA_7692(s7692, c7692, in7692_1, in7692_2, pp97[94]);
    wire[0:0] s7693, in7693_1, in7693_2;
    wire c7693;
    assign in7693_1 = {pp101[90]};
    assign in7693_2 = {pp102[89]};
    Full_Adder FA_7693(s7693, c7693, in7693_1, in7693_2, pp100[91]);
    wire[0:0] s7694, in7694_1, in7694_2;
    wire c7694;
    assign in7694_1 = {pp104[87]};
    assign in7694_2 = {pp105[86]};
    Full_Adder FA_7694(s7694, c7694, in7694_1, in7694_2, pp103[88]);
    wire[0:0] s7695, in7695_1, in7695_2;
    wire c7695;
    assign in7695_1 = {pp107[84]};
    assign in7695_2 = {pp108[83]};
    Full_Adder FA_7695(s7695, c7695, in7695_1, in7695_2, pp106[85]);
    wire[0:0] s7696, in7696_1, in7696_2;
    wire c7696;
    assign in7696_1 = {pp110[81]};
    assign in7696_2 = {pp111[80]};
    Full_Adder FA_7696(s7696, c7696, in7696_1, in7696_2, pp109[82]);
    wire[0:0] s7697, in7697_1, in7697_2;
    wire c7697;
    assign in7697_1 = {pp113[78]};
    assign in7697_2 = {pp114[77]};
    Full_Adder FA_7697(s7697, c7697, in7697_1, in7697_2, pp112[79]);
    wire[0:0] s7698, in7698_1, in7698_2;
    wire c7698;
    assign in7698_1 = {pp116[75]};
    assign in7698_2 = {pp117[74]};
    Full_Adder FA_7698(s7698, c7698, in7698_1, in7698_2, pp115[76]);
    wire[0:0] s7699, in7699_1, in7699_2;
    wire c7699;
    assign in7699_1 = {pp119[72]};
    assign in7699_2 = {pp120[71]};
    Full_Adder FA_7699(s7699, c7699, in7699_1, in7699_2, pp118[73]);
    wire[0:0] s7700, in7700_1, in7700_2;
    wire c7700;
    assign in7700_1 = {pp122[69]};
    assign in7700_2 = {pp123[68]};
    Full_Adder FA_7700(s7700, c7700, in7700_1, in7700_2, pp121[70]);
    wire[0:0] s7701, in7701_1, in7701_2;
    wire c7701;
    assign in7701_1 = {pp125[66]};
    assign in7701_2 = {pp126[65]};
    Full_Adder FA_7701(s7701, c7701, in7701_1, in7701_2, pp124[67]);
    wire[0:0] s7702, in7702_1, in7702_2;
    wire c7702;
    assign in7702_1 = {c4935};
    assign in7702_2 = {c4936};
    Full_Adder FA_7702(s7702, c7702, in7702_1, in7702_2, pp127[64]);
    wire[0:0] s7703, in7703_1, in7703_2;
    wire c7703;
    assign in7703_1 = {c4938};
    assign in7703_2 = {c4939};
    Full_Adder FA_7703(s7703, c7703, in7703_1, in7703_2, c4937);
    wire[0:0] s7704, in7704_1, in7704_2;
    wire c7704;
    assign in7704_1 = {c4941};
    assign in7704_2 = {c4942};
    Full_Adder FA_7704(s7704, c7704, in7704_1, in7704_2, c4940);
    wire[0:0] s7705, in7705_1, in7705_2;
    wire c7705;
    assign in7705_1 = {s4944[0]};
    assign in7705_2 = {s4945[0]};
    Full_Adder FA_7705(s7705, c7705, in7705_1, in7705_2, s4943[0]);
    wire[0:0] s7706, in7706_1, in7706_2;
    wire c7706;
    assign in7706_1 = {s4947[0]};
    assign in7706_2 = {s4948[0]};
    Full_Adder FA_7706(s7706, c7706, in7706_1, in7706_2, s4946[0]);
    wire[0:0] s7707, in7707_1, in7707_2;
    wire c7707;
    assign in7707_1 = {pp84[108]};
    assign in7707_2 = {pp85[107]};
    Full_Adder FA_7707(s7707, c7707, in7707_1, in7707_2, pp83[109]);
    wire[0:0] s7708, in7708_1, in7708_2;
    wire c7708;
    assign in7708_1 = {pp87[105]};
    assign in7708_2 = {pp88[104]};
    Full_Adder FA_7708(s7708, c7708, in7708_1, in7708_2, pp86[106]);
    wire[0:0] s7709, in7709_1, in7709_2;
    wire c7709;
    assign in7709_1 = {pp90[102]};
    assign in7709_2 = {pp91[101]};
    Full_Adder FA_7709(s7709, c7709, in7709_1, in7709_2, pp89[103]);
    wire[0:0] s7710, in7710_1, in7710_2;
    wire c7710;
    assign in7710_1 = {pp93[99]};
    assign in7710_2 = {pp94[98]};
    Full_Adder FA_7710(s7710, c7710, in7710_1, in7710_2, pp92[100]);
    wire[0:0] s7711, in7711_1, in7711_2;
    wire c7711;
    assign in7711_1 = {pp96[96]};
    assign in7711_2 = {pp97[95]};
    Full_Adder FA_7711(s7711, c7711, in7711_1, in7711_2, pp95[97]);
    wire[0:0] s7712, in7712_1, in7712_2;
    wire c7712;
    assign in7712_1 = {pp99[93]};
    assign in7712_2 = {pp100[92]};
    Full_Adder FA_7712(s7712, c7712, in7712_1, in7712_2, pp98[94]);
    wire[0:0] s7713, in7713_1, in7713_2;
    wire c7713;
    assign in7713_1 = {pp102[90]};
    assign in7713_2 = {pp103[89]};
    Full_Adder FA_7713(s7713, c7713, in7713_1, in7713_2, pp101[91]);
    wire[0:0] s7714, in7714_1, in7714_2;
    wire c7714;
    assign in7714_1 = {pp105[87]};
    assign in7714_2 = {pp106[86]};
    Full_Adder FA_7714(s7714, c7714, in7714_1, in7714_2, pp104[88]);
    wire[0:0] s7715, in7715_1, in7715_2;
    wire c7715;
    assign in7715_1 = {pp108[84]};
    assign in7715_2 = {pp109[83]};
    Full_Adder FA_7715(s7715, c7715, in7715_1, in7715_2, pp107[85]);
    wire[0:0] s7716, in7716_1, in7716_2;
    wire c7716;
    assign in7716_1 = {pp111[81]};
    assign in7716_2 = {pp112[80]};
    Full_Adder FA_7716(s7716, c7716, in7716_1, in7716_2, pp110[82]);
    wire[0:0] s7717, in7717_1, in7717_2;
    wire c7717;
    assign in7717_1 = {pp114[78]};
    assign in7717_2 = {pp115[77]};
    Full_Adder FA_7717(s7717, c7717, in7717_1, in7717_2, pp113[79]);
    wire[0:0] s7718, in7718_1, in7718_2;
    wire c7718;
    assign in7718_1 = {pp117[75]};
    assign in7718_2 = {pp118[74]};
    Full_Adder FA_7718(s7718, c7718, in7718_1, in7718_2, pp116[76]);
    wire[0:0] s7719, in7719_1, in7719_2;
    wire c7719;
    assign in7719_1 = {pp120[72]};
    assign in7719_2 = {pp121[71]};
    Full_Adder FA_7719(s7719, c7719, in7719_1, in7719_2, pp119[73]);
    wire[0:0] s7720, in7720_1, in7720_2;
    wire c7720;
    assign in7720_1 = {pp123[69]};
    assign in7720_2 = {pp124[68]};
    Full_Adder FA_7720(s7720, c7720, in7720_1, in7720_2, pp122[70]);
    wire[0:0] s7721, in7721_1, in7721_2;
    wire c7721;
    assign in7721_1 = {pp126[66]};
    assign in7721_2 = {pp127[65]};
    Full_Adder FA_7721(s7721, c7721, in7721_1, in7721_2, pp125[67]);
    wire[0:0] s7722, in7722_1, in7722_2;
    wire c7722;
    assign in7722_1 = {c4944};
    assign in7722_2 = {c4945};
    Full_Adder FA_7722(s7722, c7722, in7722_1, in7722_2, c4943);
    wire[0:0] s7723, in7723_1, in7723_2;
    wire c7723;
    assign in7723_1 = {c4947};
    assign in7723_2 = {c4948};
    Full_Adder FA_7723(s7723, c7723, in7723_1, in7723_2, c4946);
    wire[0:0] s7724, in7724_1, in7724_2;
    wire c7724;
    assign in7724_1 = {s4950[0]};
    assign in7724_2 = {s4951[0]};
    Full_Adder FA_7724(s7724, c7724, in7724_1, in7724_2, c4949);
    wire[0:0] s7725, in7725_1, in7725_2;
    wire c7725;
    assign in7725_1 = {s4953[0]};
    assign in7725_2 = {s4954[0]};
    Full_Adder FA_7725(s7725, c7725, in7725_1, in7725_2, s4952[0]);
    wire[0:0] s7726, in7726_1, in7726_2;
    wire c7726;
    assign in7726_1 = {pp82[111]};
    assign in7726_2 = {pp83[110]};
    Full_Adder FA_7726(s7726, c7726, in7726_1, in7726_2, pp81[112]);
    wire[0:0] s7727, in7727_1, in7727_2;
    wire c7727;
    assign in7727_1 = {pp85[108]};
    assign in7727_2 = {pp86[107]};
    Full_Adder FA_7727(s7727, c7727, in7727_1, in7727_2, pp84[109]);
    wire[0:0] s7728, in7728_1, in7728_2;
    wire c7728;
    assign in7728_1 = {pp88[105]};
    assign in7728_2 = {pp89[104]};
    Full_Adder FA_7728(s7728, c7728, in7728_1, in7728_2, pp87[106]);
    wire[0:0] s7729, in7729_1, in7729_2;
    wire c7729;
    assign in7729_1 = {pp91[102]};
    assign in7729_2 = {pp92[101]};
    Full_Adder FA_7729(s7729, c7729, in7729_1, in7729_2, pp90[103]);
    wire[0:0] s7730, in7730_1, in7730_2;
    wire c7730;
    assign in7730_1 = {pp94[99]};
    assign in7730_2 = {pp95[98]};
    Full_Adder FA_7730(s7730, c7730, in7730_1, in7730_2, pp93[100]);
    wire[0:0] s7731, in7731_1, in7731_2;
    wire c7731;
    assign in7731_1 = {pp97[96]};
    assign in7731_2 = {pp98[95]};
    Full_Adder FA_7731(s7731, c7731, in7731_1, in7731_2, pp96[97]);
    wire[0:0] s7732, in7732_1, in7732_2;
    wire c7732;
    assign in7732_1 = {pp100[93]};
    assign in7732_2 = {pp101[92]};
    Full_Adder FA_7732(s7732, c7732, in7732_1, in7732_2, pp99[94]);
    wire[0:0] s7733, in7733_1, in7733_2;
    wire c7733;
    assign in7733_1 = {pp103[90]};
    assign in7733_2 = {pp104[89]};
    Full_Adder FA_7733(s7733, c7733, in7733_1, in7733_2, pp102[91]);
    wire[0:0] s7734, in7734_1, in7734_2;
    wire c7734;
    assign in7734_1 = {pp106[87]};
    assign in7734_2 = {pp107[86]};
    Full_Adder FA_7734(s7734, c7734, in7734_1, in7734_2, pp105[88]);
    wire[0:0] s7735, in7735_1, in7735_2;
    wire c7735;
    assign in7735_1 = {pp109[84]};
    assign in7735_2 = {pp110[83]};
    Full_Adder FA_7735(s7735, c7735, in7735_1, in7735_2, pp108[85]);
    wire[0:0] s7736, in7736_1, in7736_2;
    wire c7736;
    assign in7736_1 = {pp112[81]};
    assign in7736_2 = {pp113[80]};
    Full_Adder FA_7736(s7736, c7736, in7736_1, in7736_2, pp111[82]);
    wire[0:0] s7737, in7737_1, in7737_2;
    wire c7737;
    assign in7737_1 = {pp115[78]};
    assign in7737_2 = {pp116[77]};
    Full_Adder FA_7737(s7737, c7737, in7737_1, in7737_2, pp114[79]);
    wire[0:0] s7738, in7738_1, in7738_2;
    wire c7738;
    assign in7738_1 = {pp118[75]};
    assign in7738_2 = {pp119[74]};
    Full_Adder FA_7738(s7738, c7738, in7738_1, in7738_2, pp117[76]);
    wire[0:0] s7739, in7739_1, in7739_2;
    wire c7739;
    assign in7739_1 = {pp121[72]};
    assign in7739_2 = {pp122[71]};
    Full_Adder FA_7739(s7739, c7739, in7739_1, in7739_2, pp120[73]);
    wire[0:0] s7740, in7740_1, in7740_2;
    wire c7740;
    assign in7740_1 = {pp124[69]};
    assign in7740_2 = {pp125[68]};
    Full_Adder FA_7740(s7740, c7740, in7740_1, in7740_2, pp123[70]);
    wire[0:0] s7741, in7741_1, in7741_2;
    wire c7741;
    assign in7741_1 = {pp127[66]};
    assign in7741_2 = {c4950};
    Full_Adder FA_7741(s7741, c7741, in7741_1, in7741_2, pp126[67]);
    wire[0:0] s7742, in7742_1, in7742_2;
    wire c7742;
    assign in7742_1 = {c4952};
    assign in7742_2 = {c4953};
    Full_Adder FA_7742(s7742, c7742, in7742_1, in7742_2, c4951);
    wire[0:0] s7743, in7743_1, in7743_2;
    wire c7743;
    assign in7743_1 = {c4955};
    assign in7743_2 = {s4956[0]};
    Full_Adder FA_7743(s7743, c7743, in7743_1, in7743_2, c4954);
    wire[0:0] s7744, in7744_1, in7744_2;
    wire c7744;
    assign in7744_1 = {s4958[0]};
    assign in7744_2 = {s4959[0]};
    Full_Adder FA_7744(s7744, c7744, in7744_1, in7744_2, s4957[0]);
    wire[0:0] s7745, in7745_1, in7745_2;
    wire c7745;
    assign in7745_1 = {pp80[114]};
    assign in7745_2 = {pp81[113]};
    Full_Adder FA_7745(s7745, c7745, in7745_1, in7745_2, pp79[115]);
    wire[0:0] s7746, in7746_1, in7746_2;
    wire c7746;
    assign in7746_1 = {pp83[111]};
    assign in7746_2 = {pp84[110]};
    Full_Adder FA_7746(s7746, c7746, in7746_1, in7746_2, pp82[112]);
    wire[0:0] s7747, in7747_1, in7747_2;
    wire c7747;
    assign in7747_1 = {pp86[108]};
    assign in7747_2 = {pp87[107]};
    Full_Adder FA_7747(s7747, c7747, in7747_1, in7747_2, pp85[109]);
    wire[0:0] s7748, in7748_1, in7748_2;
    wire c7748;
    assign in7748_1 = {pp89[105]};
    assign in7748_2 = {pp90[104]};
    Full_Adder FA_7748(s7748, c7748, in7748_1, in7748_2, pp88[106]);
    wire[0:0] s7749, in7749_1, in7749_2;
    wire c7749;
    assign in7749_1 = {pp92[102]};
    assign in7749_2 = {pp93[101]};
    Full_Adder FA_7749(s7749, c7749, in7749_1, in7749_2, pp91[103]);
    wire[0:0] s7750, in7750_1, in7750_2;
    wire c7750;
    assign in7750_1 = {pp95[99]};
    assign in7750_2 = {pp96[98]};
    Full_Adder FA_7750(s7750, c7750, in7750_1, in7750_2, pp94[100]);
    wire[0:0] s7751, in7751_1, in7751_2;
    wire c7751;
    assign in7751_1 = {pp98[96]};
    assign in7751_2 = {pp99[95]};
    Full_Adder FA_7751(s7751, c7751, in7751_1, in7751_2, pp97[97]);
    wire[0:0] s7752, in7752_1, in7752_2;
    wire c7752;
    assign in7752_1 = {pp101[93]};
    assign in7752_2 = {pp102[92]};
    Full_Adder FA_7752(s7752, c7752, in7752_1, in7752_2, pp100[94]);
    wire[0:0] s7753, in7753_1, in7753_2;
    wire c7753;
    assign in7753_1 = {pp104[90]};
    assign in7753_2 = {pp105[89]};
    Full_Adder FA_7753(s7753, c7753, in7753_1, in7753_2, pp103[91]);
    wire[0:0] s7754, in7754_1, in7754_2;
    wire c7754;
    assign in7754_1 = {pp107[87]};
    assign in7754_2 = {pp108[86]};
    Full_Adder FA_7754(s7754, c7754, in7754_1, in7754_2, pp106[88]);
    wire[0:0] s7755, in7755_1, in7755_2;
    wire c7755;
    assign in7755_1 = {pp110[84]};
    assign in7755_2 = {pp111[83]};
    Full_Adder FA_7755(s7755, c7755, in7755_1, in7755_2, pp109[85]);
    wire[0:0] s7756, in7756_1, in7756_2;
    wire c7756;
    assign in7756_1 = {pp113[81]};
    assign in7756_2 = {pp114[80]};
    Full_Adder FA_7756(s7756, c7756, in7756_1, in7756_2, pp112[82]);
    wire[0:0] s7757, in7757_1, in7757_2;
    wire c7757;
    assign in7757_1 = {pp116[78]};
    assign in7757_2 = {pp117[77]};
    Full_Adder FA_7757(s7757, c7757, in7757_1, in7757_2, pp115[79]);
    wire[0:0] s7758, in7758_1, in7758_2;
    wire c7758;
    assign in7758_1 = {pp119[75]};
    assign in7758_2 = {pp120[74]};
    Full_Adder FA_7758(s7758, c7758, in7758_1, in7758_2, pp118[76]);
    wire[0:0] s7759, in7759_1, in7759_2;
    wire c7759;
    assign in7759_1 = {pp122[72]};
    assign in7759_2 = {pp123[71]};
    Full_Adder FA_7759(s7759, c7759, in7759_1, in7759_2, pp121[73]);
    wire[0:0] s7760, in7760_1, in7760_2;
    wire c7760;
    assign in7760_1 = {pp125[69]};
    assign in7760_2 = {pp126[68]};
    Full_Adder FA_7760(s7760, c7760, in7760_1, in7760_2, pp124[70]);
    wire[0:0] s7761, in7761_1, in7761_2;
    wire c7761;
    assign in7761_1 = {c4956};
    assign in7761_2 = {c4957};
    Full_Adder FA_7761(s7761, c7761, in7761_1, in7761_2, pp127[67]);
    wire[0:0] s7762, in7762_1, in7762_2;
    wire c7762;
    assign in7762_1 = {c4959};
    assign in7762_2 = {c4960};
    Full_Adder FA_7762(s7762, c7762, in7762_1, in7762_2, c4958);
    wire[0:0] s7763, in7763_1, in7763_2;
    wire c7763;
    assign in7763_1 = {s4962[0]};
    assign in7763_2 = {s4963[0]};
    Full_Adder FA_7763(s7763, c7763, in7763_1, in7763_2, s4961[0]);
    wire[0:0] s7764, in7764_1, in7764_2;
    wire c7764;
    assign in7764_1 = {pp78[117]};
    assign in7764_2 = {pp79[116]};
    Full_Adder FA_7764(s7764, c7764, in7764_1, in7764_2, pp77[118]);
    wire[0:0] s7765, in7765_1, in7765_2;
    wire c7765;
    assign in7765_1 = {pp81[114]};
    assign in7765_2 = {pp82[113]};
    Full_Adder FA_7765(s7765, c7765, in7765_1, in7765_2, pp80[115]);
    wire[0:0] s7766, in7766_1, in7766_2;
    wire c7766;
    assign in7766_1 = {pp84[111]};
    assign in7766_2 = {pp85[110]};
    Full_Adder FA_7766(s7766, c7766, in7766_1, in7766_2, pp83[112]);
    wire[0:0] s7767, in7767_1, in7767_2;
    wire c7767;
    assign in7767_1 = {pp87[108]};
    assign in7767_2 = {pp88[107]};
    Full_Adder FA_7767(s7767, c7767, in7767_1, in7767_2, pp86[109]);
    wire[0:0] s7768, in7768_1, in7768_2;
    wire c7768;
    assign in7768_1 = {pp90[105]};
    assign in7768_2 = {pp91[104]};
    Full_Adder FA_7768(s7768, c7768, in7768_1, in7768_2, pp89[106]);
    wire[0:0] s7769, in7769_1, in7769_2;
    wire c7769;
    assign in7769_1 = {pp93[102]};
    assign in7769_2 = {pp94[101]};
    Full_Adder FA_7769(s7769, c7769, in7769_1, in7769_2, pp92[103]);
    wire[0:0] s7770, in7770_1, in7770_2;
    wire c7770;
    assign in7770_1 = {pp96[99]};
    assign in7770_2 = {pp97[98]};
    Full_Adder FA_7770(s7770, c7770, in7770_1, in7770_2, pp95[100]);
    wire[0:0] s7771, in7771_1, in7771_2;
    wire c7771;
    assign in7771_1 = {pp99[96]};
    assign in7771_2 = {pp100[95]};
    Full_Adder FA_7771(s7771, c7771, in7771_1, in7771_2, pp98[97]);
    wire[0:0] s7772, in7772_1, in7772_2;
    wire c7772;
    assign in7772_1 = {pp102[93]};
    assign in7772_2 = {pp103[92]};
    Full_Adder FA_7772(s7772, c7772, in7772_1, in7772_2, pp101[94]);
    wire[0:0] s7773, in7773_1, in7773_2;
    wire c7773;
    assign in7773_1 = {pp105[90]};
    assign in7773_2 = {pp106[89]};
    Full_Adder FA_7773(s7773, c7773, in7773_1, in7773_2, pp104[91]);
    wire[0:0] s7774, in7774_1, in7774_2;
    wire c7774;
    assign in7774_1 = {pp108[87]};
    assign in7774_2 = {pp109[86]};
    Full_Adder FA_7774(s7774, c7774, in7774_1, in7774_2, pp107[88]);
    wire[0:0] s7775, in7775_1, in7775_2;
    wire c7775;
    assign in7775_1 = {pp111[84]};
    assign in7775_2 = {pp112[83]};
    Full_Adder FA_7775(s7775, c7775, in7775_1, in7775_2, pp110[85]);
    wire[0:0] s7776, in7776_1, in7776_2;
    wire c7776;
    assign in7776_1 = {pp114[81]};
    assign in7776_2 = {pp115[80]};
    Full_Adder FA_7776(s7776, c7776, in7776_1, in7776_2, pp113[82]);
    wire[0:0] s7777, in7777_1, in7777_2;
    wire c7777;
    assign in7777_1 = {pp117[78]};
    assign in7777_2 = {pp118[77]};
    Full_Adder FA_7777(s7777, c7777, in7777_1, in7777_2, pp116[79]);
    wire[0:0] s7778, in7778_1, in7778_2;
    wire c7778;
    assign in7778_1 = {pp120[75]};
    assign in7778_2 = {pp121[74]};
    Full_Adder FA_7778(s7778, c7778, in7778_1, in7778_2, pp119[76]);
    wire[0:0] s7779, in7779_1, in7779_2;
    wire c7779;
    assign in7779_1 = {pp123[72]};
    assign in7779_2 = {pp124[71]};
    Full_Adder FA_7779(s7779, c7779, in7779_1, in7779_2, pp122[73]);
    wire[0:0] s7780, in7780_1, in7780_2;
    wire c7780;
    assign in7780_1 = {pp126[69]};
    assign in7780_2 = {pp127[68]};
    Full_Adder FA_7780(s7780, c7780, in7780_1, in7780_2, pp125[70]);
    wire[0:0] s7781, in7781_1, in7781_2;
    wire c7781;
    assign in7781_1 = {c4962};
    assign in7781_2 = {c4963};
    Full_Adder FA_7781(s7781, c7781, in7781_1, in7781_2, c4961);
    wire[0:0] s7782, in7782_1, in7782_2;
    wire c7782;
    assign in7782_1 = {s4965[0]};
    assign in7782_2 = {s4966[0]};
    Full_Adder FA_7782(s7782, c7782, in7782_1, in7782_2, c4964);
    wire[0:0] s7783, in7783_1, in7783_2;
    wire c7783;
    assign in7783_1 = {pp76[120]};
    assign in7783_2 = {pp77[119]};
    Full_Adder FA_7783(s7783, c7783, in7783_1, in7783_2, pp75[121]);
    wire[0:0] s7784, in7784_1, in7784_2;
    wire c7784;
    assign in7784_1 = {pp79[117]};
    assign in7784_2 = {pp80[116]};
    Full_Adder FA_7784(s7784, c7784, in7784_1, in7784_2, pp78[118]);
    wire[0:0] s7785, in7785_1, in7785_2;
    wire c7785;
    assign in7785_1 = {pp82[114]};
    assign in7785_2 = {pp83[113]};
    Full_Adder FA_7785(s7785, c7785, in7785_1, in7785_2, pp81[115]);
    wire[0:0] s7786, in7786_1, in7786_2;
    wire c7786;
    assign in7786_1 = {pp85[111]};
    assign in7786_2 = {pp86[110]};
    Full_Adder FA_7786(s7786, c7786, in7786_1, in7786_2, pp84[112]);
    wire[0:0] s7787, in7787_1, in7787_2;
    wire c7787;
    assign in7787_1 = {pp88[108]};
    assign in7787_2 = {pp89[107]};
    Full_Adder FA_7787(s7787, c7787, in7787_1, in7787_2, pp87[109]);
    wire[0:0] s7788, in7788_1, in7788_2;
    wire c7788;
    assign in7788_1 = {pp91[105]};
    assign in7788_2 = {pp92[104]};
    Full_Adder FA_7788(s7788, c7788, in7788_1, in7788_2, pp90[106]);
    wire[0:0] s7789, in7789_1, in7789_2;
    wire c7789;
    assign in7789_1 = {pp94[102]};
    assign in7789_2 = {pp95[101]};
    Full_Adder FA_7789(s7789, c7789, in7789_1, in7789_2, pp93[103]);
    wire[0:0] s7790, in7790_1, in7790_2;
    wire c7790;
    assign in7790_1 = {pp97[99]};
    assign in7790_2 = {pp98[98]};
    Full_Adder FA_7790(s7790, c7790, in7790_1, in7790_2, pp96[100]);
    wire[0:0] s7791, in7791_1, in7791_2;
    wire c7791;
    assign in7791_1 = {pp100[96]};
    assign in7791_2 = {pp101[95]};
    Full_Adder FA_7791(s7791, c7791, in7791_1, in7791_2, pp99[97]);
    wire[0:0] s7792, in7792_1, in7792_2;
    wire c7792;
    assign in7792_1 = {pp103[93]};
    assign in7792_2 = {pp104[92]};
    Full_Adder FA_7792(s7792, c7792, in7792_1, in7792_2, pp102[94]);
    wire[0:0] s7793, in7793_1, in7793_2;
    wire c7793;
    assign in7793_1 = {pp106[90]};
    assign in7793_2 = {pp107[89]};
    Full_Adder FA_7793(s7793, c7793, in7793_1, in7793_2, pp105[91]);
    wire[0:0] s7794, in7794_1, in7794_2;
    wire c7794;
    assign in7794_1 = {pp109[87]};
    assign in7794_2 = {pp110[86]};
    Full_Adder FA_7794(s7794, c7794, in7794_1, in7794_2, pp108[88]);
    wire[0:0] s7795, in7795_1, in7795_2;
    wire c7795;
    assign in7795_1 = {pp112[84]};
    assign in7795_2 = {pp113[83]};
    Full_Adder FA_7795(s7795, c7795, in7795_1, in7795_2, pp111[85]);
    wire[0:0] s7796, in7796_1, in7796_2;
    wire c7796;
    assign in7796_1 = {pp115[81]};
    assign in7796_2 = {pp116[80]};
    Full_Adder FA_7796(s7796, c7796, in7796_1, in7796_2, pp114[82]);
    wire[0:0] s7797, in7797_1, in7797_2;
    wire c7797;
    assign in7797_1 = {pp118[78]};
    assign in7797_2 = {pp119[77]};
    Full_Adder FA_7797(s7797, c7797, in7797_1, in7797_2, pp117[79]);
    wire[0:0] s7798, in7798_1, in7798_2;
    wire c7798;
    assign in7798_1 = {pp121[75]};
    assign in7798_2 = {pp122[74]};
    Full_Adder FA_7798(s7798, c7798, in7798_1, in7798_2, pp120[76]);
    wire[0:0] s7799, in7799_1, in7799_2;
    wire c7799;
    assign in7799_1 = {pp124[72]};
    assign in7799_2 = {pp125[71]};
    Full_Adder FA_7799(s7799, c7799, in7799_1, in7799_2, pp123[73]);
    wire[0:0] s7800, in7800_1, in7800_2;
    wire c7800;
    assign in7800_1 = {pp127[69]};
    assign in7800_2 = {c4965};
    Full_Adder FA_7800(s7800, c7800, in7800_1, in7800_2, pp126[70]);
    wire[0:0] s7801, in7801_1, in7801_2;
    wire c7801;
    assign in7801_1 = {c4967};
    assign in7801_2 = {s4968[0]};
    Full_Adder FA_7801(s7801, c7801, in7801_1, in7801_2, c4966);
    wire[0:0] s7802, in7802_1, in7802_2;
    wire c7802;
    assign in7802_1 = {pp74[123]};
    assign in7802_2 = {pp75[122]};
    Full_Adder FA_7802(s7802, c7802, in7802_1, in7802_2, pp73[124]);
    wire[0:0] s7803, in7803_1, in7803_2;
    wire c7803;
    assign in7803_1 = {pp77[120]};
    assign in7803_2 = {pp78[119]};
    Full_Adder FA_7803(s7803, c7803, in7803_1, in7803_2, pp76[121]);
    wire[0:0] s7804, in7804_1, in7804_2;
    wire c7804;
    assign in7804_1 = {pp80[117]};
    assign in7804_2 = {pp81[116]};
    Full_Adder FA_7804(s7804, c7804, in7804_1, in7804_2, pp79[118]);
    wire[0:0] s7805, in7805_1, in7805_2;
    wire c7805;
    assign in7805_1 = {pp83[114]};
    assign in7805_2 = {pp84[113]};
    Full_Adder FA_7805(s7805, c7805, in7805_1, in7805_2, pp82[115]);
    wire[0:0] s7806, in7806_1, in7806_2;
    wire c7806;
    assign in7806_1 = {pp86[111]};
    assign in7806_2 = {pp87[110]};
    Full_Adder FA_7806(s7806, c7806, in7806_1, in7806_2, pp85[112]);
    wire[0:0] s7807, in7807_1, in7807_2;
    wire c7807;
    assign in7807_1 = {pp89[108]};
    assign in7807_2 = {pp90[107]};
    Full_Adder FA_7807(s7807, c7807, in7807_1, in7807_2, pp88[109]);
    wire[0:0] s7808, in7808_1, in7808_2;
    wire c7808;
    assign in7808_1 = {pp92[105]};
    assign in7808_2 = {pp93[104]};
    Full_Adder FA_7808(s7808, c7808, in7808_1, in7808_2, pp91[106]);
    wire[0:0] s7809, in7809_1, in7809_2;
    wire c7809;
    assign in7809_1 = {pp95[102]};
    assign in7809_2 = {pp96[101]};
    Full_Adder FA_7809(s7809, c7809, in7809_1, in7809_2, pp94[103]);
    wire[0:0] s7810, in7810_1, in7810_2;
    wire c7810;
    assign in7810_1 = {pp98[99]};
    assign in7810_2 = {pp99[98]};
    Full_Adder FA_7810(s7810, c7810, in7810_1, in7810_2, pp97[100]);
    wire[0:0] s7811, in7811_1, in7811_2;
    wire c7811;
    assign in7811_1 = {pp101[96]};
    assign in7811_2 = {pp102[95]};
    Full_Adder FA_7811(s7811, c7811, in7811_1, in7811_2, pp100[97]);
    wire[0:0] s7812, in7812_1, in7812_2;
    wire c7812;
    assign in7812_1 = {pp104[93]};
    assign in7812_2 = {pp105[92]};
    Full_Adder FA_7812(s7812, c7812, in7812_1, in7812_2, pp103[94]);
    wire[0:0] s7813, in7813_1, in7813_2;
    wire c7813;
    assign in7813_1 = {pp107[90]};
    assign in7813_2 = {pp108[89]};
    Full_Adder FA_7813(s7813, c7813, in7813_1, in7813_2, pp106[91]);
    wire[0:0] s7814, in7814_1, in7814_2;
    wire c7814;
    assign in7814_1 = {pp110[87]};
    assign in7814_2 = {pp111[86]};
    Full_Adder FA_7814(s7814, c7814, in7814_1, in7814_2, pp109[88]);
    wire[0:0] s7815, in7815_1, in7815_2;
    wire c7815;
    assign in7815_1 = {pp113[84]};
    assign in7815_2 = {pp114[83]};
    Full_Adder FA_7815(s7815, c7815, in7815_1, in7815_2, pp112[85]);
    wire[0:0] s7816, in7816_1, in7816_2;
    wire c7816;
    assign in7816_1 = {pp116[81]};
    assign in7816_2 = {pp117[80]};
    Full_Adder FA_7816(s7816, c7816, in7816_1, in7816_2, pp115[82]);
    wire[0:0] s7817, in7817_1, in7817_2;
    wire c7817;
    assign in7817_1 = {pp119[78]};
    assign in7817_2 = {pp120[77]};
    Full_Adder FA_7817(s7817, c7817, in7817_1, in7817_2, pp118[79]);
    wire[0:0] s7818, in7818_1, in7818_2;
    wire c7818;
    assign in7818_1 = {pp122[75]};
    assign in7818_2 = {pp123[74]};
    Full_Adder FA_7818(s7818, c7818, in7818_1, in7818_2, pp121[76]);
    wire[0:0] s7819, in7819_1, in7819_2;
    wire c7819;
    assign in7819_1 = {pp125[72]};
    assign in7819_2 = {pp126[71]};
    Full_Adder FA_7819(s7819, c7819, in7819_1, in7819_2, pp124[73]);
    wire[0:0] s7820, in7820_1, in7820_2;
    wire c7820;
    assign in7820_1 = {c4968};
    assign in7820_2 = {c4969};
    Full_Adder FA_7820(s7820, c7820, in7820_1, in7820_2, pp127[70]);
    wire[0:0] s7821, in7821_1, in7821_2;
    wire c7821;
    assign in7821_1 = {pp72[126]};
    assign in7821_2 = {pp73[125]};
    Full_Adder FA_7821(s7821, c7821, in7821_1, in7821_2, pp71[127]);
    wire[0:0] s7822, in7822_1, in7822_2;
    wire c7822;
    assign in7822_1 = {pp75[123]};
    assign in7822_2 = {pp76[122]};
    Full_Adder FA_7822(s7822, c7822, in7822_1, in7822_2, pp74[124]);
    wire[0:0] s7823, in7823_1, in7823_2;
    wire c7823;
    assign in7823_1 = {pp78[120]};
    assign in7823_2 = {pp79[119]};
    Full_Adder FA_7823(s7823, c7823, in7823_1, in7823_2, pp77[121]);
    wire[0:0] s7824, in7824_1, in7824_2;
    wire c7824;
    assign in7824_1 = {pp81[117]};
    assign in7824_2 = {pp82[116]};
    Full_Adder FA_7824(s7824, c7824, in7824_1, in7824_2, pp80[118]);
    wire[0:0] s7825, in7825_1, in7825_2;
    wire c7825;
    assign in7825_1 = {pp84[114]};
    assign in7825_2 = {pp85[113]};
    Full_Adder FA_7825(s7825, c7825, in7825_1, in7825_2, pp83[115]);
    wire[0:0] s7826, in7826_1, in7826_2;
    wire c7826;
    assign in7826_1 = {pp87[111]};
    assign in7826_2 = {pp88[110]};
    Full_Adder FA_7826(s7826, c7826, in7826_1, in7826_2, pp86[112]);
    wire[0:0] s7827, in7827_1, in7827_2;
    wire c7827;
    assign in7827_1 = {pp90[108]};
    assign in7827_2 = {pp91[107]};
    Full_Adder FA_7827(s7827, c7827, in7827_1, in7827_2, pp89[109]);
    wire[0:0] s7828, in7828_1, in7828_2;
    wire c7828;
    assign in7828_1 = {pp93[105]};
    assign in7828_2 = {pp94[104]};
    Full_Adder FA_7828(s7828, c7828, in7828_1, in7828_2, pp92[106]);
    wire[0:0] s7829, in7829_1, in7829_2;
    wire c7829;
    assign in7829_1 = {pp96[102]};
    assign in7829_2 = {pp97[101]};
    Full_Adder FA_7829(s7829, c7829, in7829_1, in7829_2, pp95[103]);
    wire[0:0] s7830, in7830_1, in7830_2;
    wire c7830;
    assign in7830_1 = {pp99[99]};
    assign in7830_2 = {pp100[98]};
    Full_Adder FA_7830(s7830, c7830, in7830_1, in7830_2, pp98[100]);
    wire[0:0] s7831, in7831_1, in7831_2;
    wire c7831;
    assign in7831_1 = {pp102[96]};
    assign in7831_2 = {pp103[95]};
    Full_Adder FA_7831(s7831, c7831, in7831_1, in7831_2, pp101[97]);
    wire[0:0] s7832, in7832_1, in7832_2;
    wire c7832;
    assign in7832_1 = {pp105[93]};
    assign in7832_2 = {pp106[92]};
    Full_Adder FA_7832(s7832, c7832, in7832_1, in7832_2, pp104[94]);
    wire[0:0] s7833, in7833_1, in7833_2;
    wire c7833;
    assign in7833_1 = {pp108[90]};
    assign in7833_2 = {pp109[89]};
    Full_Adder FA_7833(s7833, c7833, in7833_1, in7833_2, pp107[91]);
    wire[0:0] s7834, in7834_1, in7834_2;
    wire c7834;
    assign in7834_1 = {pp111[87]};
    assign in7834_2 = {pp112[86]};
    Full_Adder FA_7834(s7834, c7834, in7834_1, in7834_2, pp110[88]);
    wire[0:0] s7835, in7835_1, in7835_2;
    wire c7835;
    assign in7835_1 = {pp114[84]};
    assign in7835_2 = {pp115[83]};
    Full_Adder FA_7835(s7835, c7835, in7835_1, in7835_2, pp113[85]);
    wire[0:0] s7836, in7836_1, in7836_2;
    wire c7836;
    assign in7836_1 = {pp117[81]};
    assign in7836_2 = {pp118[80]};
    Full_Adder FA_7836(s7836, c7836, in7836_1, in7836_2, pp116[82]);
    wire[0:0] s7837, in7837_1, in7837_2;
    wire c7837;
    assign in7837_1 = {pp120[78]};
    assign in7837_2 = {pp121[77]};
    Full_Adder FA_7837(s7837, c7837, in7837_1, in7837_2, pp119[79]);
    wire[0:0] s7838, in7838_1, in7838_2;
    wire c7838;
    assign in7838_1 = {pp123[75]};
    assign in7838_2 = {pp124[74]};
    Full_Adder FA_7838(s7838, c7838, in7838_1, in7838_2, pp122[76]);
    wire[0:0] s7839, in7839_1, in7839_2;
    wire c7839;
    assign in7839_1 = {pp126[72]};
    assign in7839_2 = {pp127[71]};
    Full_Adder FA_7839(s7839, c7839, in7839_1, in7839_2, pp125[73]);
    wire[0:0] s7840, in7840_1, in7840_2;
    wire c7840;
    assign in7840_1 = {pp73[126]};
    assign in7840_2 = {pp74[125]};
    Full_Adder FA_7840(s7840, c7840, in7840_1, in7840_2, pp72[127]);
    wire[0:0] s7841, in7841_1, in7841_2;
    wire c7841;
    assign in7841_1 = {pp76[123]};
    assign in7841_2 = {pp77[122]};
    Full_Adder FA_7841(s7841, c7841, in7841_1, in7841_2, pp75[124]);
    wire[0:0] s7842, in7842_1, in7842_2;
    wire c7842;
    assign in7842_1 = {pp79[120]};
    assign in7842_2 = {pp80[119]};
    Full_Adder FA_7842(s7842, c7842, in7842_1, in7842_2, pp78[121]);
    wire[0:0] s7843, in7843_1, in7843_2;
    wire c7843;
    assign in7843_1 = {pp82[117]};
    assign in7843_2 = {pp83[116]};
    Full_Adder FA_7843(s7843, c7843, in7843_1, in7843_2, pp81[118]);
    wire[0:0] s7844, in7844_1, in7844_2;
    wire c7844;
    assign in7844_1 = {pp85[114]};
    assign in7844_2 = {pp86[113]};
    Full_Adder FA_7844(s7844, c7844, in7844_1, in7844_2, pp84[115]);
    wire[0:0] s7845, in7845_1, in7845_2;
    wire c7845;
    assign in7845_1 = {pp88[111]};
    assign in7845_2 = {pp89[110]};
    Full_Adder FA_7845(s7845, c7845, in7845_1, in7845_2, pp87[112]);
    wire[0:0] s7846, in7846_1, in7846_2;
    wire c7846;
    assign in7846_1 = {pp91[108]};
    assign in7846_2 = {pp92[107]};
    Full_Adder FA_7846(s7846, c7846, in7846_1, in7846_2, pp90[109]);
    wire[0:0] s7847, in7847_1, in7847_2;
    wire c7847;
    assign in7847_1 = {pp94[105]};
    assign in7847_2 = {pp95[104]};
    Full_Adder FA_7847(s7847, c7847, in7847_1, in7847_2, pp93[106]);
    wire[0:0] s7848, in7848_1, in7848_2;
    wire c7848;
    assign in7848_1 = {pp97[102]};
    assign in7848_2 = {pp98[101]};
    Full_Adder FA_7848(s7848, c7848, in7848_1, in7848_2, pp96[103]);
    wire[0:0] s7849, in7849_1, in7849_2;
    wire c7849;
    assign in7849_1 = {pp100[99]};
    assign in7849_2 = {pp101[98]};
    Full_Adder FA_7849(s7849, c7849, in7849_1, in7849_2, pp99[100]);
    wire[0:0] s7850, in7850_1, in7850_2;
    wire c7850;
    assign in7850_1 = {pp103[96]};
    assign in7850_2 = {pp104[95]};
    Full_Adder FA_7850(s7850, c7850, in7850_1, in7850_2, pp102[97]);
    wire[0:0] s7851, in7851_1, in7851_2;
    wire c7851;
    assign in7851_1 = {pp106[93]};
    assign in7851_2 = {pp107[92]};
    Full_Adder FA_7851(s7851, c7851, in7851_1, in7851_2, pp105[94]);
    wire[0:0] s7852, in7852_1, in7852_2;
    wire c7852;
    assign in7852_1 = {pp109[90]};
    assign in7852_2 = {pp110[89]};
    Full_Adder FA_7852(s7852, c7852, in7852_1, in7852_2, pp108[91]);
    wire[0:0] s7853, in7853_1, in7853_2;
    wire c7853;
    assign in7853_1 = {pp112[87]};
    assign in7853_2 = {pp113[86]};
    Full_Adder FA_7853(s7853, c7853, in7853_1, in7853_2, pp111[88]);
    wire[0:0] s7854, in7854_1, in7854_2;
    wire c7854;
    assign in7854_1 = {pp115[84]};
    assign in7854_2 = {pp116[83]};
    Full_Adder FA_7854(s7854, c7854, in7854_1, in7854_2, pp114[85]);
    wire[0:0] s7855, in7855_1, in7855_2;
    wire c7855;
    assign in7855_1 = {pp118[81]};
    assign in7855_2 = {pp119[80]};
    Full_Adder FA_7855(s7855, c7855, in7855_1, in7855_2, pp117[82]);
    wire[0:0] s7856, in7856_1, in7856_2;
    wire c7856;
    assign in7856_1 = {pp121[78]};
    assign in7856_2 = {pp122[77]};
    Full_Adder FA_7856(s7856, c7856, in7856_1, in7856_2, pp120[79]);
    wire[0:0] s7857, in7857_1, in7857_2;
    wire c7857;
    assign in7857_1 = {pp124[75]};
    assign in7857_2 = {pp125[74]};
    Full_Adder FA_7857(s7857, c7857, in7857_1, in7857_2, pp123[76]);
    wire[0:0] s7858, in7858_1, in7858_2;
    wire c7858;
    assign in7858_1 = {pp74[126]};
    assign in7858_2 = {pp75[125]};
    Full_Adder FA_7858(s7858, c7858, in7858_1, in7858_2, pp73[127]);
    wire[0:0] s7859, in7859_1, in7859_2;
    wire c7859;
    assign in7859_1 = {pp77[123]};
    assign in7859_2 = {pp78[122]};
    Full_Adder FA_7859(s7859, c7859, in7859_1, in7859_2, pp76[124]);
    wire[0:0] s7860, in7860_1, in7860_2;
    wire c7860;
    assign in7860_1 = {pp80[120]};
    assign in7860_2 = {pp81[119]};
    Full_Adder FA_7860(s7860, c7860, in7860_1, in7860_2, pp79[121]);
    wire[0:0] s7861, in7861_1, in7861_2;
    wire c7861;
    assign in7861_1 = {pp83[117]};
    assign in7861_2 = {pp84[116]};
    Full_Adder FA_7861(s7861, c7861, in7861_1, in7861_2, pp82[118]);
    wire[0:0] s7862, in7862_1, in7862_2;
    wire c7862;
    assign in7862_1 = {pp86[114]};
    assign in7862_2 = {pp87[113]};
    Full_Adder FA_7862(s7862, c7862, in7862_1, in7862_2, pp85[115]);
    wire[0:0] s7863, in7863_1, in7863_2;
    wire c7863;
    assign in7863_1 = {pp89[111]};
    assign in7863_2 = {pp90[110]};
    Full_Adder FA_7863(s7863, c7863, in7863_1, in7863_2, pp88[112]);
    wire[0:0] s7864, in7864_1, in7864_2;
    wire c7864;
    assign in7864_1 = {pp92[108]};
    assign in7864_2 = {pp93[107]};
    Full_Adder FA_7864(s7864, c7864, in7864_1, in7864_2, pp91[109]);
    wire[0:0] s7865, in7865_1, in7865_2;
    wire c7865;
    assign in7865_1 = {pp95[105]};
    assign in7865_2 = {pp96[104]};
    Full_Adder FA_7865(s7865, c7865, in7865_1, in7865_2, pp94[106]);
    wire[0:0] s7866, in7866_1, in7866_2;
    wire c7866;
    assign in7866_1 = {pp98[102]};
    assign in7866_2 = {pp99[101]};
    Full_Adder FA_7866(s7866, c7866, in7866_1, in7866_2, pp97[103]);
    wire[0:0] s7867, in7867_1, in7867_2;
    wire c7867;
    assign in7867_1 = {pp101[99]};
    assign in7867_2 = {pp102[98]};
    Full_Adder FA_7867(s7867, c7867, in7867_1, in7867_2, pp100[100]);
    wire[0:0] s7868, in7868_1, in7868_2;
    wire c7868;
    assign in7868_1 = {pp104[96]};
    assign in7868_2 = {pp105[95]};
    Full_Adder FA_7868(s7868, c7868, in7868_1, in7868_2, pp103[97]);
    wire[0:0] s7869, in7869_1, in7869_2;
    wire c7869;
    assign in7869_1 = {pp107[93]};
    assign in7869_2 = {pp108[92]};
    Full_Adder FA_7869(s7869, c7869, in7869_1, in7869_2, pp106[94]);
    wire[0:0] s7870, in7870_1, in7870_2;
    wire c7870;
    assign in7870_1 = {pp110[90]};
    assign in7870_2 = {pp111[89]};
    Full_Adder FA_7870(s7870, c7870, in7870_1, in7870_2, pp109[91]);
    wire[0:0] s7871, in7871_1, in7871_2;
    wire c7871;
    assign in7871_1 = {pp113[87]};
    assign in7871_2 = {pp114[86]};
    Full_Adder FA_7871(s7871, c7871, in7871_1, in7871_2, pp112[88]);
    wire[0:0] s7872, in7872_1, in7872_2;
    wire c7872;
    assign in7872_1 = {pp116[84]};
    assign in7872_2 = {pp117[83]};
    Full_Adder FA_7872(s7872, c7872, in7872_1, in7872_2, pp115[85]);
    wire[0:0] s7873, in7873_1, in7873_2;
    wire c7873;
    assign in7873_1 = {pp119[81]};
    assign in7873_2 = {pp120[80]};
    Full_Adder FA_7873(s7873, c7873, in7873_1, in7873_2, pp118[82]);
    wire[0:0] s7874, in7874_1, in7874_2;
    wire c7874;
    assign in7874_1 = {pp122[78]};
    assign in7874_2 = {pp123[77]};
    Full_Adder FA_7874(s7874, c7874, in7874_1, in7874_2, pp121[79]);
    wire[0:0] s7875, in7875_1, in7875_2;
    wire c7875;
    assign in7875_1 = {pp75[126]};
    assign in7875_2 = {pp76[125]};
    Full_Adder FA_7875(s7875, c7875, in7875_1, in7875_2, pp74[127]);
    wire[0:0] s7876, in7876_1, in7876_2;
    wire c7876;
    assign in7876_1 = {pp78[123]};
    assign in7876_2 = {pp79[122]};
    Full_Adder FA_7876(s7876, c7876, in7876_1, in7876_2, pp77[124]);
    wire[0:0] s7877, in7877_1, in7877_2;
    wire c7877;
    assign in7877_1 = {pp81[120]};
    assign in7877_2 = {pp82[119]};
    Full_Adder FA_7877(s7877, c7877, in7877_1, in7877_2, pp80[121]);
    wire[0:0] s7878, in7878_1, in7878_2;
    wire c7878;
    assign in7878_1 = {pp84[117]};
    assign in7878_2 = {pp85[116]};
    Full_Adder FA_7878(s7878, c7878, in7878_1, in7878_2, pp83[118]);
    wire[0:0] s7879, in7879_1, in7879_2;
    wire c7879;
    assign in7879_1 = {pp87[114]};
    assign in7879_2 = {pp88[113]};
    Full_Adder FA_7879(s7879, c7879, in7879_1, in7879_2, pp86[115]);
    wire[0:0] s7880, in7880_1, in7880_2;
    wire c7880;
    assign in7880_1 = {pp90[111]};
    assign in7880_2 = {pp91[110]};
    Full_Adder FA_7880(s7880, c7880, in7880_1, in7880_2, pp89[112]);
    wire[0:0] s7881, in7881_1, in7881_2;
    wire c7881;
    assign in7881_1 = {pp93[108]};
    assign in7881_2 = {pp94[107]};
    Full_Adder FA_7881(s7881, c7881, in7881_1, in7881_2, pp92[109]);
    wire[0:0] s7882, in7882_1, in7882_2;
    wire c7882;
    assign in7882_1 = {pp96[105]};
    assign in7882_2 = {pp97[104]};
    Full_Adder FA_7882(s7882, c7882, in7882_1, in7882_2, pp95[106]);
    wire[0:0] s7883, in7883_1, in7883_2;
    wire c7883;
    assign in7883_1 = {pp99[102]};
    assign in7883_2 = {pp100[101]};
    Full_Adder FA_7883(s7883, c7883, in7883_1, in7883_2, pp98[103]);
    wire[0:0] s7884, in7884_1, in7884_2;
    wire c7884;
    assign in7884_1 = {pp102[99]};
    assign in7884_2 = {pp103[98]};
    Full_Adder FA_7884(s7884, c7884, in7884_1, in7884_2, pp101[100]);
    wire[0:0] s7885, in7885_1, in7885_2;
    wire c7885;
    assign in7885_1 = {pp105[96]};
    assign in7885_2 = {pp106[95]};
    Full_Adder FA_7885(s7885, c7885, in7885_1, in7885_2, pp104[97]);
    wire[0:0] s7886, in7886_1, in7886_2;
    wire c7886;
    assign in7886_1 = {pp108[93]};
    assign in7886_2 = {pp109[92]};
    Full_Adder FA_7886(s7886, c7886, in7886_1, in7886_2, pp107[94]);
    wire[0:0] s7887, in7887_1, in7887_2;
    wire c7887;
    assign in7887_1 = {pp111[90]};
    assign in7887_2 = {pp112[89]};
    Full_Adder FA_7887(s7887, c7887, in7887_1, in7887_2, pp110[91]);
    wire[0:0] s7888, in7888_1, in7888_2;
    wire c7888;
    assign in7888_1 = {pp114[87]};
    assign in7888_2 = {pp115[86]};
    Full_Adder FA_7888(s7888, c7888, in7888_1, in7888_2, pp113[88]);
    wire[0:0] s7889, in7889_1, in7889_2;
    wire c7889;
    assign in7889_1 = {pp117[84]};
    assign in7889_2 = {pp118[83]};
    Full_Adder FA_7889(s7889, c7889, in7889_1, in7889_2, pp116[85]);
    wire[0:0] s7890, in7890_1, in7890_2;
    wire c7890;
    assign in7890_1 = {pp120[81]};
    assign in7890_2 = {pp121[80]};
    Full_Adder FA_7890(s7890, c7890, in7890_1, in7890_2, pp119[82]);
    wire[0:0] s7891, in7891_1, in7891_2;
    wire c7891;
    assign in7891_1 = {pp76[126]};
    assign in7891_2 = {pp77[125]};
    Full_Adder FA_7891(s7891, c7891, in7891_1, in7891_2, pp75[127]);
    wire[0:0] s7892, in7892_1, in7892_2;
    wire c7892;
    assign in7892_1 = {pp79[123]};
    assign in7892_2 = {pp80[122]};
    Full_Adder FA_7892(s7892, c7892, in7892_1, in7892_2, pp78[124]);
    wire[0:0] s7893, in7893_1, in7893_2;
    wire c7893;
    assign in7893_1 = {pp82[120]};
    assign in7893_2 = {pp83[119]};
    Full_Adder FA_7893(s7893, c7893, in7893_1, in7893_2, pp81[121]);
    wire[0:0] s7894, in7894_1, in7894_2;
    wire c7894;
    assign in7894_1 = {pp85[117]};
    assign in7894_2 = {pp86[116]};
    Full_Adder FA_7894(s7894, c7894, in7894_1, in7894_2, pp84[118]);
    wire[0:0] s7895, in7895_1, in7895_2;
    wire c7895;
    assign in7895_1 = {pp88[114]};
    assign in7895_2 = {pp89[113]};
    Full_Adder FA_7895(s7895, c7895, in7895_1, in7895_2, pp87[115]);
    wire[0:0] s7896, in7896_1, in7896_2;
    wire c7896;
    assign in7896_1 = {pp91[111]};
    assign in7896_2 = {pp92[110]};
    Full_Adder FA_7896(s7896, c7896, in7896_1, in7896_2, pp90[112]);
    wire[0:0] s7897, in7897_1, in7897_2;
    wire c7897;
    assign in7897_1 = {pp94[108]};
    assign in7897_2 = {pp95[107]};
    Full_Adder FA_7897(s7897, c7897, in7897_1, in7897_2, pp93[109]);
    wire[0:0] s7898, in7898_1, in7898_2;
    wire c7898;
    assign in7898_1 = {pp97[105]};
    assign in7898_2 = {pp98[104]};
    Full_Adder FA_7898(s7898, c7898, in7898_1, in7898_2, pp96[106]);
    wire[0:0] s7899, in7899_1, in7899_2;
    wire c7899;
    assign in7899_1 = {pp100[102]};
    assign in7899_2 = {pp101[101]};
    Full_Adder FA_7899(s7899, c7899, in7899_1, in7899_2, pp99[103]);
    wire[0:0] s7900, in7900_1, in7900_2;
    wire c7900;
    assign in7900_1 = {pp103[99]};
    assign in7900_2 = {pp104[98]};
    Full_Adder FA_7900(s7900, c7900, in7900_1, in7900_2, pp102[100]);
    wire[0:0] s7901, in7901_1, in7901_2;
    wire c7901;
    assign in7901_1 = {pp106[96]};
    assign in7901_2 = {pp107[95]};
    Full_Adder FA_7901(s7901, c7901, in7901_1, in7901_2, pp105[97]);
    wire[0:0] s7902, in7902_1, in7902_2;
    wire c7902;
    assign in7902_1 = {pp109[93]};
    assign in7902_2 = {pp110[92]};
    Full_Adder FA_7902(s7902, c7902, in7902_1, in7902_2, pp108[94]);
    wire[0:0] s7903, in7903_1, in7903_2;
    wire c7903;
    assign in7903_1 = {pp112[90]};
    assign in7903_2 = {pp113[89]};
    Full_Adder FA_7903(s7903, c7903, in7903_1, in7903_2, pp111[91]);
    wire[0:0] s7904, in7904_1, in7904_2;
    wire c7904;
    assign in7904_1 = {pp115[87]};
    assign in7904_2 = {pp116[86]};
    Full_Adder FA_7904(s7904, c7904, in7904_1, in7904_2, pp114[88]);
    wire[0:0] s7905, in7905_1, in7905_2;
    wire c7905;
    assign in7905_1 = {pp118[84]};
    assign in7905_2 = {pp119[83]};
    Full_Adder FA_7905(s7905, c7905, in7905_1, in7905_2, pp117[85]);
    wire[0:0] s7906, in7906_1, in7906_2;
    wire c7906;
    assign in7906_1 = {pp77[126]};
    assign in7906_2 = {pp78[125]};
    Full_Adder FA_7906(s7906, c7906, in7906_1, in7906_2, pp76[127]);
    wire[0:0] s7907, in7907_1, in7907_2;
    wire c7907;
    assign in7907_1 = {pp80[123]};
    assign in7907_2 = {pp81[122]};
    Full_Adder FA_7907(s7907, c7907, in7907_1, in7907_2, pp79[124]);
    wire[0:0] s7908, in7908_1, in7908_2;
    wire c7908;
    assign in7908_1 = {pp83[120]};
    assign in7908_2 = {pp84[119]};
    Full_Adder FA_7908(s7908, c7908, in7908_1, in7908_2, pp82[121]);
    wire[0:0] s7909, in7909_1, in7909_2;
    wire c7909;
    assign in7909_1 = {pp86[117]};
    assign in7909_2 = {pp87[116]};
    Full_Adder FA_7909(s7909, c7909, in7909_1, in7909_2, pp85[118]);
    wire[0:0] s7910, in7910_1, in7910_2;
    wire c7910;
    assign in7910_1 = {pp89[114]};
    assign in7910_2 = {pp90[113]};
    Full_Adder FA_7910(s7910, c7910, in7910_1, in7910_2, pp88[115]);
    wire[0:0] s7911, in7911_1, in7911_2;
    wire c7911;
    assign in7911_1 = {pp92[111]};
    assign in7911_2 = {pp93[110]};
    Full_Adder FA_7911(s7911, c7911, in7911_1, in7911_2, pp91[112]);
    wire[0:0] s7912, in7912_1, in7912_2;
    wire c7912;
    assign in7912_1 = {pp95[108]};
    assign in7912_2 = {pp96[107]};
    Full_Adder FA_7912(s7912, c7912, in7912_1, in7912_2, pp94[109]);
    wire[0:0] s7913, in7913_1, in7913_2;
    wire c7913;
    assign in7913_1 = {pp98[105]};
    assign in7913_2 = {pp99[104]};
    Full_Adder FA_7913(s7913, c7913, in7913_1, in7913_2, pp97[106]);
    wire[0:0] s7914, in7914_1, in7914_2;
    wire c7914;
    assign in7914_1 = {pp101[102]};
    assign in7914_2 = {pp102[101]};
    Full_Adder FA_7914(s7914, c7914, in7914_1, in7914_2, pp100[103]);
    wire[0:0] s7915, in7915_1, in7915_2;
    wire c7915;
    assign in7915_1 = {pp104[99]};
    assign in7915_2 = {pp105[98]};
    Full_Adder FA_7915(s7915, c7915, in7915_1, in7915_2, pp103[100]);
    wire[0:0] s7916, in7916_1, in7916_2;
    wire c7916;
    assign in7916_1 = {pp107[96]};
    assign in7916_2 = {pp108[95]};
    Full_Adder FA_7916(s7916, c7916, in7916_1, in7916_2, pp106[97]);
    wire[0:0] s7917, in7917_1, in7917_2;
    wire c7917;
    assign in7917_1 = {pp110[93]};
    assign in7917_2 = {pp111[92]};
    Full_Adder FA_7917(s7917, c7917, in7917_1, in7917_2, pp109[94]);
    wire[0:0] s7918, in7918_1, in7918_2;
    wire c7918;
    assign in7918_1 = {pp113[90]};
    assign in7918_2 = {pp114[89]};
    Full_Adder FA_7918(s7918, c7918, in7918_1, in7918_2, pp112[91]);
    wire[0:0] s7919, in7919_1, in7919_2;
    wire c7919;
    assign in7919_1 = {pp116[87]};
    assign in7919_2 = {pp117[86]};
    Full_Adder FA_7919(s7919, c7919, in7919_1, in7919_2, pp115[88]);
    wire[0:0] s7920, in7920_1, in7920_2;
    wire c7920;
    assign in7920_1 = {pp78[126]};
    assign in7920_2 = {pp79[125]};
    Full_Adder FA_7920(s7920, c7920, in7920_1, in7920_2, pp77[127]);
    wire[0:0] s7921, in7921_1, in7921_2;
    wire c7921;
    assign in7921_1 = {pp81[123]};
    assign in7921_2 = {pp82[122]};
    Full_Adder FA_7921(s7921, c7921, in7921_1, in7921_2, pp80[124]);
    wire[0:0] s7922, in7922_1, in7922_2;
    wire c7922;
    assign in7922_1 = {pp84[120]};
    assign in7922_2 = {pp85[119]};
    Full_Adder FA_7922(s7922, c7922, in7922_1, in7922_2, pp83[121]);
    wire[0:0] s7923, in7923_1, in7923_2;
    wire c7923;
    assign in7923_1 = {pp87[117]};
    assign in7923_2 = {pp88[116]};
    Full_Adder FA_7923(s7923, c7923, in7923_1, in7923_2, pp86[118]);
    wire[0:0] s7924, in7924_1, in7924_2;
    wire c7924;
    assign in7924_1 = {pp90[114]};
    assign in7924_2 = {pp91[113]};
    Full_Adder FA_7924(s7924, c7924, in7924_1, in7924_2, pp89[115]);
    wire[0:0] s7925, in7925_1, in7925_2;
    wire c7925;
    assign in7925_1 = {pp93[111]};
    assign in7925_2 = {pp94[110]};
    Full_Adder FA_7925(s7925, c7925, in7925_1, in7925_2, pp92[112]);
    wire[0:0] s7926, in7926_1, in7926_2;
    wire c7926;
    assign in7926_1 = {pp96[108]};
    assign in7926_2 = {pp97[107]};
    Full_Adder FA_7926(s7926, c7926, in7926_1, in7926_2, pp95[109]);
    wire[0:0] s7927, in7927_1, in7927_2;
    wire c7927;
    assign in7927_1 = {pp99[105]};
    assign in7927_2 = {pp100[104]};
    Full_Adder FA_7927(s7927, c7927, in7927_1, in7927_2, pp98[106]);
    wire[0:0] s7928, in7928_1, in7928_2;
    wire c7928;
    assign in7928_1 = {pp102[102]};
    assign in7928_2 = {pp103[101]};
    Full_Adder FA_7928(s7928, c7928, in7928_1, in7928_2, pp101[103]);
    wire[0:0] s7929, in7929_1, in7929_2;
    wire c7929;
    assign in7929_1 = {pp105[99]};
    assign in7929_2 = {pp106[98]};
    Full_Adder FA_7929(s7929, c7929, in7929_1, in7929_2, pp104[100]);
    wire[0:0] s7930, in7930_1, in7930_2;
    wire c7930;
    assign in7930_1 = {pp108[96]};
    assign in7930_2 = {pp109[95]};
    Full_Adder FA_7930(s7930, c7930, in7930_1, in7930_2, pp107[97]);
    wire[0:0] s7931, in7931_1, in7931_2;
    wire c7931;
    assign in7931_1 = {pp111[93]};
    assign in7931_2 = {pp112[92]};
    Full_Adder FA_7931(s7931, c7931, in7931_1, in7931_2, pp110[94]);
    wire[0:0] s7932, in7932_1, in7932_2;
    wire c7932;
    assign in7932_1 = {pp114[90]};
    assign in7932_2 = {pp115[89]};
    Full_Adder FA_7932(s7932, c7932, in7932_1, in7932_2, pp113[91]);
    wire[0:0] s7933, in7933_1, in7933_2;
    wire c7933;
    assign in7933_1 = {pp79[126]};
    assign in7933_2 = {pp80[125]};
    Full_Adder FA_7933(s7933, c7933, in7933_1, in7933_2, pp78[127]);
    wire[0:0] s7934, in7934_1, in7934_2;
    wire c7934;
    assign in7934_1 = {pp82[123]};
    assign in7934_2 = {pp83[122]};
    Full_Adder FA_7934(s7934, c7934, in7934_1, in7934_2, pp81[124]);
    wire[0:0] s7935, in7935_1, in7935_2;
    wire c7935;
    assign in7935_1 = {pp85[120]};
    assign in7935_2 = {pp86[119]};
    Full_Adder FA_7935(s7935, c7935, in7935_1, in7935_2, pp84[121]);
    wire[0:0] s7936, in7936_1, in7936_2;
    wire c7936;
    assign in7936_1 = {pp88[117]};
    assign in7936_2 = {pp89[116]};
    Full_Adder FA_7936(s7936, c7936, in7936_1, in7936_2, pp87[118]);
    wire[0:0] s7937, in7937_1, in7937_2;
    wire c7937;
    assign in7937_1 = {pp91[114]};
    assign in7937_2 = {pp92[113]};
    Full_Adder FA_7937(s7937, c7937, in7937_1, in7937_2, pp90[115]);
    wire[0:0] s7938, in7938_1, in7938_2;
    wire c7938;
    assign in7938_1 = {pp94[111]};
    assign in7938_2 = {pp95[110]};
    Full_Adder FA_7938(s7938, c7938, in7938_1, in7938_2, pp93[112]);
    wire[0:0] s7939, in7939_1, in7939_2;
    wire c7939;
    assign in7939_1 = {pp97[108]};
    assign in7939_2 = {pp98[107]};
    Full_Adder FA_7939(s7939, c7939, in7939_1, in7939_2, pp96[109]);
    wire[0:0] s7940, in7940_1, in7940_2;
    wire c7940;
    assign in7940_1 = {pp100[105]};
    assign in7940_2 = {pp101[104]};
    Full_Adder FA_7940(s7940, c7940, in7940_1, in7940_2, pp99[106]);
    wire[0:0] s7941, in7941_1, in7941_2;
    wire c7941;
    assign in7941_1 = {pp103[102]};
    assign in7941_2 = {pp104[101]};
    Full_Adder FA_7941(s7941, c7941, in7941_1, in7941_2, pp102[103]);
    wire[0:0] s7942, in7942_1, in7942_2;
    wire c7942;
    assign in7942_1 = {pp106[99]};
    assign in7942_2 = {pp107[98]};
    Full_Adder FA_7942(s7942, c7942, in7942_1, in7942_2, pp105[100]);
    wire[0:0] s7943, in7943_1, in7943_2;
    wire c7943;
    assign in7943_1 = {pp109[96]};
    assign in7943_2 = {pp110[95]};
    Full_Adder FA_7943(s7943, c7943, in7943_1, in7943_2, pp108[97]);
    wire[0:0] s7944, in7944_1, in7944_2;
    wire c7944;
    assign in7944_1 = {pp112[93]};
    assign in7944_2 = {pp113[92]};
    Full_Adder FA_7944(s7944, c7944, in7944_1, in7944_2, pp111[94]);
    wire[0:0] s7945, in7945_1, in7945_2;
    wire c7945;
    assign in7945_1 = {pp80[126]};
    assign in7945_2 = {pp81[125]};
    Full_Adder FA_7945(s7945, c7945, in7945_1, in7945_2, pp79[127]);
    wire[0:0] s7946, in7946_1, in7946_2;
    wire c7946;
    assign in7946_1 = {pp83[123]};
    assign in7946_2 = {pp84[122]};
    Full_Adder FA_7946(s7946, c7946, in7946_1, in7946_2, pp82[124]);
    wire[0:0] s7947, in7947_1, in7947_2;
    wire c7947;
    assign in7947_1 = {pp86[120]};
    assign in7947_2 = {pp87[119]};
    Full_Adder FA_7947(s7947, c7947, in7947_1, in7947_2, pp85[121]);
    wire[0:0] s7948, in7948_1, in7948_2;
    wire c7948;
    assign in7948_1 = {pp89[117]};
    assign in7948_2 = {pp90[116]};
    Full_Adder FA_7948(s7948, c7948, in7948_1, in7948_2, pp88[118]);
    wire[0:0] s7949, in7949_1, in7949_2;
    wire c7949;
    assign in7949_1 = {pp92[114]};
    assign in7949_2 = {pp93[113]};
    Full_Adder FA_7949(s7949, c7949, in7949_1, in7949_2, pp91[115]);
    wire[0:0] s7950, in7950_1, in7950_2;
    wire c7950;
    assign in7950_1 = {pp95[111]};
    assign in7950_2 = {pp96[110]};
    Full_Adder FA_7950(s7950, c7950, in7950_1, in7950_2, pp94[112]);
    wire[0:0] s7951, in7951_1, in7951_2;
    wire c7951;
    assign in7951_1 = {pp98[108]};
    assign in7951_2 = {pp99[107]};
    Full_Adder FA_7951(s7951, c7951, in7951_1, in7951_2, pp97[109]);
    wire[0:0] s7952, in7952_1, in7952_2;
    wire c7952;
    assign in7952_1 = {pp101[105]};
    assign in7952_2 = {pp102[104]};
    Full_Adder FA_7952(s7952, c7952, in7952_1, in7952_2, pp100[106]);
    wire[0:0] s7953, in7953_1, in7953_2;
    wire c7953;
    assign in7953_1 = {pp104[102]};
    assign in7953_2 = {pp105[101]};
    Full_Adder FA_7953(s7953, c7953, in7953_1, in7953_2, pp103[103]);
    wire[0:0] s7954, in7954_1, in7954_2;
    wire c7954;
    assign in7954_1 = {pp107[99]};
    assign in7954_2 = {pp108[98]};
    Full_Adder FA_7954(s7954, c7954, in7954_1, in7954_2, pp106[100]);
    wire[0:0] s7955, in7955_1, in7955_2;
    wire c7955;
    assign in7955_1 = {pp110[96]};
    assign in7955_2 = {pp111[95]};
    Full_Adder FA_7955(s7955, c7955, in7955_1, in7955_2, pp109[97]);
    wire[0:0] s7956, in7956_1, in7956_2;
    wire c7956;
    assign in7956_1 = {pp81[126]};
    assign in7956_2 = {pp82[125]};
    Full_Adder FA_7956(s7956, c7956, in7956_1, in7956_2, pp80[127]);
    wire[0:0] s7957, in7957_1, in7957_2;
    wire c7957;
    assign in7957_1 = {pp84[123]};
    assign in7957_2 = {pp85[122]};
    Full_Adder FA_7957(s7957, c7957, in7957_1, in7957_2, pp83[124]);
    wire[0:0] s7958, in7958_1, in7958_2;
    wire c7958;
    assign in7958_1 = {pp87[120]};
    assign in7958_2 = {pp88[119]};
    Full_Adder FA_7958(s7958, c7958, in7958_1, in7958_2, pp86[121]);
    wire[0:0] s7959, in7959_1, in7959_2;
    wire c7959;
    assign in7959_1 = {pp90[117]};
    assign in7959_2 = {pp91[116]};
    Full_Adder FA_7959(s7959, c7959, in7959_1, in7959_2, pp89[118]);
    wire[0:0] s7960, in7960_1, in7960_2;
    wire c7960;
    assign in7960_1 = {pp93[114]};
    assign in7960_2 = {pp94[113]};
    Full_Adder FA_7960(s7960, c7960, in7960_1, in7960_2, pp92[115]);
    wire[0:0] s7961, in7961_1, in7961_2;
    wire c7961;
    assign in7961_1 = {pp96[111]};
    assign in7961_2 = {pp97[110]};
    Full_Adder FA_7961(s7961, c7961, in7961_1, in7961_2, pp95[112]);
    wire[0:0] s7962, in7962_1, in7962_2;
    wire c7962;
    assign in7962_1 = {pp99[108]};
    assign in7962_2 = {pp100[107]};
    Full_Adder FA_7962(s7962, c7962, in7962_1, in7962_2, pp98[109]);
    wire[0:0] s7963, in7963_1, in7963_2;
    wire c7963;
    assign in7963_1 = {pp102[105]};
    assign in7963_2 = {pp103[104]};
    Full_Adder FA_7963(s7963, c7963, in7963_1, in7963_2, pp101[106]);
    wire[0:0] s7964, in7964_1, in7964_2;
    wire c7964;
    assign in7964_1 = {pp105[102]};
    assign in7964_2 = {pp106[101]};
    Full_Adder FA_7964(s7964, c7964, in7964_1, in7964_2, pp104[103]);
    wire[0:0] s7965, in7965_1, in7965_2;
    wire c7965;
    assign in7965_1 = {pp108[99]};
    assign in7965_2 = {pp109[98]};
    Full_Adder FA_7965(s7965, c7965, in7965_1, in7965_2, pp107[100]);
    wire[0:0] s7966, in7966_1, in7966_2;
    wire c7966;
    assign in7966_1 = {pp82[126]};
    assign in7966_2 = {pp83[125]};
    Full_Adder FA_7966(s7966, c7966, in7966_1, in7966_2, pp81[127]);
    wire[0:0] s7967, in7967_1, in7967_2;
    wire c7967;
    assign in7967_1 = {pp85[123]};
    assign in7967_2 = {pp86[122]};
    Full_Adder FA_7967(s7967, c7967, in7967_1, in7967_2, pp84[124]);
    wire[0:0] s7968, in7968_1, in7968_2;
    wire c7968;
    assign in7968_1 = {pp88[120]};
    assign in7968_2 = {pp89[119]};
    Full_Adder FA_7968(s7968, c7968, in7968_1, in7968_2, pp87[121]);
    wire[0:0] s7969, in7969_1, in7969_2;
    wire c7969;
    assign in7969_1 = {pp91[117]};
    assign in7969_2 = {pp92[116]};
    Full_Adder FA_7969(s7969, c7969, in7969_1, in7969_2, pp90[118]);
    wire[0:0] s7970, in7970_1, in7970_2;
    wire c7970;
    assign in7970_1 = {pp94[114]};
    assign in7970_2 = {pp95[113]};
    Full_Adder FA_7970(s7970, c7970, in7970_1, in7970_2, pp93[115]);
    wire[0:0] s7971, in7971_1, in7971_2;
    wire c7971;
    assign in7971_1 = {pp97[111]};
    assign in7971_2 = {pp98[110]};
    Full_Adder FA_7971(s7971, c7971, in7971_1, in7971_2, pp96[112]);
    wire[0:0] s7972, in7972_1, in7972_2;
    wire c7972;
    assign in7972_1 = {pp100[108]};
    assign in7972_2 = {pp101[107]};
    Full_Adder FA_7972(s7972, c7972, in7972_1, in7972_2, pp99[109]);
    wire[0:0] s7973, in7973_1, in7973_2;
    wire c7973;
    assign in7973_1 = {pp103[105]};
    assign in7973_2 = {pp104[104]};
    Full_Adder FA_7973(s7973, c7973, in7973_1, in7973_2, pp102[106]);
    wire[0:0] s7974, in7974_1, in7974_2;
    wire c7974;
    assign in7974_1 = {pp106[102]};
    assign in7974_2 = {pp107[101]};
    Full_Adder FA_7974(s7974, c7974, in7974_1, in7974_2, pp105[103]);
    wire[0:0] s7975, in7975_1, in7975_2;
    wire c7975;
    assign in7975_1 = {pp83[126]};
    assign in7975_2 = {pp84[125]};
    Full_Adder FA_7975(s7975, c7975, in7975_1, in7975_2, pp82[127]);
    wire[0:0] s7976, in7976_1, in7976_2;
    wire c7976;
    assign in7976_1 = {pp86[123]};
    assign in7976_2 = {pp87[122]};
    Full_Adder FA_7976(s7976, c7976, in7976_1, in7976_2, pp85[124]);
    wire[0:0] s7977, in7977_1, in7977_2;
    wire c7977;
    assign in7977_1 = {pp89[120]};
    assign in7977_2 = {pp90[119]};
    Full_Adder FA_7977(s7977, c7977, in7977_1, in7977_2, pp88[121]);
    wire[0:0] s7978, in7978_1, in7978_2;
    wire c7978;
    assign in7978_1 = {pp92[117]};
    assign in7978_2 = {pp93[116]};
    Full_Adder FA_7978(s7978, c7978, in7978_1, in7978_2, pp91[118]);
    wire[0:0] s7979, in7979_1, in7979_2;
    wire c7979;
    assign in7979_1 = {pp95[114]};
    assign in7979_2 = {pp96[113]};
    Full_Adder FA_7979(s7979, c7979, in7979_1, in7979_2, pp94[115]);
    wire[0:0] s7980, in7980_1, in7980_2;
    wire c7980;
    assign in7980_1 = {pp98[111]};
    assign in7980_2 = {pp99[110]};
    Full_Adder FA_7980(s7980, c7980, in7980_1, in7980_2, pp97[112]);
    wire[0:0] s7981, in7981_1, in7981_2;
    wire c7981;
    assign in7981_1 = {pp101[108]};
    assign in7981_2 = {pp102[107]};
    Full_Adder FA_7981(s7981, c7981, in7981_1, in7981_2, pp100[109]);
    wire[0:0] s7982, in7982_1, in7982_2;
    wire c7982;
    assign in7982_1 = {pp104[105]};
    assign in7982_2 = {pp105[104]};
    Full_Adder FA_7982(s7982, c7982, in7982_1, in7982_2, pp103[106]);
    wire[0:0] s7983, in7983_1, in7983_2;
    wire c7983;
    assign in7983_1 = {pp84[126]};
    assign in7983_2 = {pp85[125]};
    Full_Adder FA_7983(s7983, c7983, in7983_1, in7983_2, pp83[127]);
    wire[0:0] s7984, in7984_1, in7984_2;
    wire c7984;
    assign in7984_1 = {pp87[123]};
    assign in7984_2 = {pp88[122]};
    Full_Adder FA_7984(s7984, c7984, in7984_1, in7984_2, pp86[124]);
    wire[0:0] s7985, in7985_1, in7985_2;
    wire c7985;
    assign in7985_1 = {pp90[120]};
    assign in7985_2 = {pp91[119]};
    Full_Adder FA_7985(s7985, c7985, in7985_1, in7985_2, pp89[121]);
    wire[0:0] s7986, in7986_1, in7986_2;
    wire c7986;
    assign in7986_1 = {pp93[117]};
    assign in7986_2 = {pp94[116]};
    Full_Adder FA_7986(s7986, c7986, in7986_1, in7986_2, pp92[118]);
    wire[0:0] s7987, in7987_1, in7987_2;
    wire c7987;
    assign in7987_1 = {pp96[114]};
    assign in7987_2 = {pp97[113]};
    Full_Adder FA_7987(s7987, c7987, in7987_1, in7987_2, pp95[115]);
    wire[0:0] s7988, in7988_1, in7988_2;
    wire c7988;
    assign in7988_1 = {pp99[111]};
    assign in7988_2 = {pp100[110]};
    Full_Adder FA_7988(s7988, c7988, in7988_1, in7988_2, pp98[112]);
    wire[0:0] s7989, in7989_1, in7989_2;
    wire c7989;
    assign in7989_1 = {pp102[108]};
    assign in7989_2 = {pp103[107]};
    Full_Adder FA_7989(s7989, c7989, in7989_1, in7989_2, pp101[109]);
    wire[0:0] s7990, in7990_1, in7990_2;
    wire c7990;
    assign in7990_1 = {pp85[126]};
    assign in7990_2 = {pp86[125]};
    Full_Adder FA_7990(s7990, c7990, in7990_1, in7990_2, pp84[127]);
    wire[0:0] s7991, in7991_1, in7991_2;
    wire c7991;
    assign in7991_1 = {pp88[123]};
    assign in7991_2 = {pp89[122]};
    Full_Adder FA_7991(s7991, c7991, in7991_1, in7991_2, pp87[124]);
    wire[0:0] s7992, in7992_1, in7992_2;
    wire c7992;
    assign in7992_1 = {pp91[120]};
    assign in7992_2 = {pp92[119]};
    Full_Adder FA_7992(s7992, c7992, in7992_1, in7992_2, pp90[121]);
    wire[0:0] s7993, in7993_1, in7993_2;
    wire c7993;
    assign in7993_1 = {pp94[117]};
    assign in7993_2 = {pp95[116]};
    Full_Adder FA_7993(s7993, c7993, in7993_1, in7993_2, pp93[118]);
    wire[0:0] s7994, in7994_1, in7994_2;
    wire c7994;
    assign in7994_1 = {pp97[114]};
    assign in7994_2 = {pp98[113]};
    Full_Adder FA_7994(s7994, c7994, in7994_1, in7994_2, pp96[115]);
    wire[0:0] s7995, in7995_1, in7995_2;
    wire c7995;
    assign in7995_1 = {pp100[111]};
    assign in7995_2 = {pp101[110]};
    Full_Adder FA_7995(s7995, c7995, in7995_1, in7995_2, pp99[112]);
    wire[0:0] s7996, in7996_1, in7996_2;
    wire c7996;
    assign in7996_1 = {pp86[126]};
    assign in7996_2 = {pp87[125]};
    Full_Adder FA_7996(s7996, c7996, in7996_1, in7996_2, pp85[127]);
    wire[0:0] s7997, in7997_1, in7997_2;
    wire c7997;
    assign in7997_1 = {pp89[123]};
    assign in7997_2 = {pp90[122]};
    Full_Adder FA_7997(s7997, c7997, in7997_1, in7997_2, pp88[124]);
    wire[0:0] s7998, in7998_1, in7998_2;
    wire c7998;
    assign in7998_1 = {pp92[120]};
    assign in7998_2 = {pp93[119]};
    Full_Adder FA_7998(s7998, c7998, in7998_1, in7998_2, pp91[121]);
    wire[0:0] s7999, in7999_1, in7999_2;
    wire c7999;
    assign in7999_1 = {pp95[117]};
    assign in7999_2 = {pp96[116]};
    Full_Adder FA_7999(s7999, c7999, in7999_1, in7999_2, pp94[118]);
    wire[0:0] s8000, in8000_1, in8000_2;
    wire c8000;
    assign in8000_1 = {pp98[114]};
    assign in8000_2 = {pp99[113]};
    Full_Adder FA_8000(s8000, c8000, in8000_1, in8000_2, pp97[115]);
    wire[0:0] s8001, in8001_1, in8001_2;
    wire c8001;
    assign in8001_1 = {pp87[126]};
    assign in8001_2 = {pp88[125]};
    Full_Adder FA_8001(s8001, c8001, in8001_1, in8001_2, pp86[127]);
    wire[0:0] s8002, in8002_1, in8002_2;
    wire c8002;
    assign in8002_1 = {pp90[123]};
    assign in8002_2 = {pp91[122]};
    Full_Adder FA_8002(s8002, c8002, in8002_1, in8002_2, pp89[124]);
    wire[0:0] s8003, in8003_1, in8003_2;
    wire c8003;
    assign in8003_1 = {pp93[120]};
    assign in8003_2 = {pp94[119]};
    Full_Adder FA_8003(s8003, c8003, in8003_1, in8003_2, pp92[121]);
    wire[0:0] s8004, in8004_1, in8004_2;
    wire c8004;
    assign in8004_1 = {pp96[117]};
    assign in8004_2 = {pp97[116]};
    Full_Adder FA_8004(s8004, c8004, in8004_1, in8004_2, pp95[118]);
    wire[0:0] s8005, in8005_1, in8005_2;
    wire c8005;
    assign in8005_1 = {pp88[126]};
    assign in8005_2 = {pp89[125]};
    Full_Adder FA_8005(s8005, c8005, in8005_1, in8005_2, pp87[127]);
    wire[0:0] s8006, in8006_1, in8006_2;
    wire c8006;
    assign in8006_1 = {pp91[123]};
    assign in8006_2 = {pp92[122]};
    Full_Adder FA_8006(s8006, c8006, in8006_1, in8006_2, pp90[124]);
    wire[0:0] s8007, in8007_1, in8007_2;
    wire c8007;
    assign in8007_1 = {pp94[120]};
    assign in8007_2 = {pp95[119]};
    Full_Adder FA_8007(s8007, c8007, in8007_1, in8007_2, pp93[121]);
    wire[0:0] s8008, in8008_1, in8008_2;
    wire c8008;
    assign in8008_1 = {pp89[126]};
    assign in8008_2 = {pp90[125]};
    Full_Adder FA_8008(s8008, c8008, in8008_1, in8008_2, pp88[127]);
    wire[0:0] s8009, in8009_1, in8009_2;
    wire c8009;
    assign in8009_1 = {pp92[123]};
    assign in8009_2 = {pp93[122]};
    Full_Adder FA_8009(s8009, c8009, in8009_1, in8009_2, pp91[124]);
    wire[0:0] s8010, in8010_1, in8010_2;
    wire c8010;
    assign in8010_1 = {pp90[126]};
    assign in8010_2 = {pp91[125]};
    Full_Adder FA_8010(s8010, c8010, in8010_1, in8010_2, pp89[127]);

    /*Stage 4*/
    wire[0:0] s8011, in8011_1, in8011_2;
    wire c8011;
    assign in8011_1 = {pp0[26]};
    assign in8011_2 = {pp1[25]};
    Half_Adder HA_8011(s8011, c8011, in8011_1, in8011_2);
    wire[0:0] s8012, in8012_1, in8012_2;
    wire c8012;
    assign in8012_1 = {pp1[26]};
    assign in8012_2 = {pp2[25]};
    Full_Adder FA_8012(s8012, c8012, in8012_1, in8012_2, pp0[27]);
    wire[0:0] s8013, in8013_1, in8013_2;
    wire c8013;
    assign in8013_1 = {pp3[24]};
    assign in8013_2 = {pp4[23]};
    Half_Adder HA_8013(s8013, c8013, in8013_1, in8013_2);
    wire[0:0] s8014, in8014_1, in8014_2;
    wire c8014;
    assign in8014_1 = {pp1[27]};
    assign in8014_2 = {pp2[26]};
    Full_Adder FA_8014(s8014, c8014, in8014_1, in8014_2, pp0[28]);
    wire[0:0] s8015, in8015_1, in8015_2;
    wire c8015;
    assign in8015_1 = {pp4[24]};
    assign in8015_2 = {pp5[23]};
    Full_Adder FA_8015(s8015, c8015, in8015_1, in8015_2, pp3[25]);
    wire[0:0] s8016, in8016_1, in8016_2;
    wire c8016;
    assign in8016_1 = {pp6[22]};
    assign in8016_2 = {pp7[21]};
    Half_Adder HA_8016(s8016, c8016, in8016_1, in8016_2);
    wire[0:0] s8017, in8017_1, in8017_2;
    wire c8017;
    assign in8017_1 = {pp1[28]};
    assign in8017_2 = {pp2[27]};
    Full_Adder FA_8017(s8017, c8017, in8017_1, in8017_2, pp0[29]);
    wire[0:0] s8018, in8018_1, in8018_2;
    wire c8018;
    assign in8018_1 = {pp4[25]};
    assign in8018_2 = {pp5[24]};
    Full_Adder FA_8018(s8018, c8018, in8018_1, in8018_2, pp3[26]);
    wire[0:0] s8019, in8019_1, in8019_2;
    wire c8019;
    assign in8019_1 = {pp7[22]};
    assign in8019_2 = {pp8[21]};
    Full_Adder FA_8019(s8019, c8019, in8019_1, in8019_2, pp6[23]);
    wire[0:0] s8020, in8020_1, in8020_2;
    wire c8020;
    assign in8020_1 = {pp9[20]};
    assign in8020_2 = {pp10[19]};
    Half_Adder HA_8020(s8020, c8020, in8020_1, in8020_2);
    wire[0:0] s8021, in8021_1, in8021_2;
    wire c8021;
    assign in8021_1 = {pp1[29]};
    assign in8021_2 = {pp2[28]};
    Full_Adder FA_8021(s8021, c8021, in8021_1, in8021_2, pp0[30]);
    wire[0:0] s8022, in8022_1, in8022_2;
    wire c8022;
    assign in8022_1 = {pp4[26]};
    assign in8022_2 = {pp5[25]};
    Full_Adder FA_8022(s8022, c8022, in8022_1, in8022_2, pp3[27]);
    wire[0:0] s8023, in8023_1, in8023_2;
    wire c8023;
    assign in8023_1 = {pp7[23]};
    assign in8023_2 = {pp8[22]};
    Full_Adder FA_8023(s8023, c8023, in8023_1, in8023_2, pp6[24]);
    wire[0:0] s8024, in8024_1, in8024_2;
    wire c8024;
    assign in8024_1 = {pp10[20]};
    assign in8024_2 = {pp11[19]};
    Full_Adder FA_8024(s8024, c8024, in8024_1, in8024_2, pp9[21]);
    wire[0:0] s8025, in8025_1, in8025_2;
    wire c8025;
    assign in8025_1 = {pp12[18]};
    assign in8025_2 = {pp13[17]};
    Half_Adder HA_8025(s8025, c8025, in8025_1, in8025_2);
    wire[0:0] s8026, in8026_1, in8026_2;
    wire c8026;
    assign in8026_1 = {pp1[30]};
    assign in8026_2 = {pp2[29]};
    Full_Adder FA_8026(s8026, c8026, in8026_1, in8026_2, pp0[31]);
    wire[0:0] s8027, in8027_1, in8027_2;
    wire c8027;
    assign in8027_1 = {pp4[27]};
    assign in8027_2 = {pp5[26]};
    Full_Adder FA_8027(s8027, c8027, in8027_1, in8027_2, pp3[28]);
    wire[0:0] s8028, in8028_1, in8028_2;
    wire c8028;
    assign in8028_1 = {pp7[24]};
    assign in8028_2 = {pp8[23]};
    Full_Adder FA_8028(s8028, c8028, in8028_1, in8028_2, pp6[25]);
    wire[0:0] s8029, in8029_1, in8029_2;
    wire c8029;
    assign in8029_1 = {pp10[21]};
    assign in8029_2 = {pp11[20]};
    Full_Adder FA_8029(s8029, c8029, in8029_1, in8029_2, pp9[22]);
    wire[0:0] s8030, in8030_1, in8030_2;
    wire c8030;
    assign in8030_1 = {pp13[18]};
    assign in8030_2 = {pp14[17]};
    Full_Adder FA_8030(s8030, c8030, in8030_1, in8030_2, pp12[19]);
    wire[0:0] s8031, in8031_1, in8031_2;
    wire c8031;
    assign in8031_1 = {pp15[16]};
    assign in8031_2 = {pp16[15]};
    Half_Adder HA_8031(s8031, c8031, in8031_1, in8031_2);
    wire[0:0] s8032, in8032_1, in8032_2;
    wire c8032;
    assign in8032_1 = {pp1[31]};
    assign in8032_2 = {pp2[30]};
    Full_Adder FA_8032(s8032, c8032, in8032_1, in8032_2, pp0[32]);
    wire[0:0] s8033, in8033_1, in8033_2;
    wire c8033;
    assign in8033_1 = {pp4[28]};
    assign in8033_2 = {pp5[27]};
    Full_Adder FA_8033(s8033, c8033, in8033_1, in8033_2, pp3[29]);
    wire[0:0] s8034, in8034_1, in8034_2;
    wire c8034;
    assign in8034_1 = {pp7[25]};
    assign in8034_2 = {pp8[24]};
    Full_Adder FA_8034(s8034, c8034, in8034_1, in8034_2, pp6[26]);
    wire[0:0] s8035, in8035_1, in8035_2;
    wire c8035;
    assign in8035_1 = {pp10[22]};
    assign in8035_2 = {pp11[21]};
    Full_Adder FA_8035(s8035, c8035, in8035_1, in8035_2, pp9[23]);
    wire[0:0] s8036, in8036_1, in8036_2;
    wire c8036;
    assign in8036_1 = {pp13[19]};
    assign in8036_2 = {pp14[18]};
    Full_Adder FA_8036(s8036, c8036, in8036_1, in8036_2, pp12[20]);
    wire[0:0] s8037, in8037_1, in8037_2;
    wire c8037;
    assign in8037_1 = {pp16[16]};
    assign in8037_2 = {pp17[15]};
    Full_Adder FA_8037(s8037, c8037, in8037_1, in8037_2, pp15[17]);
    wire[0:0] s8038, in8038_1, in8038_2;
    wire c8038;
    assign in8038_1 = {pp18[14]};
    assign in8038_2 = {pp19[13]};
    Half_Adder HA_8038(s8038, c8038, in8038_1, in8038_2);
    wire[0:0] s8039, in8039_1, in8039_2;
    wire c8039;
    assign in8039_1 = {pp1[32]};
    assign in8039_2 = {pp2[31]};
    Full_Adder FA_8039(s8039, c8039, in8039_1, in8039_2, pp0[33]);
    wire[0:0] s8040, in8040_1, in8040_2;
    wire c8040;
    assign in8040_1 = {pp4[29]};
    assign in8040_2 = {pp5[28]};
    Full_Adder FA_8040(s8040, c8040, in8040_1, in8040_2, pp3[30]);
    wire[0:0] s8041, in8041_1, in8041_2;
    wire c8041;
    assign in8041_1 = {pp7[26]};
    assign in8041_2 = {pp8[25]};
    Full_Adder FA_8041(s8041, c8041, in8041_1, in8041_2, pp6[27]);
    wire[0:0] s8042, in8042_1, in8042_2;
    wire c8042;
    assign in8042_1 = {pp10[23]};
    assign in8042_2 = {pp11[22]};
    Full_Adder FA_8042(s8042, c8042, in8042_1, in8042_2, pp9[24]);
    wire[0:0] s8043, in8043_1, in8043_2;
    wire c8043;
    assign in8043_1 = {pp13[20]};
    assign in8043_2 = {pp14[19]};
    Full_Adder FA_8043(s8043, c8043, in8043_1, in8043_2, pp12[21]);
    wire[0:0] s8044, in8044_1, in8044_2;
    wire c8044;
    assign in8044_1 = {pp16[17]};
    assign in8044_2 = {pp17[16]};
    Full_Adder FA_8044(s8044, c8044, in8044_1, in8044_2, pp15[18]);
    wire[0:0] s8045, in8045_1, in8045_2;
    wire c8045;
    assign in8045_1 = {pp19[14]};
    assign in8045_2 = {pp20[13]};
    Full_Adder FA_8045(s8045, c8045, in8045_1, in8045_2, pp18[15]);
    wire[0:0] s8046, in8046_1, in8046_2;
    wire c8046;
    assign in8046_1 = {pp21[12]};
    assign in8046_2 = {pp22[11]};
    Half_Adder HA_8046(s8046, c8046, in8046_1, in8046_2);
    wire[0:0] s8047, in8047_1, in8047_2;
    wire c8047;
    assign in8047_1 = {pp1[33]};
    assign in8047_2 = {pp2[32]};
    Full_Adder FA_8047(s8047, c8047, in8047_1, in8047_2, pp0[34]);
    wire[0:0] s8048, in8048_1, in8048_2;
    wire c8048;
    assign in8048_1 = {pp4[30]};
    assign in8048_2 = {pp5[29]};
    Full_Adder FA_8048(s8048, c8048, in8048_1, in8048_2, pp3[31]);
    wire[0:0] s8049, in8049_1, in8049_2;
    wire c8049;
    assign in8049_1 = {pp7[27]};
    assign in8049_2 = {pp8[26]};
    Full_Adder FA_8049(s8049, c8049, in8049_1, in8049_2, pp6[28]);
    wire[0:0] s8050, in8050_1, in8050_2;
    wire c8050;
    assign in8050_1 = {pp10[24]};
    assign in8050_2 = {pp11[23]};
    Full_Adder FA_8050(s8050, c8050, in8050_1, in8050_2, pp9[25]);
    wire[0:0] s8051, in8051_1, in8051_2;
    wire c8051;
    assign in8051_1 = {pp13[21]};
    assign in8051_2 = {pp14[20]};
    Full_Adder FA_8051(s8051, c8051, in8051_1, in8051_2, pp12[22]);
    wire[0:0] s8052, in8052_1, in8052_2;
    wire c8052;
    assign in8052_1 = {pp16[18]};
    assign in8052_2 = {pp17[17]};
    Full_Adder FA_8052(s8052, c8052, in8052_1, in8052_2, pp15[19]);
    wire[0:0] s8053, in8053_1, in8053_2;
    wire c8053;
    assign in8053_1 = {pp19[15]};
    assign in8053_2 = {pp20[14]};
    Full_Adder FA_8053(s8053, c8053, in8053_1, in8053_2, pp18[16]);
    wire[0:0] s8054, in8054_1, in8054_2;
    wire c8054;
    assign in8054_1 = {pp22[12]};
    assign in8054_2 = {pp23[11]};
    Full_Adder FA_8054(s8054, c8054, in8054_1, in8054_2, pp21[13]);
    wire[0:0] s8055, in8055_1, in8055_2;
    wire c8055;
    assign in8055_1 = {pp24[10]};
    assign in8055_2 = {pp25[9]};
    Half_Adder HA_8055(s8055, c8055, in8055_1, in8055_2);
    wire[0:0] s8056, in8056_1, in8056_2;
    wire c8056;
    assign in8056_1 = {pp1[34]};
    assign in8056_2 = {pp2[33]};
    Full_Adder FA_8056(s8056, c8056, in8056_1, in8056_2, pp0[35]);
    wire[0:0] s8057, in8057_1, in8057_2;
    wire c8057;
    assign in8057_1 = {pp4[31]};
    assign in8057_2 = {pp5[30]};
    Full_Adder FA_8057(s8057, c8057, in8057_1, in8057_2, pp3[32]);
    wire[0:0] s8058, in8058_1, in8058_2;
    wire c8058;
    assign in8058_1 = {pp7[28]};
    assign in8058_2 = {pp8[27]};
    Full_Adder FA_8058(s8058, c8058, in8058_1, in8058_2, pp6[29]);
    wire[0:0] s8059, in8059_1, in8059_2;
    wire c8059;
    assign in8059_1 = {pp10[25]};
    assign in8059_2 = {pp11[24]};
    Full_Adder FA_8059(s8059, c8059, in8059_1, in8059_2, pp9[26]);
    wire[0:0] s8060, in8060_1, in8060_2;
    wire c8060;
    assign in8060_1 = {pp13[22]};
    assign in8060_2 = {pp14[21]};
    Full_Adder FA_8060(s8060, c8060, in8060_1, in8060_2, pp12[23]);
    wire[0:0] s8061, in8061_1, in8061_2;
    wire c8061;
    assign in8061_1 = {pp16[19]};
    assign in8061_2 = {pp17[18]};
    Full_Adder FA_8061(s8061, c8061, in8061_1, in8061_2, pp15[20]);
    wire[0:0] s8062, in8062_1, in8062_2;
    wire c8062;
    assign in8062_1 = {pp19[16]};
    assign in8062_2 = {pp20[15]};
    Full_Adder FA_8062(s8062, c8062, in8062_1, in8062_2, pp18[17]);
    wire[0:0] s8063, in8063_1, in8063_2;
    wire c8063;
    assign in8063_1 = {pp22[13]};
    assign in8063_2 = {pp23[12]};
    Full_Adder FA_8063(s8063, c8063, in8063_1, in8063_2, pp21[14]);
    wire[0:0] s8064, in8064_1, in8064_2;
    wire c8064;
    assign in8064_1 = {pp25[10]};
    assign in8064_2 = {pp26[9]};
    Full_Adder FA_8064(s8064, c8064, in8064_1, in8064_2, pp24[11]);
    wire[0:0] s8065, in8065_1, in8065_2;
    wire c8065;
    assign in8065_1 = {pp27[8]};
    assign in8065_2 = {pp28[7]};
    Half_Adder HA_8065(s8065, c8065, in8065_1, in8065_2);
    wire[0:0] s8066, in8066_1, in8066_2;
    wire c8066;
    assign in8066_1 = {pp1[35]};
    assign in8066_2 = {pp2[34]};
    Full_Adder FA_8066(s8066, c8066, in8066_1, in8066_2, pp0[36]);
    wire[0:0] s8067, in8067_1, in8067_2;
    wire c8067;
    assign in8067_1 = {pp4[32]};
    assign in8067_2 = {pp5[31]};
    Full_Adder FA_8067(s8067, c8067, in8067_1, in8067_2, pp3[33]);
    wire[0:0] s8068, in8068_1, in8068_2;
    wire c8068;
    assign in8068_1 = {pp7[29]};
    assign in8068_2 = {pp8[28]};
    Full_Adder FA_8068(s8068, c8068, in8068_1, in8068_2, pp6[30]);
    wire[0:0] s8069, in8069_1, in8069_2;
    wire c8069;
    assign in8069_1 = {pp10[26]};
    assign in8069_2 = {pp11[25]};
    Full_Adder FA_8069(s8069, c8069, in8069_1, in8069_2, pp9[27]);
    wire[0:0] s8070, in8070_1, in8070_2;
    wire c8070;
    assign in8070_1 = {pp13[23]};
    assign in8070_2 = {pp14[22]};
    Full_Adder FA_8070(s8070, c8070, in8070_1, in8070_2, pp12[24]);
    wire[0:0] s8071, in8071_1, in8071_2;
    wire c8071;
    assign in8071_1 = {pp16[20]};
    assign in8071_2 = {pp17[19]};
    Full_Adder FA_8071(s8071, c8071, in8071_1, in8071_2, pp15[21]);
    wire[0:0] s8072, in8072_1, in8072_2;
    wire c8072;
    assign in8072_1 = {pp19[17]};
    assign in8072_2 = {pp20[16]};
    Full_Adder FA_8072(s8072, c8072, in8072_1, in8072_2, pp18[18]);
    wire[0:0] s8073, in8073_1, in8073_2;
    wire c8073;
    assign in8073_1 = {pp22[14]};
    assign in8073_2 = {pp23[13]};
    Full_Adder FA_8073(s8073, c8073, in8073_1, in8073_2, pp21[15]);
    wire[0:0] s8074, in8074_1, in8074_2;
    wire c8074;
    assign in8074_1 = {pp25[11]};
    assign in8074_2 = {pp26[10]};
    Full_Adder FA_8074(s8074, c8074, in8074_1, in8074_2, pp24[12]);
    wire[0:0] s8075, in8075_1, in8075_2;
    wire c8075;
    assign in8075_1 = {pp28[8]};
    assign in8075_2 = {pp29[7]};
    Full_Adder FA_8075(s8075, c8075, in8075_1, in8075_2, pp27[9]);
    wire[0:0] s8076, in8076_1, in8076_2;
    wire c8076;
    assign in8076_1 = {pp30[6]};
    assign in8076_2 = {pp31[5]};
    Half_Adder HA_8076(s8076, c8076, in8076_1, in8076_2);
    wire[0:0] s8077, in8077_1, in8077_2;
    wire c8077;
    assign in8077_1 = {pp1[36]};
    assign in8077_2 = {pp2[35]};
    Full_Adder FA_8077(s8077, c8077, in8077_1, in8077_2, pp0[37]);
    wire[0:0] s8078, in8078_1, in8078_2;
    wire c8078;
    assign in8078_1 = {pp4[33]};
    assign in8078_2 = {pp5[32]};
    Full_Adder FA_8078(s8078, c8078, in8078_1, in8078_2, pp3[34]);
    wire[0:0] s8079, in8079_1, in8079_2;
    wire c8079;
    assign in8079_1 = {pp7[30]};
    assign in8079_2 = {pp8[29]};
    Full_Adder FA_8079(s8079, c8079, in8079_1, in8079_2, pp6[31]);
    wire[0:0] s8080, in8080_1, in8080_2;
    wire c8080;
    assign in8080_1 = {pp10[27]};
    assign in8080_2 = {pp11[26]};
    Full_Adder FA_8080(s8080, c8080, in8080_1, in8080_2, pp9[28]);
    wire[0:0] s8081, in8081_1, in8081_2;
    wire c8081;
    assign in8081_1 = {pp13[24]};
    assign in8081_2 = {pp14[23]};
    Full_Adder FA_8081(s8081, c8081, in8081_1, in8081_2, pp12[25]);
    wire[0:0] s8082, in8082_1, in8082_2;
    wire c8082;
    assign in8082_1 = {pp16[21]};
    assign in8082_2 = {pp17[20]};
    Full_Adder FA_8082(s8082, c8082, in8082_1, in8082_2, pp15[22]);
    wire[0:0] s8083, in8083_1, in8083_2;
    wire c8083;
    assign in8083_1 = {pp19[18]};
    assign in8083_2 = {pp20[17]};
    Full_Adder FA_8083(s8083, c8083, in8083_1, in8083_2, pp18[19]);
    wire[0:0] s8084, in8084_1, in8084_2;
    wire c8084;
    assign in8084_1 = {pp22[15]};
    assign in8084_2 = {pp23[14]};
    Full_Adder FA_8084(s8084, c8084, in8084_1, in8084_2, pp21[16]);
    wire[0:0] s8085, in8085_1, in8085_2;
    wire c8085;
    assign in8085_1 = {pp25[12]};
    assign in8085_2 = {pp26[11]};
    Full_Adder FA_8085(s8085, c8085, in8085_1, in8085_2, pp24[13]);
    wire[0:0] s8086, in8086_1, in8086_2;
    wire c8086;
    assign in8086_1 = {pp28[9]};
    assign in8086_2 = {pp29[8]};
    Full_Adder FA_8086(s8086, c8086, in8086_1, in8086_2, pp27[10]);
    wire[0:0] s8087, in8087_1, in8087_2;
    wire c8087;
    assign in8087_1 = {pp31[6]};
    assign in8087_2 = {pp32[5]};
    Full_Adder FA_8087(s8087, c8087, in8087_1, in8087_2, pp30[7]);
    wire[0:0] s8088, in8088_1, in8088_2;
    wire c8088;
    assign in8088_1 = {pp33[4]};
    assign in8088_2 = {pp34[3]};
    Half_Adder HA_8088(s8088, c8088, in8088_1, in8088_2);
    wire[0:0] s8089, in8089_1, in8089_2;
    wire c8089;
    assign in8089_1 = {pp1[37]};
    assign in8089_2 = {pp2[36]};
    Full_Adder FA_8089(s8089, c8089, in8089_1, in8089_2, pp0[38]);
    wire[0:0] s8090, in8090_1, in8090_2;
    wire c8090;
    assign in8090_1 = {pp4[34]};
    assign in8090_2 = {pp5[33]};
    Full_Adder FA_8090(s8090, c8090, in8090_1, in8090_2, pp3[35]);
    wire[0:0] s8091, in8091_1, in8091_2;
    wire c8091;
    assign in8091_1 = {pp7[31]};
    assign in8091_2 = {pp8[30]};
    Full_Adder FA_8091(s8091, c8091, in8091_1, in8091_2, pp6[32]);
    wire[0:0] s8092, in8092_1, in8092_2;
    wire c8092;
    assign in8092_1 = {pp10[28]};
    assign in8092_2 = {pp11[27]};
    Full_Adder FA_8092(s8092, c8092, in8092_1, in8092_2, pp9[29]);
    wire[0:0] s8093, in8093_1, in8093_2;
    wire c8093;
    assign in8093_1 = {pp13[25]};
    assign in8093_2 = {pp14[24]};
    Full_Adder FA_8093(s8093, c8093, in8093_1, in8093_2, pp12[26]);
    wire[0:0] s8094, in8094_1, in8094_2;
    wire c8094;
    assign in8094_1 = {pp16[22]};
    assign in8094_2 = {pp17[21]};
    Full_Adder FA_8094(s8094, c8094, in8094_1, in8094_2, pp15[23]);
    wire[0:0] s8095, in8095_1, in8095_2;
    wire c8095;
    assign in8095_1 = {pp19[19]};
    assign in8095_2 = {pp20[18]};
    Full_Adder FA_8095(s8095, c8095, in8095_1, in8095_2, pp18[20]);
    wire[0:0] s8096, in8096_1, in8096_2;
    wire c8096;
    assign in8096_1 = {pp22[16]};
    assign in8096_2 = {pp23[15]};
    Full_Adder FA_8096(s8096, c8096, in8096_1, in8096_2, pp21[17]);
    wire[0:0] s8097, in8097_1, in8097_2;
    wire c8097;
    assign in8097_1 = {pp25[13]};
    assign in8097_2 = {pp26[12]};
    Full_Adder FA_8097(s8097, c8097, in8097_1, in8097_2, pp24[14]);
    wire[0:0] s8098, in8098_1, in8098_2;
    wire c8098;
    assign in8098_1 = {pp28[10]};
    assign in8098_2 = {pp29[9]};
    Full_Adder FA_8098(s8098, c8098, in8098_1, in8098_2, pp27[11]);
    wire[0:0] s8099, in8099_1, in8099_2;
    wire c8099;
    assign in8099_1 = {pp31[7]};
    assign in8099_2 = {pp32[6]};
    Full_Adder FA_8099(s8099, c8099, in8099_1, in8099_2, pp30[8]);
    wire[0:0] s8100, in8100_1, in8100_2;
    wire c8100;
    assign in8100_1 = {pp34[4]};
    assign in8100_2 = {pp35[3]};
    Full_Adder FA_8100(s8100, c8100, in8100_1, in8100_2, pp33[5]);
    wire[0:0] s8101, in8101_1, in8101_2;
    wire c8101;
    assign in8101_1 = {pp36[2]};
    assign in8101_2 = {pp37[1]};
    Half_Adder HA_8101(s8101, c8101, in8101_1, in8101_2);
    wire[0:0] s8102, in8102_1, in8102_2;
    wire c8102;
    assign in8102_1 = {pp3[36]};
    assign in8102_2 = {pp4[35]};
    Full_Adder FA_8102(s8102, c8102, in8102_1, in8102_2, pp2[37]);
    wire[0:0] s8103, in8103_1, in8103_2;
    wire c8103;
    assign in8103_1 = {pp6[33]};
    assign in8103_2 = {pp7[32]};
    Full_Adder FA_8103(s8103, c8103, in8103_1, in8103_2, pp5[34]);
    wire[0:0] s8104, in8104_1, in8104_2;
    wire c8104;
    assign in8104_1 = {pp9[30]};
    assign in8104_2 = {pp10[29]};
    Full_Adder FA_8104(s8104, c8104, in8104_1, in8104_2, pp8[31]);
    wire[0:0] s8105, in8105_1, in8105_2;
    wire c8105;
    assign in8105_1 = {pp12[27]};
    assign in8105_2 = {pp13[26]};
    Full_Adder FA_8105(s8105, c8105, in8105_1, in8105_2, pp11[28]);
    wire[0:0] s8106, in8106_1, in8106_2;
    wire c8106;
    assign in8106_1 = {pp15[24]};
    assign in8106_2 = {pp16[23]};
    Full_Adder FA_8106(s8106, c8106, in8106_1, in8106_2, pp14[25]);
    wire[0:0] s8107, in8107_1, in8107_2;
    wire c8107;
    assign in8107_1 = {pp18[21]};
    assign in8107_2 = {pp19[20]};
    Full_Adder FA_8107(s8107, c8107, in8107_1, in8107_2, pp17[22]);
    wire[0:0] s8108, in8108_1, in8108_2;
    wire c8108;
    assign in8108_1 = {pp21[18]};
    assign in8108_2 = {pp22[17]};
    Full_Adder FA_8108(s8108, c8108, in8108_1, in8108_2, pp20[19]);
    wire[0:0] s8109, in8109_1, in8109_2;
    wire c8109;
    assign in8109_1 = {pp24[15]};
    assign in8109_2 = {pp25[14]};
    Full_Adder FA_8109(s8109, c8109, in8109_1, in8109_2, pp23[16]);
    wire[0:0] s8110, in8110_1, in8110_2;
    wire c8110;
    assign in8110_1 = {pp27[12]};
    assign in8110_2 = {pp28[11]};
    Full_Adder FA_8110(s8110, c8110, in8110_1, in8110_2, pp26[13]);
    wire[0:0] s8111, in8111_1, in8111_2;
    wire c8111;
    assign in8111_1 = {pp30[9]};
    assign in8111_2 = {pp31[8]};
    Full_Adder FA_8111(s8111, c8111, in8111_1, in8111_2, pp29[10]);
    wire[0:0] s8112, in8112_1, in8112_2;
    wire c8112;
    assign in8112_1 = {pp33[6]};
    assign in8112_2 = {pp34[5]};
    Full_Adder FA_8112(s8112, c8112, in8112_1, in8112_2, pp32[7]);
    wire[0:0] s8113, in8113_1, in8113_2;
    wire c8113;
    assign in8113_1 = {pp36[3]};
    assign in8113_2 = {pp37[2]};
    Full_Adder FA_8113(s8113, c8113, in8113_1, in8113_2, pp35[4]);
    wire[0:0] s8114, in8114_1, in8114_2;
    wire c8114;
    assign in8114_1 = {pp39[0]};
    assign in8114_2 = {s4971[0]};
    Full_Adder FA_8114(s8114, c8114, in8114_1, in8114_2, pp38[1]);
    wire[0:0] s8115, in8115_1, in8115_2;
    wire c8115;
    assign in8115_1 = {pp6[34]};
    assign in8115_2 = {pp7[33]};
    Full_Adder FA_8115(s8115, c8115, in8115_1, in8115_2, pp5[35]);
    wire[0:0] s8116, in8116_1, in8116_2;
    wire c8116;
    assign in8116_1 = {pp9[31]};
    assign in8116_2 = {pp10[30]};
    Full_Adder FA_8116(s8116, c8116, in8116_1, in8116_2, pp8[32]);
    wire[0:0] s8117, in8117_1, in8117_2;
    wire c8117;
    assign in8117_1 = {pp12[28]};
    assign in8117_2 = {pp13[27]};
    Full_Adder FA_8117(s8117, c8117, in8117_1, in8117_2, pp11[29]);
    wire[0:0] s8118, in8118_1, in8118_2;
    wire c8118;
    assign in8118_1 = {pp15[25]};
    assign in8118_2 = {pp16[24]};
    Full_Adder FA_8118(s8118, c8118, in8118_1, in8118_2, pp14[26]);
    wire[0:0] s8119, in8119_1, in8119_2;
    wire c8119;
    assign in8119_1 = {pp18[22]};
    assign in8119_2 = {pp19[21]};
    Full_Adder FA_8119(s8119, c8119, in8119_1, in8119_2, pp17[23]);
    wire[0:0] s8120, in8120_1, in8120_2;
    wire c8120;
    assign in8120_1 = {pp21[19]};
    assign in8120_2 = {pp22[18]};
    Full_Adder FA_8120(s8120, c8120, in8120_1, in8120_2, pp20[20]);
    wire[0:0] s8121, in8121_1, in8121_2;
    wire c8121;
    assign in8121_1 = {pp24[16]};
    assign in8121_2 = {pp25[15]};
    Full_Adder FA_8121(s8121, c8121, in8121_1, in8121_2, pp23[17]);
    wire[0:0] s8122, in8122_1, in8122_2;
    wire c8122;
    assign in8122_1 = {pp27[13]};
    assign in8122_2 = {pp28[12]};
    Full_Adder FA_8122(s8122, c8122, in8122_1, in8122_2, pp26[14]);
    wire[0:0] s8123, in8123_1, in8123_2;
    wire c8123;
    assign in8123_1 = {pp30[10]};
    assign in8123_2 = {pp31[9]};
    Full_Adder FA_8123(s8123, c8123, in8123_1, in8123_2, pp29[11]);
    wire[0:0] s8124, in8124_1, in8124_2;
    wire c8124;
    assign in8124_1 = {pp33[7]};
    assign in8124_2 = {pp34[6]};
    Full_Adder FA_8124(s8124, c8124, in8124_1, in8124_2, pp32[8]);
    wire[0:0] s8125, in8125_1, in8125_2;
    wire c8125;
    assign in8125_1 = {pp36[4]};
    assign in8125_2 = {pp37[3]};
    Full_Adder FA_8125(s8125, c8125, in8125_1, in8125_2, pp35[5]);
    wire[0:0] s8126, in8126_1, in8126_2;
    wire c8126;
    assign in8126_1 = {pp39[1]};
    assign in8126_2 = {pp40[0]};
    Full_Adder FA_8126(s8126, c8126, in8126_1, in8126_2, pp38[2]);
    wire[0:0] s8127, in8127_1, in8127_2;
    wire c8127;
    assign in8127_1 = {s4972[0]};
    assign in8127_2 = {s4973[0]};
    Full_Adder FA_8127(s8127, c8127, in8127_1, in8127_2, c4971);
    wire[0:0] s8128, in8128_1, in8128_2;
    wire c8128;
    assign in8128_1 = {pp9[32]};
    assign in8128_2 = {pp10[31]};
    Full_Adder FA_8128(s8128, c8128, in8128_1, in8128_2, pp8[33]);
    wire[0:0] s8129, in8129_1, in8129_2;
    wire c8129;
    assign in8129_1 = {pp12[29]};
    assign in8129_2 = {pp13[28]};
    Full_Adder FA_8129(s8129, c8129, in8129_1, in8129_2, pp11[30]);
    wire[0:0] s8130, in8130_1, in8130_2;
    wire c8130;
    assign in8130_1 = {pp15[26]};
    assign in8130_2 = {pp16[25]};
    Full_Adder FA_8130(s8130, c8130, in8130_1, in8130_2, pp14[27]);
    wire[0:0] s8131, in8131_1, in8131_2;
    wire c8131;
    assign in8131_1 = {pp18[23]};
    assign in8131_2 = {pp19[22]};
    Full_Adder FA_8131(s8131, c8131, in8131_1, in8131_2, pp17[24]);
    wire[0:0] s8132, in8132_1, in8132_2;
    wire c8132;
    assign in8132_1 = {pp21[20]};
    assign in8132_2 = {pp22[19]};
    Full_Adder FA_8132(s8132, c8132, in8132_1, in8132_2, pp20[21]);
    wire[0:0] s8133, in8133_1, in8133_2;
    wire c8133;
    assign in8133_1 = {pp24[17]};
    assign in8133_2 = {pp25[16]};
    Full_Adder FA_8133(s8133, c8133, in8133_1, in8133_2, pp23[18]);
    wire[0:0] s8134, in8134_1, in8134_2;
    wire c8134;
    assign in8134_1 = {pp27[14]};
    assign in8134_2 = {pp28[13]};
    Full_Adder FA_8134(s8134, c8134, in8134_1, in8134_2, pp26[15]);
    wire[0:0] s8135, in8135_1, in8135_2;
    wire c8135;
    assign in8135_1 = {pp30[11]};
    assign in8135_2 = {pp31[10]};
    Full_Adder FA_8135(s8135, c8135, in8135_1, in8135_2, pp29[12]);
    wire[0:0] s8136, in8136_1, in8136_2;
    wire c8136;
    assign in8136_1 = {pp33[8]};
    assign in8136_2 = {pp34[7]};
    Full_Adder FA_8136(s8136, c8136, in8136_1, in8136_2, pp32[9]);
    wire[0:0] s8137, in8137_1, in8137_2;
    wire c8137;
    assign in8137_1 = {pp36[5]};
    assign in8137_2 = {pp37[4]};
    Full_Adder FA_8137(s8137, c8137, in8137_1, in8137_2, pp35[6]);
    wire[0:0] s8138, in8138_1, in8138_2;
    wire c8138;
    assign in8138_1 = {pp39[2]};
    assign in8138_2 = {pp40[1]};
    Full_Adder FA_8138(s8138, c8138, in8138_1, in8138_2, pp38[3]);
    wire[0:0] s8139, in8139_1, in8139_2;
    wire c8139;
    assign in8139_1 = {c4972};
    assign in8139_2 = {c4973};
    Full_Adder FA_8139(s8139, c8139, in8139_1, in8139_2, pp41[0]);
    wire[0:0] s8140, in8140_1, in8140_2;
    wire c8140;
    assign in8140_1 = {s4975[0]};
    assign in8140_2 = {s4976[0]};
    Full_Adder FA_8140(s8140, c8140, in8140_1, in8140_2, s4974[0]);
    wire[0:0] s8141, in8141_1, in8141_2;
    wire c8141;
    assign in8141_1 = {pp12[30]};
    assign in8141_2 = {pp13[29]};
    Full_Adder FA_8141(s8141, c8141, in8141_1, in8141_2, pp11[31]);
    wire[0:0] s8142, in8142_1, in8142_2;
    wire c8142;
    assign in8142_1 = {pp15[27]};
    assign in8142_2 = {pp16[26]};
    Full_Adder FA_8142(s8142, c8142, in8142_1, in8142_2, pp14[28]);
    wire[0:0] s8143, in8143_1, in8143_2;
    wire c8143;
    assign in8143_1 = {pp18[24]};
    assign in8143_2 = {pp19[23]};
    Full_Adder FA_8143(s8143, c8143, in8143_1, in8143_2, pp17[25]);
    wire[0:0] s8144, in8144_1, in8144_2;
    wire c8144;
    assign in8144_1 = {pp21[21]};
    assign in8144_2 = {pp22[20]};
    Full_Adder FA_8144(s8144, c8144, in8144_1, in8144_2, pp20[22]);
    wire[0:0] s8145, in8145_1, in8145_2;
    wire c8145;
    assign in8145_1 = {pp24[18]};
    assign in8145_2 = {pp25[17]};
    Full_Adder FA_8145(s8145, c8145, in8145_1, in8145_2, pp23[19]);
    wire[0:0] s8146, in8146_1, in8146_2;
    wire c8146;
    assign in8146_1 = {pp27[15]};
    assign in8146_2 = {pp28[14]};
    Full_Adder FA_8146(s8146, c8146, in8146_1, in8146_2, pp26[16]);
    wire[0:0] s8147, in8147_1, in8147_2;
    wire c8147;
    assign in8147_1 = {pp30[12]};
    assign in8147_2 = {pp31[11]};
    Full_Adder FA_8147(s8147, c8147, in8147_1, in8147_2, pp29[13]);
    wire[0:0] s8148, in8148_1, in8148_2;
    wire c8148;
    assign in8148_1 = {pp33[9]};
    assign in8148_2 = {pp34[8]};
    Full_Adder FA_8148(s8148, c8148, in8148_1, in8148_2, pp32[10]);
    wire[0:0] s8149, in8149_1, in8149_2;
    wire c8149;
    assign in8149_1 = {pp36[6]};
    assign in8149_2 = {pp37[5]};
    Full_Adder FA_8149(s8149, c8149, in8149_1, in8149_2, pp35[7]);
    wire[0:0] s8150, in8150_1, in8150_2;
    wire c8150;
    assign in8150_1 = {pp39[3]};
    assign in8150_2 = {pp40[2]};
    Full_Adder FA_8150(s8150, c8150, in8150_1, in8150_2, pp38[4]);
    wire[0:0] s8151, in8151_1, in8151_2;
    wire c8151;
    assign in8151_1 = {pp42[0]};
    assign in8151_2 = {c4974};
    Full_Adder FA_8151(s8151, c8151, in8151_1, in8151_2, pp41[1]);
    wire[0:0] s8152, in8152_1, in8152_2;
    wire c8152;
    assign in8152_1 = {c4976};
    assign in8152_2 = {s4977[0]};
    Full_Adder FA_8152(s8152, c8152, in8152_1, in8152_2, c4975);
    wire[0:0] s8153, in8153_1, in8153_2;
    wire c8153;
    assign in8153_1 = {s4979[0]};
    assign in8153_2 = {s4980[0]};
    Full_Adder FA_8153(s8153, c8153, in8153_1, in8153_2, s4978[0]);
    wire[0:0] s8154, in8154_1, in8154_2;
    wire c8154;
    assign in8154_1 = {pp15[28]};
    assign in8154_2 = {pp16[27]};
    Full_Adder FA_8154(s8154, c8154, in8154_1, in8154_2, pp14[29]);
    wire[0:0] s8155, in8155_1, in8155_2;
    wire c8155;
    assign in8155_1 = {pp18[25]};
    assign in8155_2 = {pp19[24]};
    Full_Adder FA_8155(s8155, c8155, in8155_1, in8155_2, pp17[26]);
    wire[0:0] s8156, in8156_1, in8156_2;
    wire c8156;
    assign in8156_1 = {pp21[22]};
    assign in8156_2 = {pp22[21]};
    Full_Adder FA_8156(s8156, c8156, in8156_1, in8156_2, pp20[23]);
    wire[0:0] s8157, in8157_1, in8157_2;
    wire c8157;
    assign in8157_1 = {pp24[19]};
    assign in8157_2 = {pp25[18]};
    Full_Adder FA_8157(s8157, c8157, in8157_1, in8157_2, pp23[20]);
    wire[0:0] s8158, in8158_1, in8158_2;
    wire c8158;
    assign in8158_1 = {pp27[16]};
    assign in8158_2 = {pp28[15]};
    Full_Adder FA_8158(s8158, c8158, in8158_1, in8158_2, pp26[17]);
    wire[0:0] s8159, in8159_1, in8159_2;
    wire c8159;
    assign in8159_1 = {pp30[13]};
    assign in8159_2 = {pp31[12]};
    Full_Adder FA_8159(s8159, c8159, in8159_1, in8159_2, pp29[14]);
    wire[0:0] s8160, in8160_1, in8160_2;
    wire c8160;
    assign in8160_1 = {pp33[10]};
    assign in8160_2 = {pp34[9]};
    Full_Adder FA_8160(s8160, c8160, in8160_1, in8160_2, pp32[11]);
    wire[0:0] s8161, in8161_1, in8161_2;
    wire c8161;
    assign in8161_1 = {pp36[7]};
    assign in8161_2 = {pp37[6]};
    Full_Adder FA_8161(s8161, c8161, in8161_1, in8161_2, pp35[8]);
    wire[0:0] s8162, in8162_1, in8162_2;
    wire c8162;
    assign in8162_1 = {pp39[4]};
    assign in8162_2 = {pp40[3]};
    Full_Adder FA_8162(s8162, c8162, in8162_1, in8162_2, pp38[5]);
    wire[0:0] s8163, in8163_1, in8163_2;
    wire c8163;
    assign in8163_1 = {pp42[1]};
    assign in8163_2 = {pp43[0]};
    Full_Adder FA_8163(s8163, c8163, in8163_1, in8163_2, pp41[2]);
    wire[0:0] s8164, in8164_1, in8164_2;
    wire c8164;
    assign in8164_1 = {c4978};
    assign in8164_2 = {c4979};
    Full_Adder FA_8164(s8164, c8164, in8164_1, in8164_2, c4977);
    wire[0:0] s8165, in8165_1, in8165_2;
    wire c8165;
    assign in8165_1 = {s4981[0]};
    assign in8165_2 = {s4982[0]};
    Full_Adder FA_8165(s8165, c8165, in8165_1, in8165_2, c4980);
    wire[0:0] s8166, in8166_1, in8166_2;
    wire c8166;
    assign in8166_1 = {s4984[0]};
    assign in8166_2 = {s4985[0]};
    Full_Adder FA_8166(s8166, c8166, in8166_1, in8166_2, s4983[0]);
    wire[0:0] s8167, in8167_1, in8167_2;
    wire c8167;
    assign in8167_1 = {pp18[26]};
    assign in8167_2 = {pp19[25]};
    Full_Adder FA_8167(s8167, c8167, in8167_1, in8167_2, pp17[27]);
    wire[0:0] s8168, in8168_1, in8168_2;
    wire c8168;
    assign in8168_1 = {pp21[23]};
    assign in8168_2 = {pp22[22]};
    Full_Adder FA_8168(s8168, c8168, in8168_1, in8168_2, pp20[24]);
    wire[0:0] s8169, in8169_1, in8169_2;
    wire c8169;
    assign in8169_1 = {pp24[20]};
    assign in8169_2 = {pp25[19]};
    Full_Adder FA_8169(s8169, c8169, in8169_1, in8169_2, pp23[21]);
    wire[0:0] s8170, in8170_1, in8170_2;
    wire c8170;
    assign in8170_1 = {pp27[17]};
    assign in8170_2 = {pp28[16]};
    Full_Adder FA_8170(s8170, c8170, in8170_1, in8170_2, pp26[18]);
    wire[0:0] s8171, in8171_1, in8171_2;
    wire c8171;
    assign in8171_1 = {pp30[14]};
    assign in8171_2 = {pp31[13]};
    Full_Adder FA_8171(s8171, c8171, in8171_1, in8171_2, pp29[15]);
    wire[0:0] s8172, in8172_1, in8172_2;
    wire c8172;
    assign in8172_1 = {pp33[11]};
    assign in8172_2 = {pp34[10]};
    Full_Adder FA_8172(s8172, c8172, in8172_1, in8172_2, pp32[12]);
    wire[0:0] s8173, in8173_1, in8173_2;
    wire c8173;
    assign in8173_1 = {pp36[8]};
    assign in8173_2 = {pp37[7]};
    Full_Adder FA_8173(s8173, c8173, in8173_1, in8173_2, pp35[9]);
    wire[0:0] s8174, in8174_1, in8174_2;
    wire c8174;
    assign in8174_1 = {pp39[5]};
    assign in8174_2 = {pp40[4]};
    Full_Adder FA_8174(s8174, c8174, in8174_1, in8174_2, pp38[6]);
    wire[0:0] s8175, in8175_1, in8175_2;
    wire c8175;
    assign in8175_1 = {pp42[2]};
    assign in8175_2 = {pp43[1]};
    Full_Adder FA_8175(s8175, c8175, in8175_1, in8175_2, pp41[3]);
    wire[0:0] s8176, in8176_1, in8176_2;
    wire c8176;
    assign in8176_1 = {c4981};
    assign in8176_2 = {c4982};
    Full_Adder FA_8176(s8176, c8176, in8176_1, in8176_2, pp44[0]);
    wire[0:0] s8177, in8177_1, in8177_2;
    wire c8177;
    assign in8177_1 = {c4984};
    assign in8177_2 = {c4985};
    Full_Adder FA_8177(s8177, c8177, in8177_1, in8177_2, c4983);
    wire[0:0] s8178, in8178_1, in8178_2;
    wire c8178;
    assign in8178_1 = {s4987[0]};
    assign in8178_2 = {s4988[0]};
    Full_Adder FA_8178(s8178, c8178, in8178_1, in8178_2, s4986[0]);
    wire[0:0] s8179, in8179_1, in8179_2;
    wire c8179;
    assign in8179_1 = {s4990[0]};
    assign in8179_2 = {s4991[0]};
    Full_Adder FA_8179(s8179, c8179, in8179_1, in8179_2, s4989[0]);
    wire[0:0] s8180, in8180_1, in8180_2;
    wire c8180;
    assign in8180_1 = {pp21[24]};
    assign in8180_2 = {pp22[23]};
    Full_Adder FA_8180(s8180, c8180, in8180_1, in8180_2, pp20[25]);
    wire[0:0] s8181, in8181_1, in8181_2;
    wire c8181;
    assign in8181_1 = {pp24[21]};
    assign in8181_2 = {pp25[20]};
    Full_Adder FA_8181(s8181, c8181, in8181_1, in8181_2, pp23[22]);
    wire[0:0] s8182, in8182_1, in8182_2;
    wire c8182;
    assign in8182_1 = {pp27[18]};
    assign in8182_2 = {pp28[17]};
    Full_Adder FA_8182(s8182, c8182, in8182_1, in8182_2, pp26[19]);
    wire[0:0] s8183, in8183_1, in8183_2;
    wire c8183;
    assign in8183_1 = {pp30[15]};
    assign in8183_2 = {pp31[14]};
    Full_Adder FA_8183(s8183, c8183, in8183_1, in8183_2, pp29[16]);
    wire[0:0] s8184, in8184_1, in8184_2;
    wire c8184;
    assign in8184_1 = {pp33[12]};
    assign in8184_2 = {pp34[11]};
    Full_Adder FA_8184(s8184, c8184, in8184_1, in8184_2, pp32[13]);
    wire[0:0] s8185, in8185_1, in8185_2;
    wire c8185;
    assign in8185_1 = {pp36[9]};
    assign in8185_2 = {pp37[8]};
    Full_Adder FA_8185(s8185, c8185, in8185_1, in8185_2, pp35[10]);
    wire[0:0] s8186, in8186_1, in8186_2;
    wire c8186;
    assign in8186_1 = {pp39[6]};
    assign in8186_2 = {pp40[5]};
    Full_Adder FA_8186(s8186, c8186, in8186_1, in8186_2, pp38[7]);
    wire[0:0] s8187, in8187_1, in8187_2;
    wire c8187;
    assign in8187_1 = {pp42[3]};
    assign in8187_2 = {pp43[2]};
    Full_Adder FA_8187(s8187, c8187, in8187_1, in8187_2, pp41[4]);
    wire[0:0] s8188, in8188_1, in8188_2;
    wire c8188;
    assign in8188_1 = {pp45[0]};
    assign in8188_2 = {c4986};
    Full_Adder FA_8188(s8188, c8188, in8188_1, in8188_2, pp44[1]);
    wire[0:0] s8189, in8189_1, in8189_2;
    wire c8189;
    assign in8189_1 = {c4988};
    assign in8189_2 = {c4989};
    Full_Adder FA_8189(s8189, c8189, in8189_1, in8189_2, c4987);
    wire[0:0] s8190, in8190_1, in8190_2;
    wire c8190;
    assign in8190_1 = {c4991};
    assign in8190_2 = {s4992[0]};
    Full_Adder FA_8190(s8190, c8190, in8190_1, in8190_2, c4990);
    wire[0:0] s8191, in8191_1, in8191_2;
    wire c8191;
    assign in8191_1 = {s4994[0]};
    assign in8191_2 = {s4995[0]};
    Full_Adder FA_8191(s8191, c8191, in8191_1, in8191_2, s4993[0]);
    wire[0:0] s8192, in8192_1, in8192_2;
    wire c8192;
    assign in8192_1 = {s4997[0]};
    assign in8192_2 = {s4998[0]};
    Full_Adder FA_8192(s8192, c8192, in8192_1, in8192_2, s4996[0]);
    wire[0:0] s8193, in8193_1, in8193_2;
    wire c8193;
    assign in8193_1 = {pp24[22]};
    assign in8193_2 = {pp25[21]};
    Full_Adder FA_8193(s8193, c8193, in8193_1, in8193_2, pp23[23]);
    wire[0:0] s8194, in8194_1, in8194_2;
    wire c8194;
    assign in8194_1 = {pp27[19]};
    assign in8194_2 = {pp28[18]};
    Full_Adder FA_8194(s8194, c8194, in8194_1, in8194_2, pp26[20]);
    wire[0:0] s8195, in8195_1, in8195_2;
    wire c8195;
    assign in8195_1 = {pp30[16]};
    assign in8195_2 = {pp31[15]};
    Full_Adder FA_8195(s8195, c8195, in8195_1, in8195_2, pp29[17]);
    wire[0:0] s8196, in8196_1, in8196_2;
    wire c8196;
    assign in8196_1 = {pp33[13]};
    assign in8196_2 = {pp34[12]};
    Full_Adder FA_8196(s8196, c8196, in8196_1, in8196_2, pp32[14]);
    wire[0:0] s8197, in8197_1, in8197_2;
    wire c8197;
    assign in8197_1 = {pp36[10]};
    assign in8197_2 = {pp37[9]};
    Full_Adder FA_8197(s8197, c8197, in8197_1, in8197_2, pp35[11]);
    wire[0:0] s8198, in8198_1, in8198_2;
    wire c8198;
    assign in8198_1 = {pp39[7]};
    assign in8198_2 = {pp40[6]};
    Full_Adder FA_8198(s8198, c8198, in8198_1, in8198_2, pp38[8]);
    wire[0:0] s8199, in8199_1, in8199_2;
    wire c8199;
    assign in8199_1 = {pp42[4]};
    assign in8199_2 = {pp43[3]};
    Full_Adder FA_8199(s8199, c8199, in8199_1, in8199_2, pp41[5]);
    wire[0:0] s8200, in8200_1, in8200_2;
    wire c8200;
    assign in8200_1 = {pp45[1]};
    assign in8200_2 = {pp46[0]};
    Full_Adder FA_8200(s8200, c8200, in8200_1, in8200_2, pp44[2]);
    wire[0:0] s8201, in8201_1, in8201_2;
    wire c8201;
    assign in8201_1 = {c4993};
    assign in8201_2 = {c4994};
    Full_Adder FA_8201(s8201, c8201, in8201_1, in8201_2, c4992);
    wire[0:0] s8202, in8202_1, in8202_2;
    wire c8202;
    assign in8202_1 = {c4996};
    assign in8202_2 = {c4997};
    Full_Adder FA_8202(s8202, c8202, in8202_1, in8202_2, c4995);
    wire[0:0] s8203, in8203_1, in8203_2;
    wire c8203;
    assign in8203_1 = {s4999[0]};
    assign in8203_2 = {s5000[0]};
    Full_Adder FA_8203(s8203, c8203, in8203_1, in8203_2, c4998);
    wire[0:0] s8204, in8204_1, in8204_2;
    wire c8204;
    assign in8204_1 = {s5002[0]};
    assign in8204_2 = {s5003[0]};
    Full_Adder FA_8204(s8204, c8204, in8204_1, in8204_2, s5001[0]);
    wire[0:0] s8205, in8205_1, in8205_2;
    wire c8205;
    assign in8205_1 = {s5005[0]};
    assign in8205_2 = {s5006[0]};
    Full_Adder FA_8205(s8205, c8205, in8205_1, in8205_2, s5004[0]);
    wire[0:0] s8206, in8206_1, in8206_2;
    wire c8206;
    assign in8206_1 = {pp27[20]};
    assign in8206_2 = {pp28[19]};
    Full_Adder FA_8206(s8206, c8206, in8206_1, in8206_2, pp26[21]);
    wire[0:0] s8207, in8207_1, in8207_2;
    wire c8207;
    assign in8207_1 = {pp30[17]};
    assign in8207_2 = {pp31[16]};
    Full_Adder FA_8207(s8207, c8207, in8207_1, in8207_2, pp29[18]);
    wire[0:0] s8208, in8208_1, in8208_2;
    wire c8208;
    assign in8208_1 = {pp33[14]};
    assign in8208_2 = {pp34[13]};
    Full_Adder FA_8208(s8208, c8208, in8208_1, in8208_2, pp32[15]);
    wire[0:0] s8209, in8209_1, in8209_2;
    wire c8209;
    assign in8209_1 = {pp36[11]};
    assign in8209_2 = {pp37[10]};
    Full_Adder FA_8209(s8209, c8209, in8209_1, in8209_2, pp35[12]);
    wire[0:0] s8210, in8210_1, in8210_2;
    wire c8210;
    assign in8210_1 = {pp39[8]};
    assign in8210_2 = {pp40[7]};
    Full_Adder FA_8210(s8210, c8210, in8210_1, in8210_2, pp38[9]);
    wire[0:0] s8211, in8211_1, in8211_2;
    wire c8211;
    assign in8211_1 = {pp42[5]};
    assign in8211_2 = {pp43[4]};
    Full_Adder FA_8211(s8211, c8211, in8211_1, in8211_2, pp41[6]);
    wire[0:0] s8212, in8212_1, in8212_2;
    wire c8212;
    assign in8212_1 = {pp45[2]};
    assign in8212_2 = {pp46[1]};
    Full_Adder FA_8212(s8212, c8212, in8212_1, in8212_2, pp44[3]);
    wire[0:0] s8213, in8213_1, in8213_2;
    wire c8213;
    assign in8213_1 = {c4999};
    assign in8213_2 = {c5000};
    Full_Adder FA_8213(s8213, c8213, in8213_1, in8213_2, pp47[0]);
    wire[0:0] s8214, in8214_1, in8214_2;
    wire c8214;
    assign in8214_1 = {c5002};
    assign in8214_2 = {c5003};
    Full_Adder FA_8214(s8214, c8214, in8214_1, in8214_2, c5001);
    wire[0:0] s8215, in8215_1, in8215_2;
    wire c8215;
    assign in8215_1 = {c5005};
    assign in8215_2 = {c5006};
    Full_Adder FA_8215(s8215, c8215, in8215_1, in8215_2, c5004);
    wire[0:0] s8216, in8216_1, in8216_2;
    wire c8216;
    assign in8216_1 = {s5008[0]};
    assign in8216_2 = {s5009[0]};
    Full_Adder FA_8216(s8216, c8216, in8216_1, in8216_2, s5007[0]);
    wire[0:0] s8217, in8217_1, in8217_2;
    wire c8217;
    assign in8217_1 = {s5011[0]};
    assign in8217_2 = {s5012[0]};
    Full_Adder FA_8217(s8217, c8217, in8217_1, in8217_2, s5010[0]);
    wire[0:0] s8218, in8218_1, in8218_2;
    wire c8218;
    assign in8218_1 = {s5014[0]};
    assign in8218_2 = {s5015[0]};
    Full_Adder FA_8218(s8218, c8218, in8218_1, in8218_2, s5013[0]);
    wire[0:0] s8219, in8219_1, in8219_2;
    wire c8219;
    assign in8219_1 = {pp30[18]};
    assign in8219_2 = {pp31[17]};
    Full_Adder FA_8219(s8219, c8219, in8219_1, in8219_2, pp29[19]);
    wire[0:0] s8220, in8220_1, in8220_2;
    wire c8220;
    assign in8220_1 = {pp33[15]};
    assign in8220_2 = {pp34[14]};
    Full_Adder FA_8220(s8220, c8220, in8220_1, in8220_2, pp32[16]);
    wire[0:0] s8221, in8221_1, in8221_2;
    wire c8221;
    assign in8221_1 = {pp36[12]};
    assign in8221_2 = {pp37[11]};
    Full_Adder FA_8221(s8221, c8221, in8221_1, in8221_2, pp35[13]);
    wire[0:0] s8222, in8222_1, in8222_2;
    wire c8222;
    assign in8222_1 = {pp39[9]};
    assign in8222_2 = {pp40[8]};
    Full_Adder FA_8222(s8222, c8222, in8222_1, in8222_2, pp38[10]);
    wire[0:0] s8223, in8223_1, in8223_2;
    wire c8223;
    assign in8223_1 = {pp42[6]};
    assign in8223_2 = {pp43[5]};
    Full_Adder FA_8223(s8223, c8223, in8223_1, in8223_2, pp41[7]);
    wire[0:0] s8224, in8224_1, in8224_2;
    wire c8224;
    assign in8224_1 = {pp45[3]};
    assign in8224_2 = {pp46[2]};
    Full_Adder FA_8224(s8224, c8224, in8224_1, in8224_2, pp44[4]);
    wire[0:0] s8225, in8225_1, in8225_2;
    wire c8225;
    assign in8225_1 = {pp48[0]};
    assign in8225_2 = {c5007};
    Full_Adder FA_8225(s8225, c8225, in8225_1, in8225_2, pp47[1]);
    wire[0:0] s8226, in8226_1, in8226_2;
    wire c8226;
    assign in8226_1 = {c5009};
    assign in8226_2 = {c5010};
    Full_Adder FA_8226(s8226, c8226, in8226_1, in8226_2, c5008);
    wire[0:0] s8227, in8227_1, in8227_2;
    wire c8227;
    assign in8227_1 = {c5012};
    assign in8227_2 = {c5013};
    Full_Adder FA_8227(s8227, c8227, in8227_1, in8227_2, c5011);
    wire[0:0] s8228, in8228_1, in8228_2;
    wire c8228;
    assign in8228_1 = {c5015};
    assign in8228_2 = {s5016[0]};
    Full_Adder FA_8228(s8228, c8228, in8228_1, in8228_2, c5014);
    wire[0:0] s8229, in8229_1, in8229_2;
    wire c8229;
    assign in8229_1 = {s5018[0]};
    assign in8229_2 = {s5019[0]};
    Full_Adder FA_8229(s8229, c8229, in8229_1, in8229_2, s5017[0]);
    wire[0:0] s8230, in8230_1, in8230_2;
    wire c8230;
    assign in8230_1 = {s5021[0]};
    assign in8230_2 = {s5022[0]};
    Full_Adder FA_8230(s8230, c8230, in8230_1, in8230_2, s5020[0]);
    wire[0:0] s8231, in8231_1, in8231_2;
    wire c8231;
    assign in8231_1 = {s5024[0]};
    assign in8231_2 = {s5025[0]};
    Full_Adder FA_8231(s8231, c8231, in8231_1, in8231_2, s5023[0]);
    wire[0:0] s8232, in8232_1, in8232_2;
    wire c8232;
    assign in8232_1 = {pp33[16]};
    assign in8232_2 = {pp34[15]};
    Full_Adder FA_8232(s8232, c8232, in8232_1, in8232_2, pp32[17]);
    wire[0:0] s8233, in8233_1, in8233_2;
    wire c8233;
    assign in8233_1 = {pp36[13]};
    assign in8233_2 = {pp37[12]};
    Full_Adder FA_8233(s8233, c8233, in8233_1, in8233_2, pp35[14]);
    wire[0:0] s8234, in8234_1, in8234_2;
    wire c8234;
    assign in8234_1 = {pp39[10]};
    assign in8234_2 = {pp40[9]};
    Full_Adder FA_8234(s8234, c8234, in8234_1, in8234_2, pp38[11]);
    wire[0:0] s8235, in8235_1, in8235_2;
    wire c8235;
    assign in8235_1 = {pp42[7]};
    assign in8235_2 = {pp43[6]};
    Full_Adder FA_8235(s8235, c8235, in8235_1, in8235_2, pp41[8]);
    wire[0:0] s8236, in8236_1, in8236_2;
    wire c8236;
    assign in8236_1 = {pp45[4]};
    assign in8236_2 = {pp46[3]};
    Full_Adder FA_8236(s8236, c8236, in8236_1, in8236_2, pp44[5]);
    wire[0:0] s8237, in8237_1, in8237_2;
    wire c8237;
    assign in8237_1 = {pp48[1]};
    assign in8237_2 = {pp49[0]};
    Full_Adder FA_8237(s8237, c8237, in8237_1, in8237_2, pp47[2]);
    wire[0:0] s8238, in8238_1, in8238_2;
    wire c8238;
    assign in8238_1 = {c5017};
    assign in8238_2 = {c5018};
    Full_Adder FA_8238(s8238, c8238, in8238_1, in8238_2, c5016);
    wire[0:0] s8239, in8239_1, in8239_2;
    wire c8239;
    assign in8239_1 = {c5020};
    assign in8239_2 = {c5021};
    Full_Adder FA_8239(s8239, c8239, in8239_1, in8239_2, c5019);
    wire[0:0] s8240, in8240_1, in8240_2;
    wire c8240;
    assign in8240_1 = {c5023};
    assign in8240_2 = {c5024};
    Full_Adder FA_8240(s8240, c8240, in8240_1, in8240_2, c5022);
    wire[0:0] s8241, in8241_1, in8241_2;
    wire c8241;
    assign in8241_1 = {s5026[0]};
    assign in8241_2 = {s5027[0]};
    Full_Adder FA_8241(s8241, c8241, in8241_1, in8241_2, c5025);
    wire[0:0] s8242, in8242_1, in8242_2;
    wire c8242;
    assign in8242_1 = {s5029[0]};
    assign in8242_2 = {s5030[0]};
    Full_Adder FA_8242(s8242, c8242, in8242_1, in8242_2, s5028[0]);
    wire[0:0] s8243, in8243_1, in8243_2;
    wire c8243;
    assign in8243_1 = {s5032[0]};
    assign in8243_2 = {s5033[0]};
    Full_Adder FA_8243(s8243, c8243, in8243_1, in8243_2, s5031[0]);
    wire[0:0] s8244, in8244_1, in8244_2;
    wire c8244;
    assign in8244_1 = {s5035[0]};
    assign in8244_2 = {s5036[0]};
    Full_Adder FA_8244(s8244, c8244, in8244_1, in8244_2, s5034[0]);
    wire[0:0] s8245, in8245_1, in8245_2;
    wire c8245;
    assign in8245_1 = {pp36[14]};
    assign in8245_2 = {pp37[13]};
    Full_Adder FA_8245(s8245, c8245, in8245_1, in8245_2, pp35[15]);
    wire[0:0] s8246, in8246_1, in8246_2;
    wire c8246;
    assign in8246_1 = {pp39[11]};
    assign in8246_2 = {pp40[10]};
    Full_Adder FA_8246(s8246, c8246, in8246_1, in8246_2, pp38[12]);
    wire[0:0] s8247, in8247_1, in8247_2;
    wire c8247;
    assign in8247_1 = {pp42[8]};
    assign in8247_2 = {pp43[7]};
    Full_Adder FA_8247(s8247, c8247, in8247_1, in8247_2, pp41[9]);
    wire[0:0] s8248, in8248_1, in8248_2;
    wire c8248;
    assign in8248_1 = {pp45[5]};
    assign in8248_2 = {pp46[4]};
    Full_Adder FA_8248(s8248, c8248, in8248_1, in8248_2, pp44[6]);
    wire[0:0] s8249, in8249_1, in8249_2;
    wire c8249;
    assign in8249_1 = {pp48[2]};
    assign in8249_2 = {pp49[1]};
    Full_Adder FA_8249(s8249, c8249, in8249_1, in8249_2, pp47[3]);
    wire[0:0] s8250, in8250_1, in8250_2;
    wire c8250;
    assign in8250_1 = {c5026};
    assign in8250_2 = {c5027};
    Full_Adder FA_8250(s8250, c8250, in8250_1, in8250_2, pp50[0]);
    wire[0:0] s8251, in8251_1, in8251_2;
    wire c8251;
    assign in8251_1 = {c5029};
    assign in8251_2 = {c5030};
    Full_Adder FA_8251(s8251, c8251, in8251_1, in8251_2, c5028);
    wire[0:0] s8252, in8252_1, in8252_2;
    wire c8252;
    assign in8252_1 = {c5032};
    assign in8252_2 = {c5033};
    Full_Adder FA_8252(s8252, c8252, in8252_1, in8252_2, c5031);
    wire[0:0] s8253, in8253_1, in8253_2;
    wire c8253;
    assign in8253_1 = {c5035};
    assign in8253_2 = {c5036};
    Full_Adder FA_8253(s8253, c8253, in8253_1, in8253_2, c5034);
    wire[0:0] s8254, in8254_1, in8254_2;
    wire c8254;
    assign in8254_1 = {s5038[0]};
    assign in8254_2 = {s5039[0]};
    Full_Adder FA_8254(s8254, c8254, in8254_1, in8254_2, s5037[0]);
    wire[0:0] s8255, in8255_1, in8255_2;
    wire c8255;
    assign in8255_1 = {s5041[0]};
    assign in8255_2 = {s5042[0]};
    Full_Adder FA_8255(s8255, c8255, in8255_1, in8255_2, s5040[0]);
    wire[0:0] s8256, in8256_1, in8256_2;
    wire c8256;
    assign in8256_1 = {s5044[0]};
    assign in8256_2 = {s5045[0]};
    Full_Adder FA_8256(s8256, c8256, in8256_1, in8256_2, s5043[0]);
    wire[0:0] s8257, in8257_1, in8257_2;
    wire c8257;
    assign in8257_1 = {s5047[0]};
    assign in8257_2 = {s5048[0]};
    Full_Adder FA_8257(s8257, c8257, in8257_1, in8257_2, s5046[0]);
    wire[0:0] s8258, in8258_1, in8258_2;
    wire c8258;
    assign in8258_1 = {pp39[12]};
    assign in8258_2 = {pp40[11]};
    Full_Adder FA_8258(s8258, c8258, in8258_1, in8258_2, pp38[13]);
    wire[0:0] s8259, in8259_1, in8259_2;
    wire c8259;
    assign in8259_1 = {pp42[9]};
    assign in8259_2 = {pp43[8]};
    Full_Adder FA_8259(s8259, c8259, in8259_1, in8259_2, pp41[10]);
    wire[0:0] s8260, in8260_1, in8260_2;
    wire c8260;
    assign in8260_1 = {pp45[6]};
    assign in8260_2 = {pp46[5]};
    Full_Adder FA_8260(s8260, c8260, in8260_1, in8260_2, pp44[7]);
    wire[0:0] s8261, in8261_1, in8261_2;
    wire c8261;
    assign in8261_1 = {pp48[3]};
    assign in8261_2 = {pp49[2]};
    Full_Adder FA_8261(s8261, c8261, in8261_1, in8261_2, pp47[4]);
    wire[0:0] s8262, in8262_1, in8262_2;
    wire c8262;
    assign in8262_1 = {pp51[0]};
    assign in8262_2 = {c5037};
    Full_Adder FA_8262(s8262, c8262, in8262_1, in8262_2, pp50[1]);
    wire[0:0] s8263, in8263_1, in8263_2;
    wire c8263;
    assign in8263_1 = {c5039};
    assign in8263_2 = {c5040};
    Full_Adder FA_8263(s8263, c8263, in8263_1, in8263_2, c5038);
    wire[0:0] s8264, in8264_1, in8264_2;
    wire c8264;
    assign in8264_1 = {c5042};
    assign in8264_2 = {c5043};
    Full_Adder FA_8264(s8264, c8264, in8264_1, in8264_2, c5041);
    wire[0:0] s8265, in8265_1, in8265_2;
    wire c8265;
    assign in8265_1 = {c5045};
    assign in8265_2 = {c5046};
    Full_Adder FA_8265(s8265, c8265, in8265_1, in8265_2, c5044);
    wire[0:0] s8266, in8266_1, in8266_2;
    wire c8266;
    assign in8266_1 = {c5048};
    assign in8266_2 = {s5049[0]};
    Full_Adder FA_8266(s8266, c8266, in8266_1, in8266_2, c5047);
    wire[0:0] s8267, in8267_1, in8267_2;
    wire c8267;
    assign in8267_1 = {s5051[0]};
    assign in8267_2 = {s5052[0]};
    Full_Adder FA_8267(s8267, c8267, in8267_1, in8267_2, s5050[0]);
    wire[0:0] s8268, in8268_1, in8268_2;
    wire c8268;
    assign in8268_1 = {s5054[0]};
    assign in8268_2 = {s5055[0]};
    Full_Adder FA_8268(s8268, c8268, in8268_1, in8268_2, s5053[0]);
    wire[0:0] s8269, in8269_1, in8269_2;
    wire c8269;
    assign in8269_1 = {s5057[0]};
    assign in8269_2 = {s5058[0]};
    Full_Adder FA_8269(s8269, c8269, in8269_1, in8269_2, s5056[0]);
    wire[0:0] s8270, in8270_1, in8270_2;
    wire c8270;
    assign in8270_1 = {s5060[0]};
    assign in8270_2 = {s5061[0]};
    Full_Adder FA_8270(s8270, c8270, in8270_1, in8270_2, s5059[0]);
    wire[0:0] s8271, in8271_1, in8271_2;
    wire c8271;
    assign in8271_1 = {pp42[10]};
    assign in8271_2 = {pp43[9]};
    Full_Adder FA_8271(s8271, c8271, in8271_1, in8271_2, pp41[11]);
    wire[0:0] s8272, in8272_1, in8272_2;
    wire c8272;
    assign in8272_1 = {pp45[7]};
    assign in8272_2 = {pp46[6]};
    Full_Adder FA_8272(s8272, c8272, in8272_1, in8272_2, pp44[8]);
    wire[0:0] s8273, in8273_1, in8273_2;
    wire c8273;
    assign in8273_1 = {pp48[4]};
    assign in8273_2 = {pp49[3]};
    Full_Adder FA_8273(s8273, c8273, in8273_1, in8273_2, pp47[5]);
    wire[0:0] s8274, in8274_1, in8274_2;
    wire c8274;
    assign in8274_1 = {pp51[1]};
    assign in8274_2 = {pp52[0]};
    Full_Adder FA_8274(s8274, c8274, in8274_1, in8274_2, pp50[2]);
    wire[0:0] s8275, in8275_1, in8275_2;
    wire c8275;
    assign in8275_1 = {c5050};
    assign in8275_2 = {c5051};
    Full_Adder FA_8275(s8275, c8275, in8275_1, in8275_2, c5049);
    wire[0:0] s8276, in8276_1, in8276_2;
    wire c8276;
    assign in8276_1 = {c5053};
    assign in8276_2 = {c5054};
    Full_Adder FA_8276(s8276, c8276, in8276_1, in8276_2, c5052);
    wire[0:0] s8277, in8277_1, in8277_2;
    wire c8277;
    assign in8277_1 = {c5056};
    assign in8277_2 = {c5057};
    Full_Adder FA_8277(s8277, c8277, in8277_1, in8277_2, c5055);
    wire[0:0] s8278, in8278_1, in8278_2;
    wire c8278;
    assign in8278_1 = {c5059};
    assign in8278_2 = {c5060};
    Full_Adder FA_8278(s8278, c8278, in8278_1, in8278_2, c5058);
    wire[0:0] s8279, in8279_1, in8279_2;
    wire c8279;
    assign in8279_1 = {s5062[0]};
    assign in8279_2 = {s5063[0]};
    Full_Adder FA_8279(s8279, c8279, in8279_1, in8279_2, c5061);
    wire[0:0] s8280, in8280_1, in8280_2;
    wire c8280;
    assign in8280_1 = {s5065[0]};
    assign in8280_2 = {s5066[0]};
    Full_Adder FA_8280(s8280, c8280, in8280_1, in8280_2, s5064[0]);
    wire[0:0] s8281, in8281_1, in8281_2;
    wire c8281;
    assign in8281_1 = {s5068[0]};
    assign in8281_2 = {s5069[0]};
    Full_Adder FA_8281(s8281, c8281, in8281_1, in8281_2, s5067[0]);
    wire[0:0] s8282, in8282_1, in8282_2;
    wire c8282;
    assign in8282_1 = {s5071[0]};
    assign in8282_2 = {s5072[0]};
    Full_Adder FA_8282(s8282, c8282, in8282_1, in8282_2, s5070[0]);
    wire[0:0] s8283, in8283_1, in8283_2;
    wire c8283;
    assign in8283_1 = {s5074[0]};
    assign in8283_2 = {s5075[0]};
    Full_Adder FA_8283(s8283, c8283, in8283_1, in8283_2, s5073[0]);
    wire[0:0] s8284, in8284_1, in8284_2;
    wire c8284;
    assign in8284_1 = {pp45[8]};
    assign in8284_2 = {pp46[7]};
    Full_Adder FA_8284(s8284, c8284, in8284_1, in8284_2, pp44[9]);
    wire[0:0] s8285, in8285_1, in8285_2;
    wire c8285;
    assign in8285_1 = {pp48[5]};
    assign in8285_2 = {pp49[4]};
    Full_Adder FA_8285(s8285, c8285, in8285_1, in8285_2, pp47[6]);
    wire[0:0] s8286, in8286_1, in8286_2;
    wire c8286;
    assign in8286_1 = {pp51[2]};
    assign in8286_2 = {pp52[1]};
    Full_Adder FA_8286(s8286, c8286, in8286_1, in8286_2, pp50[3]);
    wire[0:0] s8287, in8287_1, in8287_2;
    wire c8287;
    assign in8287_1 = {c5062};
    assign in8287_2 = {c5063};
    Full_Adder FA_8287(s8287, c8287, in8287_1, in8287_2, pp53[0]);
    wire[0:0] s8288, in8288_1, in8288_2;
    wire c8288;
    assign in8288_1 = {c5065};
    assign in8288_2 = {c5066};
    Full_Adder FA_8288(s8288, c8288, in8288_1, in8288_2, c5064);
    wire[0:0] s8289, in8289_1, in8289_2;
    wire c8289;
    assign in8289_1 = {c5068};
    assign in8289_2 = {c5069};
    Full_Adder FA_8289(s8289, c8289, in8289_1, in8289_2, c5067);
    wire[0:0] s8290, in8290_1, in8290_2;
    wire c8290;
    assign in8290_1 = {c5071};
    assign in8290_2 = {c5072};
    Full_Adder FA_8290(s8290, c8290, in8290_1, in8290_2, c5070);
    wire[0:0] s8291, in8291_1, in8291_2;
    wire c8291;
    assign in8291_1 = {c5074};
    assign in8291_2 = {c5075};
    Full_Adder FA_8291(s8291, c8291, in8291_1, in8291_2, c5073);
    wire[0:0] s8292, in8292_1, in8292_2;
    wire c8292;
    assign in8292_1 = {s5077[0]};
    assign in8292_2 = {s5078[0]};
    Full_Adder FA_8292(s8292, c8292, in8292_1, in8292_2, s5076[0]);
    wire[0:0] s8293, in8293_1, in8293_2;
    wire c8293;
    assign in8293_1 = {s5080[0]};
    assign in8293_2 = {s5081[0]};
    Full_Adder FA_8293(s8293, c8293, in8293_1, in8293_2, s5079[0]);
    wire[0:0] s8294, in8294_1, in8294_2;
    wire c8294;
    assign in8294_1 = {s5083[0]};
    assign in8294_2 = {s5084[0]};
    Full_Adder FA_8294(s8294, c8294, in8294_1, in8294_2, s5082[0]);
    wire[0:0] s8295, in8295_1, in8295_2;
    wire c8295;
    assign in8295_1 = {s5086[0]};
    assign in8295_2 = {s5087[0]};
    Full_Adder FA_8295(s8295, c8295, in8295_1, in8295_2, s5085[0]);
    wire[0:0] s8296, in8296_1, in8296_2;
    wire c8296;
    assign in8296_1 = {s5089[0]};
    assign in8296_2 = {s5090[0]};
    Full_Adder FA_8296(s8296, c8296, in8296_1, in8296_2, s5088[0]);
    wire[0:0] s8297, in8297_1, in8297_2;
    wire c8297;
    assign in8297_1 = {pp48[6]};
    assign in8297_2 = {pp49[5]};
    Full_Adder FA_8297(s8297, c8297, in8297_1, in8297_2, pp47[7]);
    wire[0:0] s8298, in8298_1, in8298_2;
    wire c8298;
    assign in8298_1 = {pp51[3]};
    assign in8298_2 = {pp52[2]};
    Full_Adder FA_8298(s8298, c8298, in8298_1, in8298_2, pp50[4]);
    wire[0:0] s8299, in8299_1, in8299_2;
    wire c8299;
    assign in8299_1 = {pp54[0]};
    assign in8299_2 = {c5076};
    Full_Adder FA_8299(s8299, c8299, in8299_1, in8299_2, pp53[1]);
    wire[0:0] s8300, in8300_1, in8300_2;
    wire c8300;
    assign in8300_1 = {c5078};
    assign in8300_2 = {c5079};
    Full_Adder FA_8300(s8300, c8300, in8300_1, in8300_2, c5077);
    wire[0:0] s8301, in8301_1, in8301_2;
    wire c8301;
    assign in8301_1 = {c5081};
    assign in8301_2 = {c5082};
    Full_Adder FA_8301(s8301, c8301, in8301_1, in8301_2, c5080);
    wire[0:0] s8302, in8302_1, in8302_2;
    wire c8302;
    assign in8302_1 = {c5084};
    assign in8302_2 = {c5085};
    Full_Adder FA_8302(s8302, c8302, in8302_1, in8302_2, c5083);
    wire[0:0] s8303, in8303_1, in8303_2;
    wire c8303;
    assign in8303_1 = {c5087};
    assign in8303_2 = {c5088};
    Full_Adder FA_8303(s8303, c8303, in8303_1, in8303_2, c5086);
    wire[0:0] s8304, in8304_1, in8304_2;
    wire c8304;
    assign in8304_1 = {c5090};
    assign in8304_2 = {s5091[0]};
    Full_Adder FA_8304(s8304, c8304, in8304_1, in8304_2, c5089);
    wire[0:0] s8305, in8305_1, in8305_2;
    wire c8305;
    assign in8305_1 = {s5093[0]};
    assign in8305_2 = {s5094[0]};
    Full_Adder FA_8305(s8305, c8305, in8305_1, in8305_2, s5092[0]);
    wire[0:0] s8306, in8306_1, in8306_2;
    wire c8306;
    assign in8306_1 = {s5096[0]};
    assign in8306_2 = {s5097[0]};
    Full_Adder FA_8306(s8306, c8306, in8306_1, in8306_2, s5095[0]);
    wire[0:0] s8307, in8307_1, in8307_2;
    wire c8307;
    assign in8307_1 = {s5099[0]};
    assign in8307_2 = {s5100[0]};
    Full_Adder FA_8307(s8307, c8307, in8307_1, in8307_2, s5098[0]);
    wire[0:0] s8308, in8308_1, in8308_2;
    wire c8308;
    assign in8308_1 = {s5102[0]};
    assign in8308_2 = {s5103[0]};
    Full_Adder FA_8308(s8308, c8308, in8308_1, in8308_2, s5101[0]);
    wire[0:0] s8309, in8309_1, in8309_2;
    wire c8309;
    assign in8309_1 = {s5105[0]};
    assign in8309_2 = {s5106[0]};
    Full_Adder FA_8309(s8309, c8309, in8309_1, in8309_2, s5104[0]);
    wire[0:0] s8310, in8310_1, in8310_2;
    wire c8310;
    assign in8310_1 = {pp51[4]};
    assign in8310_2 = {pp52[3]};
    Full_Adder FA_8310(s8310, c8310, in8310_1, in8310_2, pp50[5]);
    wire[0:0] s8311, in8311_1, in8311_2;
    wire c8311;
    assign in8311_1 = {pp54[1]};
    assign in8311_2 = {pp55[0]};
    Full_Adder FA_8311(s8311, c8311, in8311_1, in8311_2, pp53[2]);
    wire[0:0] s8312, in8312_1, in8312_2;
    wire c8312;
    assign in8312_1 = {c5092};
    assign in8312_2 = {c5093};
    Full_Adder FA_8312(s8312, c8312, in8312_1, in8312_2, c5091);
    wire[0:0] s8313, in8313_1, in8313_2;
    wire c8313;
    assign in8313_1 = {c5095};
    assign in8313_2 = {c5096};
    Full_Adder FA_8313(s8313, c8313, in8313_1, in8313_2, c5094);
    wire[0:0] s8314, in8314_1, in8314_2;
    wire c8314;
    assign in8314_1 = {c5098};
    assign in8314_2 = {c5099};
    Full_Adder FA_8314(s8314, c8314, in8314_1, in8314_2, c5097);
    wire[0:0] s8315, in8315_1, in8315_2;
    wire c8315;
    assign in8315_1 = {c5101};
    assign in8315_2 = {c5102};
    Full_Adder FA_8315(s8315, c8315, in8315_1, in8315_2, c5100);
    wire[0:0] s8316, in8316_1, in8316_2;
    wire c8316;
    assign in8316_1 = {c5104};
    assign in8316_2 = {c5105};
    Full_Adder FA_8316(s8316, c8316, in8316_1, in8316_2, c5103);
    wire[0:0] s8317, in8317_1, in8317_2;
    wire c8317;
    assign in8317_1 = {s5107[0]};
    assign in8317_2 = {s5108[0]};
    Full_Adder FA_8317(s8317, c8317, in8317_1, in8317_2, c5106);
    wire[0:0] s8318, in8318_1, in8318_2;
    wire c8318;
    assign in8318_1 = {s5110[0]};
    assign in8318_2 = {s5111[0]};
    Full_Adder FA_8318(s8318, c8318, in8318_1, in8318_2, s5109[0]);
    wire[0:0] s8319, in8319_1, in8319_2;
    wire c8319;
    assign in8319_1 = {s5113[0]};
    assign in8319_2 = {s5114[0]};
    Full_Adder FA_8319(s8319, c8319, in8319_1, in8319_2, s5112[0]);
    wire[0:0] s8320, in8320_1, in8320_2;
    wire c8320;
    assign in8320_1 = {s5116[0]};
    assign in8320_2 = {s5117[0]};
    Full_Adder FA_8320(s8320, c8320, in8320_1, in8320_2, s5115[0]);
    wire[0:0] s8321, in8321_1, in8321_2;
    wire c8321;
    assign in8321_1 = {s5119[0]};
    assign in8321_2 = {s5120[0]};
    Full_Adder FA_8321(s8321, c8321, in8321_1, in8321_2, s5118[0]);
    wire[0:0] s8322, in8322_1, in8322_2;
    wire c8322;
    assign in8322_1 = {s5122[0]};
    assign in8322_2 = {s5123[0]};
    Full_Adder FA_8322(s8322, c8322, in8322_1, in8322_2, s5121[0]);
    wire[0:0] s8323, in8323_1, in8323_2;
    wire c8323;
    assign in8323_1 = {pp54[2]};
    assign in8323_2 = {pp55[1]};
    Full_Adder FA_8323(s8323, c8323, in8323_1, in8323_2, pp53[3]);
    wire[0:0] s8324, in8324_1, in8324_2;
    wire c8324;
    assign in8324_1 = {c5107};
    assign in8324_2 = {c5108};
    Full_Adder FA_8324(s8324, c8324, in8324_1, in8324_2, pp56[0]);
    wire[0:0] s8325, in8325_1, in8325_2;
    wire c8325;
    assign in8325_1 = {c5110};
    assign in8325_2 = {c5111};
    Full_Adder FA_8325(s8325, c8325, in8325_1, in8325_2, c5109);
    wire[0:0] s8326, in8326_1, in8326_2;
    wire c8326;
    assign in8326_1 = {c5113};
    assign in8326_2 = {c5114};
    Full_Adder FA_8326(s8326, c8326, in8326_1, in8326_2, c5112);
    wire[0:0] s8327, in8327_1, in8327_2;
    wire c8327;
    assign in8327_1 = {c5116};
    assign in8327_2 = {c5117};
    Full_Adder FA_8327(s8327, c8327, in8327_1, in8327_2, c5115);
    wire[0:0] s8328, in8328_1, in8328_2;
    wire c8328;
    assign in8328_1 = {c5119};
    assign in8328_2 = {c5120};
    Full_Adder FA_8328(s8328, c8328, in8328_1, in8328_2, c5118);
    wire[0:0] s8329, in8329_1, in8329_2;
    wire c8329;
    assign in8329_1 = {c5122};
    assign in8329_2 = {c5123};
    Full_Adder FA_8329(s8329, c8329, in8329_1, in8329_2, c5121);
    wire[0:0] s8330, in8330_1, in8330_2;
    wire c8330;
    assign in8330_1 = {s5125[0]};
    assign in8330_2 = {s5126[0]};
    Full_Adder FA_8330(s8330, c8330, in8330_1, in8330_2, s5124[0]);
    wire[0:0] s8331, in8331_1, in8331_2;
    wire c8331;
    assign in8331_1 = {s5128[0]};
    assign in8331_2 = {s5129[0]};
    Full_Adder FA_8331(s8331, c8331, in8331_1, in8331_2, s5127[0]);
    wire[0:0] s8332, in8332_1, in8332_2;
    wire c8332;
    assign in8332_1 = {s5131[0]};
    assign in8332_2 = {s5132[0]};
    Full_Adder FA_8332(s8332, c8332, in8332_1, in8332_2, s5130[0]);
    wire[0:0] s8333, in8333_1, in8333_2;
    wire c8333;
    assign in8333_1 = {s5134[0]};
    assign in8333_2 = {s5135[0]};
    Full_Adder FA_8333(s8333, c8333, in8333_1, in8333_2, s5133[0]);
    wire[0:0] s8334, in8334_1, in8334_2;
    wire c8334;
    assign in8334_1 = {s5137[0]};
    assign in8334_2 = {s5138[0]};
    Full_Adder FA_8334(s8334, c8334, in8334_1, in8334_2, s5136[0]);
    wire[0:0] s8335, in8335_1, in8335_2;
    wire c8335;
    assign in8335_1 = {s5140[0]};
    assign in8335_2 = {s5141[0]};
    Full_Adder FA_8335(s8335, c8335, in8335_1, in8335_2, s5139[0]);
    wire[0:0] s8336, in8336_1, in8336_2;
    wire c8336;
    assign in8336_1 = {pp57[0]};
    assign in8336_2 = {c5124};
    Full_Adder FA_8336(s8336, c8336, in8336_1, in8336_2, pp56[1]);
    wire[0:0] s8337, in8337_1, in8337_2;
    wire c8337;
    assign in8337_1 = {c5126};
    assign in8337_2 = {c5127};
    Full_Adder FA_8337(s8337, c8337, in8337_1, in8337_2, c5125);
    wire[0:0] s8338, in8338_1, in8338_2;
    wire c8338;
    assign in8338_1 = {c5129};
    assign in8338_2 = {c5130};
    Full_Adder FA_8338(s8338, c8338, in8338_1, in8338_2, c5128);
    wire[0:0] s8339, in8339_1, in8339_2;
    wire c8339;
    assign in8339_1 = {c5132};
    assign in8339_2 = {c5133};
    Full_Adder FA_8339(s8339, c8339, in8339_1, in8339_2, c5131);
    wire[0:0] s8340, in8340_1, in8340_2;
    wire c8340;
    assign in8340_1 = {c5135};
    assign in8340_2 = {c5136};
    Full_Adder FA_8340(s8340, c8340, in8340_1, in8340_2, c5134);
    wire[0:0] s8341, in8341_1, in8341_2;
    wire c8341;
    assign in8341_1 = {c5138};
    assign in8341_2 = {c5139};
    Full_Adder FA_8341(s8341, c8341, in8341_1, in8341_2, c5137);
    wire[0:0] s8342, in8342_1, in8342_2;
    wire c8342;
    assign in8342_1 = {c5141};
    assign in8342_2 = {s5142[0]};
    Full_Adder FA_8342(s8342, c8342, in8342_1, in8342_2, c5140);
    wire[0:0] s8343, in8343_1, in8343_2;
    wire c8343;
    assign in8343_1 = {s5144[0]};
    assign in8343_2 = {s5145[0]};
    Full_Adder FA_8343(s8343, c8343, in8343_1, in8343_2, s5143[0]);
    wire[0:0] s8344, in8344_1, in8344_2;
    wire c8344;
    assign in8344_1 = {s5147[0]};
    assign in8344_2 = {s5148[0]};
    Full_Adder FA_8344(s8344, c8344, in8344_1, in8344_2, s5146[0]);
    wire[0:0] s8345, in8345_1, in8345_2;
    wire c8345;
    assign in8345_1 = {s5150[0]};
    assign in8345_2 = {s5151[0]};
    Full_Adder FA_8345(s8345, c8345, in8345_1, in8345_2, s5149[0]);
    wire[0:0] s8346, in8346_1, in8346_2;
    wire c8346;
    assign in8346_1 = {s5153[0]};
    assign in8346_2 = {s5154[0]};
    Full_Adder FA_8346(s8346, c8346, in8346_1, in8346_2, s5152[0]);
    wire[0:0] s8347, in8347_1, in8347_2;
    wire c8347;
    assign in8347_1 = {s5156[0]};
    assign in8347_2 = {s5157[0]};
    Full_Adder FA_8347(s8347, c8347, in8347_1, in8347_2, s5155[0]);
    wire[0:0] s8348, in8348_1, in8348_2;
    wire c8348;
    assign in8348_1 = {s5159[0]};
    assign in8348_2 = {s5160[0]};
    Full_Adder FA_8348(s8348, c8348, in8348_1, in8348_2, s5158[0]);
    wire[0:0] s8349, in8349_1, in8349_2;
    wire c8349;
    assign in8349_1 = {c5142};
    assign in8349_2 = {c5143};
    Full_Adder FA_8349(s8349, c8349, in8349_1, in8349_2, s1807[0]);
    wire[0:0] s8350, in8350_1, in8350_2;
    wire c8350;
    assign in8350_1 = {c5145};
    assign in8350_2 = {c5146};
    Full_Adder FA_8350(s8350, c8350, in8350_1, in8350_2, c5144);
    wire[0:0] s8351, in8351_1, in8351_2;
    wire c8351;
    assign in8351_1 = {c5148};
    assign in8351_2 = {c5149};
    Full_Adder FA_8351(s8351, c8351, in8351_1, in8351_2, c5147);
    wire[0:0] s8352, in8352_1, in8352_2;
    wire c8352;
    assign in8352_1 = {c5151};
    assign in8352_2 = {c5152};
    Full_Adder FA_8352(s8352, c8352, in8352_1, in8352_2, c5150);
    wire[0:0] s8353, in8353_1, in8353_2;
    wire c8353;
    assign in8353_1 = {c5154};
    assign in8353_2 = {c5155};
    Full_Adder FA_8353(s8353, c8353, in8353_1, in8353_2, c5153);
    wire[0:0] s8354, in8354_1, in8354_2;
    wire c8354;
    assign in8354_1 = {c5157};
    assign in8354_2 = {c5158};
    Full_Adder FA_8354(s8354, c8354, in8354_1, in8354_2, c5156);
    wire[0:0] s8355, in8355_1, in8355_2;
    wire c8355;
    assign in8355_1 = {c5160};
    assign in8355_2 = {s5161[0]};
    Full_Adder FA_8355(s8355, c8355, in8355_1, in8355_2, c5159);
    wire[0:0] s8356, in8356_1, in8356_2;
    wire c8356;
    assign in8356_1 = {s5163[0]};
    assign in8356_2 = {s5164[0]};
    Full_Adder FA_8356(s8356, c8356, in8356_1, in8356_2, s5162[0]);
    wire[0:0] s8357, in8357_1, in8357_2;
    wire c8357;
    assign in8357_1 = {s5166[0]};
    assign in8357_2 = {s5167[0]};
    Full_Adder FA_8357(s8357, c8357, in8357_1, in8357_2, s5165[0]);
    wire[0:0] s8358, in8358_1, in8358_2;
    wire c8358;
    assign in8358_1 = {s5169[0]};
    assign in8358_2 = {s5170[0]};
    Full_Adder FA_8358(s8358, c8358, in8358_1, in8358_2, s5168[0]);
    wire[0:0] s8359, in8359_1, in8359_2;
    wire c8359;
    assign in8359_1 = {s5172[0]};
    assign in8359_2 = {s5173[0]};
    Full_Adder FA_8359(s8359, c8359, in8359_1, in8359_2, s5171[0]);
    wire[0:0] s8360, in8360_1, in8360_2;
    wire c8360;
    assign in8360_1 = {s5175[0]};
    assign in8360_2 = {s5176[0]};
    Full_Adder FA_8360(s8360, c8360, in8360_1, in8360_2, s5174[0]);
    wire[0:0] s8361, in8361_1, in8361_2;
    wire c8361;
    assign in8361_1 = {s5178[0]};
    assign in8361_2 = {s5179[0]};
    Full_Adder FA_8361(s8361, c8361, in8361_1, in8361_2, s5177[0]);
    wire[0:0] s8362, in8362_1, in8362_2;
    wire c8362;
    assign in8362_1 = {c5161};
    assign in8362_2 = {c5162};
    Full_Adder FA_8362(s8362, c8362, in8362_1, in8362_2, s1809[0]);
    wire[0:0] s8363, in8363_1, in8363_2;
    wire c8363;
    assign in8363_1 = {c5164};
    assign in8363_2 = {c5165};
    Full_Adder FA_8363(s8363, c8363, in8363_1, in8363_2, c5163);
    wire[0:0] s8364, in8364_1, in8364_2;
    wire c8364;
    assign in8364_1 = {c5167};
    assign in8364_2 = {c5168};
    Full_Adder FA_8364(s8364, c8364, in8364_1, in8364_2, c5166);
    wire[0:0] s8365, in8365_1, in8365_2;
    wire c8365;
    assign in8365_1 = {c5170};
    assign in8365_2 = {c5171};
    Full_Adder FA_8365(s8365, c8365, in8365_1, in8365_2, c5169);
    wire[0:0] s8366, in8366_1, in8366_2;
    wire c8366;
    assign in8366_1 = {c5173};
    assign in8366_2 = {c5174};
    Full_Adder FA_8366(s8366, c8366, in8366_1, in8366_2, c5172);
    wire[0:0] s8367, in8367_1, in8367_2;
    wire c8367;
    assign in8367_1 = {c5176};
    assign in8367_2 = {c5177};
    Full_Adder FA_8367(s8367, c8367, in8367_1, in8367_2, c5175);
    wire[0:0] s8368, in8368_1, in8368_2;
    wire c8368;
    assign in8368_1 = {c5179};
    assign in8368_2 = {s5180[0]};
    Full_Adder FA_8368(s8368, c8368, in8368_1, in8368_2, c5178);
    wire[0:0] s8369, in8369_1, in8369_2;
    wire c8369;
    assign in8369_1 = {s5182[0]};
    assign in8369_2 = {s5183[0]};
    Full_Adder FA_8369(s8369, c8369, in8369_1, in8369_2, s5181[0]);
    wire[0:0] s8370, in8370_1, in8370_2;
    wire c8370;
    assign in8370_1 = {s5185[0]};
    assign in8370_2 = {s5186[0]};
    Full_Adder FA_8370(s8370, c8370, in8370_1, in8370_2, s5184[0]);
    wire[0:0] s8371, in8371_1, in8371_2;
    wire c8371;
    assign in8371_1 = {s5188[0]};
    assign in8371_2 = {s5189[0]};
    Full_Adder FA_8371(s8371, c8371, in8371_1, in8371_2, s5187[0]);
    wire[0:0] s8372, in8372_1, in8372_2;
    wire c8372;
    assign in8372_1 = {s5191[0]};
    assign in8372_2 = {s5192[0]};
    Full_Adder FA_8372(s8372, c8372, in8372_1, in8372_2, s5190[0]);
    wire[0:0] s8373, in8373_1, in8373_2;
    wire c8373;
    assign in8373_1 = {s5194[0]};
    assign in8373_2 = {s5195[0]};
    Full_Adder FA_8373(s8373, c8373, in8373_1, in8373_2, s5193[0]);
    wire[0:0] s8374, in8374_1, in8374_2;
    wire c8374;
    assign in8374_1 = {s5197[0]};
    assign in8374_2 = {s5198[0]};
    Full_Adder FA_8374(s8374, c8374, in8374_1, in8374_2, s5196[0]);
    wire[0:0] s8375, in8375_1, in8375_2;
    wire c8375;
    assign in8375_1 = {c5180};
    assign in8375_2 = {c5181};
    Full_Adder FA_8375(s8375, c8375, in8375_1, in8375_2, s1812[0]);
    wire[0:0] s8376, in8376_1, in8376_2;
    wire c8376;
    assign in8376_1 = {c5183};
    assign in8376_2 = {c5184};
    Full_Adder FA_8376(s8376, c8376, in8376_1, in8376_2, c5182);
    wire[0:0] s8377, in8377_1, in8377_2;
    wire c8377;
    assign in8377_1 = {c5186};
    assign in8377_2 = {c5187};
    Full_Adder FA_8377(s8377, c8377, in8377_1, in8377_2, c5185);
    wire[0:0] s8378, in8378_1, in8378_2;
    wire c8378;
    assign in8378_1 = {c5189};
    assign in8378_2 = {c5190};
    Full_Adder FA_8378(s8378, c8378, in8378_1, in8378_2, c5188);
    wire[0:0] s8379, in8379_1, in8379_2;
    wire c8379;
    assign in8379_1 = {c5192};
    assign in8379_2 = {c5193};
    Full_Adder FA_8379(s8379, c8379, in8379_1, in8379_2, c5191);
    wire[0:0] s8380, in8380_1, in8380_2;
    wire c8380;
    assign in8380_1 = {c5195};
    assign in8380_2 = {c5196};
    Full_Adder FA_8380(s8380, c8380, in8380_1, in8380_2, c5194);
    wire[0:0] s8381, in8381_1, in8381_2;
    wire c8381;
    assign in8381_1 = {c5198};
    assign in8381_2 = {s5199[0]};
    Full_Adder FA_8381(s8381, c8381, in8381_1, in8381_2, c5197);
    wire[0:0] s8382, in8382_1, in8382_2;
    wire c8382;
    assign in8382_1 = {s5201[0]};
    assign in8382_2 = {s5202[0]};
    Full_Adder FA_8382(s8382, c8382, in8382_1, in8382_2, s5200[0]);
    wire[0:0] s8383, in8383_1, in8383_2;
    wire c8383;
    assign in8383_1 = {s5204[0]};
    assign in8383_2 = {s5205[0]};
    Full_Adder FA_8383(s8383, c8383, in8383_1, in8383_2, s5203[0]);
    wire[0:0] s8384, in8384_1, in8384_2;
    wire c8384;
    assign in8384_1 = {s5207[0]};
    assign in8384_2 = {s5208[0]};
    Full_Adder FA_8384(s8384, c8384, in8384_1, in8384_2, s5206[0]);
    wire[0:0] s8385, in8385_1, in8385_2;
    wire c8385;
    assign in8385_1 = {s5210[0]};
    assign in8385_2 = {s5211[0]};
    Full_Adder FA_8385(s8385, c8385, in8385_1, in8385_2, s5209[0]);
    wire[0:0] s8386, in8386_1, in8386_2;
    wire c8386;
    assign in8386_1 = {s5213[0]};
    assign in8386_2 = {s5214[0]};
    Full_Adder FA_8386(s8386, c8386, in8386_1, in8386_2, s5212[0]);
    wire[0:0] s8387, in8387_1, in8387_2;
    wire c8387;
    assign in8387_1 = {s5216[0]};
    assign in8387_2 = {s5217[0]};
    Full_Adder FA_8387(s8387, c8387, in8387_1, in8387_2, s5215[0]);
    wire[0:0] s8388, in8388_1, in8388_2;
    wire c8388;
    assign in8388_1 = {c5199};
    assign in8388_2 = {c5200};
    Full_Adder FA_8388(s8388, c8388, in8388_1, in8388_2, s1816[0]);
    wire[0:0] s8389, in8389_1, in8389_2;
    wire c8389;
    assign in8389_1 = {c5202};
    assign in8389_2 = {c5203};
    Full_Adder FA_8389(s8389, c8389, in8389_1, in8389_2, c5201);
    wire[0:0] s8390, in8390_1, in8390_2;
    wire c8390;
    assign in8390_1 = {c5205};
    assign in8390_2 = {c5206};
    Full_Adder FA_8390(s8390, c8390, in8390_1, in8390_2, c5204);
    wire[0:0] s8391, in8391_1, in8391_2;
    wire c8391;
    assign in8391_1 = {c5208};
    assign in8391_2 = {c5209};
    Full_Adder FA_8391(s8391, c8391, in8391_1, in8391_2, c5207);
    wire[0:0] s8392, in8392_1, in8392_2;
    wire c8392;
    assign in8392_1 = {c5211};
    assign in8392_2 = {c5212};
    Full_Adder FA_8392(s8392, c8392, in8392_1, in8392_2, c5210);
    wire[0:0] s8393, in8393_1, in8393_2;
    wire c8393;
    assign in8393_1 = {c5214};
    assign in8393_2 = {c5215};
    Full_Adder FA_8393(s8393, c8393, in8393_1, in8393_2, c5213);
    wire[0:0] s8394, in8394_1, in8394_2;
    wire c8394;
    assign in8394_1 = {c5217};
    assign in8394_2 = {s5218[0]};
    Full_Adder FA_8394(s8394, c8394, in8394_1, in8394_2, c5216);
    wire[0:0] s8395, in8395_1, in8395_2;
    wire c8395;
    assign in8395_1 = {s5220[0]};
    assign in8395_2 = {s5221[0]};
    Full_Adder FA_8395(s8395, c8395, in8395_1, in8395_2, s5219[0]);
    wire[0:0] s8396, in8396_1, in8396_2;
    wire c8396;
    assign in8396_1 = {s5223[0]};
    assign in8396_2 = {s5224[0]};
    Full_Adder FA_8396(s8396, c8396, in8396_1, in8396_2, s5222[0]);
    wire[0:0] s8397, in8397_1, in8397_2;
    wire c8397;
    assign in8397_1 = {s5226[0]};
    assign in8397_2 = {s5227[0]};
    Full_Adder FA_8397(s8397, c8397, in8397_1, in8397_2, s5225[0]);
    wire[0:0] s8398, in8398_1, in8398_2;
    wire c8398;
    assign in8398_1 = {s5229[0]};
    assign in8398_2 = {s5230[0]};
    Full_Adder FA_8398(s8398, c8398, in8398_1, in8398_2, s5228[0]);
    wire[0:0] s8399, in8399_1, in8399_2;
    wire c8399;
    assign in8399_1 = {s5232[0]};
    assign in8399_2 = {s5233[0]};
    Full_Adder FA_8399(s8399, c8399, in8399_1, in8399_2, s5231[0]);
    wire[0:0] s8400, in8400_1, in8400_2;
    wire c8400;
    assign in8400_1 = {s5235[0]};
    assign in8400_2 = {s5236[0]};
    Full_Adder FA_8400(s8400, c8400, in8400_1, in8400_2, s5234[0]);
    wire[0:0] s8401, in8401_1, in8401_2;
    wire c8401;
    assign in8401_1 = {c5218};
    assign in8401_2 = {c5219};
    Full_Adder FA_8401(s8401, c8401, in8401_1, in8401_2, s1821[0]);
    wire[0:0] s8402, in8402_1, in8402_2;
    wire c8402;
    assign in8402_1 = {c5221};
    assign in8402_2 = {c5222};
    Full_Adder FA_8402(s8402, c8402, in8402_1, in8402_2, c5220);
    wire[0:0] s8403, in8403_1, in8403_2;
    wire c8403;
    assign in8403_1 = {c5224};
    assign in8403_2 = {c5225};
    Full_Adder FA_8403(s8403, c8403, in8403_1, in8403_2, c5223);
    wire[0:0] s8404, in8404_1, in8404_2;
    wire c8404;
    assign in8404_1 = {c5227};
    assign in8404_2 = {c5228};
    Full_Adder FA_8404(s8404, c8404, in8404_1, in8404_2, c5226);
    wire[0:0] s8405, in8405_1, in8405_2;
    wire c8405;
    assign in8405_1 = {c5230};
    assign in8405_2 = {c5231};
    Full_Adder FA_8405(s8405, c8405, in8405_1, in8405_2, c5229);
    wire[0:0] s8406, in8406_1, in8406_2;
    wire c8406;
    assign in8406_1 = {c5233};
    assign in8406_2 = {c5234};
    Full_Adder FA_8406(s8406, c8406, in8406_1, in8406_2, c5232);
    wire[0:0] s8407, in8407_1, in8407_2;
    wire c8407;
    assign in8407_1 = {c5236};
    assign in8407_2 = {s5237[0]};
    Full_Adder FA_8407(s8407, c8407, in8407_1, in8407_2, c5235);
    wire[0:0] s8408, in8408_1, in8408_2;
    wire c8408;
    assign in8408_1 = {s5239[0]};
    assign in8408_2 = {s5240[0]};
    Full_Adder FA_8408(s8408, c8408, in8408_1, in8408_2, s5238[0]);
    wire[0:0] s8409, in8409_1, in8409_2;
    wire c8409;
    assign in8409_1 = {s5242[0]};
    assign in8409_2 = {s5243[0]};
    Full_Adder FA_8409(s8409, c8409, in8409_1, in8409_2, s5241[0]);
    wire[0:0] s8410, in8410_1, in8410_2;
    wire c8410;
    assign in8410_1 = {s5245[0]};
    assign in8410_2 = {s5246[0]};
    Full_Adder FA_8410(s8410, c8410, in8410_1, in8410_2, s5244[0]);
    wire[0:0] s8411, in8411_1, in8411_2;
    wire c8411;
    assign in8411_1 = {s5248[0]};
    assign in8411_2 = {s5249[0]};
    Full_Adder FA_8411(s8411, c8411, in8411_1, in8411_2, s5247[0]);
    wire[0:0] s8412, in8412_1, in8412_2;
    wire c8412;
    assign in8412_1 = {s5251[0]};
    assign in8412_2 = {s5252[0]};
    Full_Adder FA_8412(s8412, c8412, in8412_1, in8412_2, s5250[0]);
    wire[0:0] s8413, in8413_1, in8413_2;
    wire c8413;
    assign in8413_1 = {s5254[0]};
    assign in8413_2 = {s5255[0]};
    Full_Adder FA_8413(s8413, c8413, in8413_1, in8413_2, s5253[0]);
    wire[0:0] s8414, in8414_1, in8414_2;
    wire c8414;
    assign in8414_1 = {c5237};
    assign in8414_2 = {c5238};
    Full_Adder FA_8414(s8414, c8414, in8414_1, in8414_2, s1827[0]);
    wire[0:0] s8415, in8415_1, in8415_2;
    wire c8415;
    assign in8415_1 = {c5240};
    assign in8415_2 = {c5241};
    Full_Adder FA_8415(s8415, c8415, in8415_1, in8415_2, c5239);
    wire[0:0] s8416, in8416_1, in8416_2;
    wire c8416;
    assign in8416_1 = {c5243};
    assign in8416_2 = {c5244};
    Full_Adder FA_8416(s8416, c8416, in8416_1, in8416_2, c5242);
    wire[0:0] s8417, in8417_1, in8417_2;
    wire c8417;
    assign in8417_1 = {c5246};
    assign in8417_2 = {c5247};
    Full_Adder FA_8417(s8417, c8417, in8417_1, in8417_2, c5245);
    wire[0:0] s8418, in8418_1, in8418_2;
    wire c8418;
    assign in8418_1 = {c5249};
    assign in8418_2 = {c5250};
    Full_Adder FA_8418(s8418, c8418, in8418_1, in8418_2, c5248);
    wire[0:0] s8419, in8419_1, in8419_2;
    wire c8419;
    assign in8419_1 = {c5252};
    assign in8419_2 = {c5253};
    Full_Adder FA_8419(s8419, c8419, in8419_1, in8419_2, c5251);
    wire[0:0] s8420, in8420_1, in8420_2;
    wire c8420;
    assign in8420_1 = {c5255};
    assign in8420_2 = {s5256[0]};
    Full_Adder FA_8420(s8420, c8420, in8420_1, in8420_2, c5254);
    wire[0:0] s8421, in8421_1, in8421_2;
    wire c8421;
    assign in8421_1 = {s5258[0]};
    assign in8421_2 = {s5259[0]};
    Full_Adder FA_8421(s8421, c8421, in8421_1, in8421_2, s5257[0]);
    wire[0:0] s8422, in8422_1, in8422_2;
    wire c8422;
    assign in8422_1 = {s5261[0]};
    assign in8422_2 = {s5262[0]};
    Full_Adder FA_8422(s8422, c8422, in8422_1, in8422_2, s5260[0]);
    wire[0:0] s8423, in8423_1, in8423_2;
    wire c8423;
    assign in8423_1 = {s5264[0]};
    assign in8423_2 = {s5265[0]};
    Full_Adder FA_8423(s8423, c8423, in8423_1, in8423_2, s5263[0]);
    wire[0:0] s8424, in8424_1, in8424_2;
    wire c8424;
    assign in8424_1 = {s5267[0]};
    assign in8424_2 = {s5268[0]};
    Full_Adder FA_8424(s8424, c8424, in8424_1, in8424_2, s5266[0]);
    wire[0:0] s8425, in8425_1, in8425_2;
    wire c8425;
    assign in8425_1 = {s5270[0]};
    assign in8425_2 = {s5271[0]};
    Full_Adder FA_8425(s8425, c8425, in8425_1, in8425_2, s5269[0]);
    wire[0:0] s8426, in8426_1, in8426_2;
    wire c8426;
    assign in8426_1 = {s5273[0]};
    assign in8426_2 = {s5274[0]};
    Full_Adder FA_8426(s8426, c8426, in8426_1, in8426_2, s5272[0]);
    wire[0:0] s8427, in8427_1, in8427_2;
    wire c8427;
    assign in8427_1 = {c5256};
    assign in8427_2 = {c5257};
    Full_Adder FA_8427(s8427, c8427, in8427_1, in8427_2, s1834[0]);
    wire[0:0] s8428, in8428_1, in8428_2;
    wire c8428;
    assign in8428_1 = {c5259};
    assign in8428_2 = {c5260};
    Full_Adder FA_8428(s8428, c8428, in8428_1, in8428_2, c5258);
    wire[0:0] s8429, in8429_1, in8429_2;
    wire c8429;
    assign in8429_1 = {c5262};
    assign in8429_2 = {c5263};
    Full_Adder FA_8429(s8429, c8429, in8429_1, in8429_2, c5261);
    wire[0:0] s8430, in8430_1, in8430_2;
    wire c8430;
    assign in8430_1 = {c5265};
    assign in8430_2 = {c5266};
    Full_Adder FA_8430(s8430, c8430, in8430_1, in8430_2, c5264);
    wire[0:0] s8431, in8431_1, in8431_2;
    wire c8431;
    assign in8431_1 = {c5268};
    assign in8431_2 = {c5269};
    Full_Adder FA_8431(s8431, c8431, in8431_1, in8431_2, c5267);
    wire[0:0] s8432, in8432_1, in8432_2;
    wire c8432;
    assign in8432_1 = {c5271};
    assign in8432_2 = {c5272};
    Full_Adder FA_8432(s8432, c8432, in8432_1, in8432_2, c5270);
    wire[0:0] s8433, in8433_1, in8433_2;
    wire c8433;
    assign in8433_1 = {c5274};
    assign in8433_2 = {s5275[0]};
    Full_Adder FA_8433(s8433, c8433, in8433_1, in8433_2, c5273);
    wire[0:0] s8434, in8434_1, in8434_2;
    wire c8434;
    assign in8434_1 = {s5277[0]};
    assign in8434_2 = {s5278[0]};
    Full_Adder FA_8434(s8434, c8434, in8434_1, in8434_2, s5276[0]);
    wire[0:0] s8435, in8435_1, in8435_2;
    wire c8435;
    assign in8435_1 = {s5280[0]};
    assign in8435_2 = {s5281[0]};
    Full_Adder FA_8435(s8435, c8435, in8435_1, in8435_2, s5279[0]);
    wire[0:0] s8436, in8436_1, in8436_2;
    wire c8436;
    assign in8436_1 = {s5283[0]};
    assign in8436_2 = {s5284[0]};
    Full_Adder FA_8436(s8436, c8436, in8436_1, in8436_2, s5282[0]);
    wire[0:0] s8437, in8437_1, in8437_2;
    wire c8437;
    assign in8437_1 = {s5286[0]};
    assign in8437_2 = {s5287[0]};
    Full_Adder FA_8437(s8437, c8437, in8437_1, in8437_2, s5285[0]);
    wire[0:0] s8438, in8438_1, in8438_2;
    wire c8438;
    assign in8438_1 = {s5289[0]};
    assign in8438_2 = {s5290[0]};
    Full_Adder FA_8438(s8438, c8438, in8438_1, in8438_2, s5288[0]);
    wire[0:0] s8439, in8439_1, in8439_2;
    wire c8439;
    assign in8439_1 = {s5292[0]};
    assign in8439_2 = {s5293[0]};
    Full_Adder FA_8439(s8439, c8439, in8439_1, in8439_2, s5291[0]);
    wire[0:0] s8440, in8440_1, in8440_2;
    wire c8440;
    assign in8440_1 = {c5275};
    assign in8440_2 = {c5276};
    Full_Adder FA_8440(s8440, c8440, in8440_1, in8440_2, s1842[0]);
    wire[0:0] s8441, in8441_1, in8441_2;
    wire c8441;
    assign in8441_1 = {c5278};
    assign in8441_2 = {c5279};
    Full_Adder FA_8441(s8441, c8441, in8441_1, in8441_2, c5277);
    wire[0:0] s8442, in8442_1, in8442_2;
    wire c8442;
    assign in8442_1 = {c5281};
    assign in8442_2 = {c5282};
    Full_Adder FA_8442(s8442, c8442, in8442_1, in8442_2, c5280);
    wire[0:0] s8443, in8443_1, in8443_2;
    wire c8443;
    assign in8443_1 = {c5284};
    assign in8443_2 = {c5285};
    Full_Adder FA_8443(s8443, c8443, in8443_1, in8443_2, c5283);
    wire[0:0] s8444, in8444_1, in8444_2;
    wire c8444;
    assign in8444_1 = {c5287};
    assign in8444_2 = {c5288};
    Full_Adder FA_8444(s8444, c8444, in8444_1, in8444_2, c5286);
    wire[0:0] s8445, in8445_1, in8445_2;
    wire c8445;
    assign in8445_1 = {c5290};
    assign in8445_2 = {c5291};
    Full_Adder FA_8445(s8445, c8445, in8445_1, in8445_2, c5289);
    wire[0:0] s8446, in8446_1, in8446_2;
    wire c8446;
    assign in8446_1 = {c5293};
    assign in8446_2 = {s5294[0]};
    Full_Adder FA_8446(s8446, c8446, in8446_1, in8446_2, c5292);
    wire[0:0] s8447, in8447_1, in8447_2;
    wire c8447;
    assign in8447_1 = {s5296[0]};
    assign in8447_2 = {s5297[0]};
    Full_Adder FA_8447(s8447, c8447, in8447_1, in8447_2, s5295[0]);
    wire[0:0] s8448, in8448_1, in8448_2;
    wire c8448;
    assign in8448_1 = {s5299[0]};
    assign in8448_2 = {s5300[0]};
    Full_Adder FA_8448(s8448, c8448, in8448_1, in8448_2, s5298[0]);
    wire[0:0] s8449, in8449_1, in8449_2;
    wire c8449;
    assign in8449_1 = {s5302[0]};
    assign in8449_2 = {s5303[0]};
    Full_Adder FA_8449(s8449, c8449, in8449_1, in8449_2, s5301[0]);
    wire[0:0] s8450, in8450_1, in8450_2;
    wire c8450;
    assign in8450_1 = {s5305[0]};
    assign in8450_2 = {s5306[0]};
    Full_Adder FA_8450(s8450, c8450, in8450_1, in8450_2, s5304[0]);
    wire[0:0] s8451, in8451_1, in8451_2;
    wire c8451;
    assign in8451_1 = {s5308[0]};
    assign in8451_2 = {s5309[0]};
    Full_Adder FA_8451(s8451, c8451, in8451_1, in8451_2, s5307[0]);
    wire[0:0] s8452, in8452_1, in8452_2;
    wire c8452;
    assign in8452_1 = {s5311[0]};
    assign in8452_2 = {s5312[0]};
    Full_Adder FA_8452(s8452, c8452, in8452_1, in8452_2, s5310[0]);
    wire[0:0] s8453, in8453_1, in8453_2;
    wire c8453;
    assign in8453_1 = {c5294};
    assign in8453_2 = {c5295};
    Full_Adder FA_8453(s8453, c8453, in8453_1, in8453_2, s1851[0]);
    wire[0:0] s8454, in8454_1, in8454_2;
    wire c8454;
    assign in8454_1 = {c5297};
    assign in8454_2 = {c5298};
    Full_Adder FA_8454(s8454, c8454, in8454_1, in8454_2, c5296);
    wire[0:0] s8455, in8455_1, in8455_2;
    wire c8455;
    assign in8455_1 = {c5300};
    assign in8455_2 = {c5301};
    Full_Adder FA_8455(s8455, c8455, in8455_1, in8455_2, c5299);
    wire[0:0] s8456, in8456_1, in8456_2;
    wire c8456;
    assign in8456_1 = {c5303};
    assign in8456_2 = {c5304};
    Full_Adder FA_8456(s8456, c8456, in8456_1, in8456_2, c5302);
    wire[0:0] s8457, in8457_1, in8457_2;
    wire c8457;
    assign in8457_1 = {c5306};
    assign in8457_2 = {c5307};
    Full_Adder FA_8457(s8457, c8457, in8457_1, in8457_2, c5305);
    wire[0:0] s8458, in8458_1, in8458_2;
    wire c8458;
    assign in8458_1 = {c5309};
    assign in8458_2 = {c5310};
    Full_Adder FA_8458(s8458, c8458, in8458_1, in8458_2, c5308);
    wire[0:0] s8459, in8459_1, in8459_2;
    wire c8459;
    assign in8459_1 = {c5312};
    assign in8459_2 = {s5313[0]};
    Full_Adder FA_8459(s8459, c8459, in8459_1, in8459_2, c5311);
    wire[0:0] s8460, in8460_1, in8460_2;
    wire c8460;
    assign in8460_1 = {s5315[0]};
    assign in8460_2 = {s5316[0]};
    Full_Adder FA_8460(s8460, c8460, in8460_1, in8460_2, s5314[0]);
    wire[0:0] s8461, in8461_1, in8461_2;
    wire c8461;
    assign in8461_1 = {s5318[0]};
    assign in8461_2 = {s5319[0]};
    Full_Adder FA_8461(s8461, c8461, in8461_1, in8461_2, s5317[0]);
    wire[0:0] s8462, in8462_1, in8462_2;
    wire c8462;
    assign in8462_1 = {s5321[0]};
    assign in8462_2 = {s5322[0]};
    Full_Adder FA_8462(s8462, c8462, in8462_1, in8462_2, s5320[0]);
    wire[0:0] s8463, in8463_1, in8463_2;
    wire c8463;
    assign in8463_1 = {s5324[0]};
    assign in8463_2 = {s5325[0]};
    Full_Adder FA_8463(s8463, c8463, in8463_1, in8463_2, s5323[0]);
    wire[0:0] s8464, in8464_1, in8464_2;
    wire c8464;
    assign in8464_1 = {s5327[0]};
    assign in8464_2 = {s5328[0]};
    Full_Adder FA_8464(s8464, c8464, in8464_1, in8464_2, s5326[0]);
    wire[0:0] s8465, in8465_1, in8465_2;
    wire c8465;
    assign in8465_1 = {s5330[0]};
    assign in8465_2 = {s5331[0]};
    Full_Adder FA_8465(s8465, c8465, in8465_1, in8465_2, s5329[0]);
    wire[0:0] s8466, in8466_1, in8466_2;
    wire c8466;
    assign in8466_1 = {c5313};
    assign in8466_2 = {c5314};
    Full_Adder FA_8466(s8466, c8466, in8466_1, in8466_2, s1861[0]);
    wire[0:0] s8467, in8467_1, in8467_2;
    wire c8467;
    assign in8467_1 = {c5316};
    assign in8467_2 = {c5317};
    Full_Adder FA_8467(s8467, c8467, in8467_1, in8467_2, c5315);
    wire[0:0] s8468, in8468_1, in8468_2;
    wire c8468;
    assign in8468_1 = {c5319};
    assign in8468_2 = {c5320};
    Full_Adder FA_8468(s8468, c8468, in8468_1, in8468_2, c5318);
    wire[0:0] s8469, in8469_1, in8469_2;
    wire c8469;
    assign in8469_1 = {c5322};
    assign in8469_2 = {c5323};
    Full_Adder FA_8469(s8469, c8469, in8469_1, in8469_2, c5321);
    wire[0:0] s8470, in8470_1, in8470_2;
    wire c8470;
    assign in8470_1 = {c5325};
    assign in8470_2 = {c5326};
    Full_Adder FA_8470(s8470, c8470, in8470_1, in8470_2, c5324);
    wire[0:0] s8471, in8471_1, in8471_2;
    wire c8471;
    assign in8471_1 = {c5328};
    assign in8471_2 = {c5329};
    Full_Adder FA_8471(s8471, c8471, in8471_1, in8471_2, c5327);
    wire[0:0] s8472, in8472_1, in8472_2;
    wire c8472;
    assign in8472_1 = {c5331};
    assign in8472_2 = {s5332[0]};
    Full_Adder FA_8472(s8472, c8472, in8472_1, in8472_2, c5330);
    wire[0:0] s8473, in8473_1, in8473_2;
    wire c8473;
    assign in8473_1 = {s5334[0]};
    assign in8473_2 = {s5335[0]};
    Full_Adder FA_8473(s8473, c8473, in8473_1, in8473_2, s5333[0]);
    wire[0:0] s8474, in8474_1, in8474_2;
    wire c8474;
    assign in8474_1 = {s5337[0]};
    assign in8474_2 = {s5338[0]};
    Full_Adder FA_8474(s8474, c8474, in8474_1, in8474_2, s5336[0]);
    wire[0:0] s8475, in8475_1, in8475_2;
    wire c8475;
    assign in8475_1 = {s5340[0]};
    assign in8475_2 = {s5341[0]};
    Full_Adder FA_8475(s8475, c8475, in8475_1, in8475_2, s5339[0]);
    wire[0:0] s8476, in8476_1, in8476_2;
    wire c8476;
    assign in8476_1 = {s5343[0]};
    assign in8476_2 = {s5344[0]};
    Full_Adder FA_8476(s8476, c8476, in8476_1, in8476_2, s5342[0]);
    wire[0:0] s8477, in8477_1, in8477_2;
    wire c8477;
    assign in8477_1 = {s5346[0]};
    assign in8477_2 = {s5347[0]};
    Full_Adder FA_8477(s8477, c8477, in8477_1, in8477_2, s5345[0]);
    wire[0:0] s8478, in8478_1, in8478_2;
    wire c8478;
    assign in8478_1 = {s5349[0]};
    assign in8478_2 = {s5350[0]};
    Full_Adder FA_8478(s8478, c8478, in8478_1, in8478_2, s5348[0]);
    wire[0:0] s8479, in8479_1, in8479_2;
    wire c8479;
    assign in8479_1 = {c5332};
    assign in8479_2 = {c5333};
    Full_Adder FA_8479(s8479, c8479, in8479_1, in8479_2, s1872[0]);
    wire[0:0] s8480, in8480_1, in8480_2;
    wire c8480;
    assign in8480_1 = {c5335};
    assign in8480_2 = {c5336};
    Full_Adder FA_8480(s8480, c8480, in8480_1, in8480_2, c5334);
    wire[0:0] s8481, in8481_1, in8481_2;
    wire c8481;
    assign in8481_1 = {c5338};
    assign in8481_2 = {c5339};
    Full_Adder FA_8481(s8481, c8481, in8481_1, in8481_2, c5337);
    wire[0:0] s8482, in8482_1, in8482_2;
    wire c8482;
    assign in8482_1 = {c5341};
    assign in8482_2 = {c5342};
    Full_Adder FA_8482(s8482, c8482, in8482_1, in8482_2, c5340);
    wire[0:0] s8483, in8483_1, in8483_2;
    wire c8483;
    assign in8483_1 = {c5344};
    assign in8483_2 = {c5345};
    Full_Adder FA_8483(s8483, c8483, in8483_1, in8483_2, c5343);
    wire[0:0] s8484, in8484_1, in8484_2;
    wire c8484;
    assign in8484_1 = {c5347};
    assign in8484_2 = {c5348};
    Full_Adder FA_8484(s8484, c8484, in8484_1, in8484_2, c5346);
    wire[0:0] s8485, in8485_1, in8485_2;
    wire c8485;
    assign in8485_1 = {c5350};
    assign in8485_2 = {s5351[0]};
    Full_Adder FA_8485(s8485, c8485, in8485_1, in8485_2, c5349);
    wire[0:0] s8486, in8486_1, in8486_2;
    wire c8486;
    assign in8486_1 = {s5353[0]};
    assign in8486_2 = {s5354[0]};
    Full_Adder FA_8486(s8486, c8486, in8486_1, in8486_2, s5352[0]);
    wire[0:0] s8487, in8487_1, in8487_2;
    wire c8487;
    assign in8487_1 = {s5356[0]};
    assign in8487_2 = {s5357[0]};
    Full_Adder FA_8487(s8487, c8487, in8487_1, in8487_2, s5355[0]);
    wire[0:0] s8488, in8488_1, in8488_2;
    wire c8488;
    assign in8488_1 = {s5359[0]};
    assign in8488_2 = {s5360[0]};
    Full_Adder FA_8488(s8488, c8488, in8488_1, in8488_2, s5358[0]);
    wire[0:0] s8489, in8489_1, in8489_2;
    wire c8489;
    assign in8489_1 = {s5362[0]};
    assign in8489_2 = {s5363[0]};
    Full_Adder FA_8489(s8489, c8489, in8489_1, in8489_2, s5361[0]);
    wire[0:0] s8490, in8490_1, in8490_2;
    wire c8490;
    assign in8490_1 = {s5365[0]};
    assign in8490_2 = {s5366[0]};
    Full_Adder FA_8490(s8490, c8490, in8490_1, in8490_2, s5364[0]);
    wire[0:0] s8491, in8491_1, in8491_2;
    wire c8491;
    assign in8491_1 = {s5368[0]};
    assign in8491_2 = {s5369[0]};
    Full_Adder FA_8491(s8491, c8491, in8491_1, in8491_2, s5367[0]);
    wire[0:0] s8492, in8492_1, in8492_2;
    wire c8492;
    assign in8492_1 = {c5351};
    assign in8492_2 = {c5352};
    Full_Adder FA_8492(s8492, c8492, in8492_1, in8492_2, s1884[0]);
    wire[0:0] s8493, in8493_1, in8493_2;
    wire c8493;
    assign in8493_1 = {c5354};
    assign in8493_2 = {c5355};
    Full_Adder FA_8493(s8493, c8493, in8493_1, in8493_2, c5353);
    wire[0:0] s8494, in8494_1, in8494_2;
    wire c8494;
    assign in8494_1 = {c5357};
    assign in8494_2 = {c5358};
    Full_Adder FA_8494(s8494, c8494, in8494_1, in8494_2, c5356);
    wire[0:0] s8495, in8495_1, in8495_2;
    wire c8495;
    assign in8495_1 = {c5360};
    assign in8495_2 = {c5361};
    Full_Adder FA_8495(s8495, c8495, in8495_1, in8495_2, c5359);
    wire[0:0] s8496, in8496_1, in8496_2;
    wire c8496;
    assign in8496_1 = {c5363};
    assign in8496_2 = {c5364};
    Full_Adder FA_8496(s8496, c8496, in8496_1, in8496_2, c5362);
    wire[0:0] s8497, in8497_1, in8497_2;
    wire c8497;
    assign in8497_1 = {c5366};
    assign in8497_2 = {c5367};
    Full_Adder FA_8497(s8497, c8497, in8497_1, in8497_2, c5365);
    wire[0:0] s8498, in8498_1, in8498_2;
    wire c8498;
    assign in8498_1 = {c5369};
    assign in8498_2 = {s5370[0]};
    Full_Adder FA_8498(s8498, c8498, in8498_1, in8498_2, c5368);
    wire[0:0] s8499, in8499_1, in8499_2;
    wire c8499;
    assign in8499_1 = {s5372[0]};
    assign in8499_2 = {s5373[0]};
    Full_Adder FA_8499(s8499, c8499, in8499_1, in8499_2, s5371[0]);
    wire[0:0] s8500, in8500_1, in8500_2;
    wire c8500;
    assign in8500_1 = {s5375[0]};
    assign in8500_2 = {s5376[0]};
    Full_Adder FA_8500(s8500, c8500, in8500_1, in8500_2, s5374[0]);
    wire[0:0] s8501, in8501_1, in8501_2;
    wire c8501;
    assign in8501_1 = {s5378[0]};
    assign in8501_2 = {s5379[0]};
    Full_Adder FA_8501(s8501, c8501, in8501_1, in8501_2, s5377[0]);
    wire[0:0] s8502, in8502_1, in8502_2;
    wire c8502;
    assign in8502_1 = {s5381[0]};
    assign in8502_2 = {s5382[0]};
    Full_Adder FA_8502(s8502, c8502, in8502_1, in8502_2, s5380[0]);
    wire[0:0] s8503, in8503_1, in8503_2;
    wire c8503;
    assign in8503_1 = {s5384[0]};
    assign in8503_2 = {s5385[0]};
    Full_Adder FA_8503(s8503, c8503, in8503_1, in8503_2, s5383[0]);
    wire[0:0] s8504, in8504_1, in8504_2;
    wire c8504;
    assign in8504_1 = {s5387[0]};
    assign in8504_2 = {s5388[0]};
    Full_Adder FA_8504(s8504, c8504, in8504_1, in8504_2, s5386[0]);
    wire[0:0] s8505, in8505_1, in8505_2;
    wire c8505;
    assign in8505_1 = {c5370};
    assign in8505_2 = {c5371};
    Full_Adder FA_8505(s8505, c8505, in8505_1, in8505_2, s1897[0]);
    wire[0:0] s8506, in8506_1, in8506_2;
    wire c8506;
    assign in8506_1 = {c5373};
    assign in8506_2 = {c5374};
    Full_Adder FA_8506(s8506, c8506, in8506_1, in8506_2, c5372);
    wire[0:0] s8507, in8507_1, in8507_2;
    wire c8507;
    assign in8507_1 = {c5376};
    assign in8507_2 = {c5377};
    Full_Adder FA_8507(s8507, c8507, in8507_1, in8507_2, c5375);
    wire[0:0] s8508, in8508_1, in8508_2;
    wire c8508;
    assign in8508_1 = {c5379};
    assign in8508_2 = {c5380};
    Full_Adder FA_8508(s8508, c8508, in8508_1, in8508_2, c5378);
    wire[0:0] s8509, in8509_1, in8509_2;
    wire c8509;
    assign in8509_1 = {c5382};
    assign in8509_2 = {c5383};
    Full_Adder FA_8509(s8509, c8509, in8509_1, in8509_2, c5381);
    wire[0:0] s8510, in8510_1, in8510_2;
    wire c8510;
    assign in8510_1 = {c5385};
    assign in8510_2 = {c5386};
    Full_Adder FA_8510(s8510, c8510, in8510_1, in8510_2, c5384);
    wire[0:0] s8511, in8511_1, in8511_2;
    wire c8511;
    assign in8511_1 = {c5388};
    assign in8511_2 = {s5389[0]};
    Full_Adder FA_8511(s8511, c8511, in8511_1, in8511_2, c5387);
    wire[0:0] s8512, in8512_1, in8512_2;
    wire c8512;
    assign in8512_1 = {s5391[0]};
    assign in8512_2 = {s5392[0]};
    Full_Adder FA_8512(s8512, c8512, in8512_1, in8512_2, s5390[0]);
    wire[0:0] s8513, in8513_1, in8513_2;
    wire c8513;
    assign in8513_1 = {s5394[0]};
    assign in8513_2 = {s5395[0]};
    Full_Adder FA_8513(s8513, c8513, in8513_1, in8513_2, s5393[0]);
    wire[0:0] s8514, in8514_1, in8514_2;
    wire c8514;
    assign in8514_1 = {s5397[0]};
    assign in8514_2 = {s5398[0]};
    Full_Adder FA_8514(s8514, c8514, in8514_1, in8514_2, s5396[0]);
    wire[0:0] s8515, in8515_1, in8515_2;
    wire c8515;
    assign in8515_1 = {s5400[0]};
    assign in8515_2 = {s5401[0]};
    Full_Adder FA_8515(s8515, c8515, in8515_1, in8515_2, s5399[0]);
    wire[0:0] s8516, in8516_1, in8516_2;
    wire c8516;
    assign in8516_1 = {s5403[0]};
    assign in8516_2 = {s5404[0]};
    Full_Adder FA_8516(s8516, c8516, in8516_1, in8516_2, s5402[0]);
    wire[0:0] s8517, in8517_1, in8517_2;
    wire c8517;
    assign in8517_1 = {s5406[0]};
    assign in8517_2 = {s5407[0]};
    Full_Adder FA_8517(s8517, c8517, in8517_1, in8517_2, s5405[0]);
    wire[0:0] s8518, in8518_1, in8518_2;
    wire c8518;
    assign in8518_1 = {c5389};
    assign in8518_2 = {c5390};
    Full_Adder FA_8518(s8518, c8518, in8518_1, in8518_2, s1911[0]);
    wire[0:0] s8519, in8519_1, in8519_2;
    wire c8519;
    assign in8519_1 = {c5392};
    assign in8519_2 = {c5393};
    Full_Adder FA_8519(s8519, c8519, in8519_1, in8519_2, c5391);
    wire[0:0] s8520, in8520_1, in8520_2;
    wire c8520;
    assign in8520_1 = {c5395};
    assign in8520_2 = {c5396};
    Full_Adder FA_8520(s8520, c8520, in8520_1, in8520_2, c5394);
    wire[0:0] s8521, in8521_1, in8521_2;
    wire c8521;
    assign in8521_1 = {c5398};
    assign in8521_2 = {c5399};
    Full_Adder FA_8521(s8521, c8521, in8521_1, in8521_2, c5397);
    wire[0:0] s8522, in8522_1, in8522_2;
    wire c8522;
    assign in8522_1 = {c5401};
    assign in8522_2 = {c5402};
    Full_Adder FA_8522(s8522, c8522, in8522_1, in8522_2, c5400);
    wire[0:0] s8523, in8523_1, in8523_2;
    wire c8523;
    assign in8523_1 = {c5404};
    assign in8523_2 = {c5405};
    Full_Adder FA_8523(s8523, c8523, in8523_1, in8523_2, c5403);
    wire[0:0] s8524, in8524_1, in8524_2;
    wire c8524;
    assign in8524_1 = {c5407};
    assign in8524_2 = {s5408[0]};
    Full_Adder FA_8524(s8524, c8524, in8524_1, in8524_2, c5406);
    wire[0:0] s8525, in8525_1, in8525_2;
    wire c8525;
    assign in8525_1 = {s5410[0]};
    assign in8525_2 = {s5411[0]};
    Full_Adder FA_8525(s8525, c8525, in8525_1, in8525_2, s5409[0]);
    wire[0:0] s8526, in8526_1, in8526_2;
    wire c8526;
    assign in8526_1 = {s5413[0]};
    assign in8526_2 = {s5414[0]};
    Full_Adder FA_8526(s8526, c8526, in8526_1, in8526_2, s5412[0]);
    wire[0:0] s8527, in8527_1, in8527_2;
    wire c8527;
    assign in8527_1 = {s5416[0]};
    assign in8527_2 = {s5417[0]};
    Full_Adder FA_8527(s8527, c8527, in8527_1, in8527_2, s5415[0]);
    wire[0:0] s8528, in8528_1, in8528_2;
    wire c8528;
    assign in8528_1 = {s5419[0]};
    assign in8528_2 = {s5420[0]};
    Full_Adder FA_8528(s8528, c8528, in8528_1, in8528_2, s5418[0]);
    wire[0:0] s8529, in8529_1, in8529_2;
    wire c8529;
    assign in8529_1 = {s5422[0]};
    assign in8529_2 = {s5423[0]};
    Full_Adder FA_8529(s8529, c8529, in8529_1, in8529_2, s5421[0]);
    wire[0:0] s8530, in8530_1, in8530_2;
    wire c8530;
    assign in8530_1 = {s5425[0]};
    assign in8530_2 = {s5426[0]};
    Full_Adder FA_8530(s8530, c8530, in8530_1, in8530_2, s5424[0]);
    wire[0:0] s8531, in8531_1, in8531_2;
    wire c8531;
    assign in8531_1 = {c5408};
    assign in8531_2 = {c5409};
    Full_Adder FA_8531(s8531, c8531, in8531_1, in8531_2, s1926[0]);
    wire[0:0] s8532, in8532_1, in8532_2;
    wire c8532;
    assign in8532_1 = {c5411};
    assign in8532_2 = {c5412};
    Full_Adder FA_8532(s8532, c8532, in8532_1, in8532_2, c5410);
    wire[0:0] s8533, in8533_1, in8533_2;
    wire c8533;
    assign in8533_1 = {c5414};
    assign in8533_2 = {c5415};
    Full_Adder FA_8533(s8533, c8533, in8533_1, in8533_2, c5413);
    wire[0:0] s8534, in8534_1, in8534_2;
    wire c8534;
    assign in8534_1 = {c5417};
    assign in8534_2 = {c5418};
    Full_Adder FA_8534(s8534, c8534, in8534_1, in8534_2, c5416);
    wire[0:0] s8535, in8535_1, in8535_2;
    wire c8535;
    assign in8535_1 = {c5420};
    assign in8535_2 = {c5421};
    Full_Adder FA_8535(s8535, c8535, in8535_1, in8535_2, c5419);
    wire[0:0] s8536, in8536_1, in8536_2;
    wire c8536;
    assign in8536_1 = {c5423};
    assign in8536_2 = {c5424};
    Full_Adder FA_8536(s8536, c8536, in8536_1, in8536_2, c5422);
    wire[0:0] s8537, in8537_1, in8537_2;
    wire c8537;
    assign in8537_1 = {c5426};
    assign in8537_2 = {s5427[0]};
    Full_Adder FA_8537(s8537, c8537, in8537_1, in8537_2, c5425);
    wire[0:0] s8538, in8538_1, in8538_2;
    wire c8538;
    assign in8538_1 = {s5429[0]};
    assign in8538_2 = {s5430[0]};
    Full_Adder FA_8538(s8538, c8538, in8538_1, in8538_2, s5428[0]);
    wire[0:0] s8539, in8539_1, in8539_2;
    wire c8539;
    assign in8539_1 = {s5432[0]};
    assign in8539_2 = {s5433[0]};
    Full_Adder FA_8539(s8539, c8539, in8539_1, in8539_2, s5431[0]);
    wire[0:0] s8540, in8540_1, in8540_2;
    wire c8540;
    assign in8540_1 = {s5435[0]};
    assign in8540_2 = {s5436[0]};
    Full_Adder FA_8540(s8540, c8540, in8540_1, in8540_2, s5434[0]);
    wire[0:0] s8541, in8541_1, in8541_2;
    wire c8541;
    assign in8541_1 = {s5438[0]};
    assign in8541_2 = {s5439[0]};
    Full_Adder FA_8541(s8541, c8541, in8541_1, in8541_2, s5437[0]);
    wire[0:0] s8542, in8542_1, in8542_2;
    wire c8542;
    assign in8542_1 = {s5441[0]};
    assign in8542_2 = {s5442[0]};
    Full_Adder FA_8542(s8542, c8542, in8542_1, in8542_2, s5440[0]);
    wire[0:0] s8543, in8543_1, in8543_2;
    wire c8543;
    assign in8543_1 = {s5444[0]};
    assign in8543_2 = {s5445[0]};
    Full_Adder FA_8543(s8543, c8543, in8543_1, in8543_2, s5443[0]);
    wire[0:0] s8544, in8544_1, in8544_2;
    wire c8544;
    assign in8544_1 = {c5427};
    assign in8544_2 = {c5428};
    Full_Adder FA_8544(s8544, c8544, in8544_1, in8544_2, s1942[0]);
    wire[0:0] s8545, in8545_1, in8545_2;
    wire c8545;
    assign in8545_1 = {c5430};
    assign in8545_2 = {c5431};
    Full_Adder FA_8545(s8545, c8545, in8545_1, in8545_2, c5429);
    wire[0:0] s8546, in8546_1, in8546_2;
    wire c8546;
    assign in8546_1 = {c5433};
    assign in8546_2 = {c5434};
    Full_Adder FA_8546(s8546, c8546, in8546_1, in8546_2, c5432);
    wire[0:0] s8547, in8547_1, in8547_2;
    wire c8547;
    assign in8547_1 = {c5436};
    assign in8547_2 = {c5437};
    Full_Adder FA_8547(s8547, c8547, in8547_1, in8547_2, c5435);
    wire[0:0] s8548, in8548_1, in8548_2;
    wire c8548;
    assign in8548_1 = {c5439};
    assign in8548_2 = {c5440};
    Full_Adder FA_8548(s8548, c8548, in8548_1, in8548_2, c5438);
    wire[0:0] s8549, in8549_1, in8549_2;
    wire c8549;
    assign in8549_1 = {c5442};
    assign in8549_2 = {c5443};
    Full_Adder FA_8549(s8549, c8549, in8549_1, in8549_2, c5441);
    wire[0:0] s8550, in8550_1, in8550_2;
    wire c8550;
    assign in8550_1 = {c5445};
    assign in8550_2 = {s5446[0]};
    Full_Adder FA_8550(s8550, c8550, in8550_1, in8550_2, c5444);
    wire[0:0] s8551, in8551_1, in8551_2;
    wire c8551;
    assign in8551_1 = {s5448[0]};
    assign in8551_2 = {s5449[0]};
    Full_Adder FA_8551(s8551, c8551, in8551_1, in8551_2, s5447[0]);
    wire[0:0] s8552, in8552_1, in8552_2;
    wire c8552;
    assign in8552_1 = {s5451[0]};
    assign in8552_2 = {s5452[0]};
    Full_Adder FA_8552(s8552, c8552, in8552_1, in8552_2, s5450[0]);
    wire[0:0] s8553, in8553_1, in8553_2;
    wire c8553;
    assign in8553_1 = {s5454[0]};
    assign in8553_2 = {s5455[0]};
    Full_Adder FA_8553(s8553, c8553, in8553_1, in8553_2, s5453[0]);
    wire[0:0] s8554, in8554_1, in8554_2;
    wire c8554;
    assign in8554_1 = {s5457[0]};
    assign in8554_2 = {s5458[0]};
    Full_Adder FA_8554(s8554, c8554, in8554_1, in8554_2, s5456[0]);
    wire[0:0] s8555, in8555_1, in8555_2;
    wire c8555;
    assign in8555_1 = {s5460[0]};
    assign in8555_2 = {s5461[0]};
    Full_Adder FA_8555(s8555, c8555, in8555_1, in8555_2, s5459[0]);
    wire[0:0] s8556, in8556_1, in8556_2;
    wire c8556;
    assign in8556_1 = {s5463[0]};
    assign in8556_2 = {s5464[0]};
    Full_Adder FA_8556(s8556, c8556, in8556_1, in8556_2, s5462[0]);
    wire[0:0] s8557, in8557_1, in8557_2;
    wire c8557;
    assign in8557_1 = {c5446};
    assign in8557_2 = {c5447};
    Full_Adder FA_8557(s8557, c8557, in8557_1, in8557_2, s1959[0]);
    wire[0:0] s8558, in8558_1, in8558_2;
    wire c8558;
    assign in8558_1 = {c5449};
    assign in8558_2 = {c5450};
    Full_Adder FA_8558(s8558, c8558, in8558_1, in8558_2, c5448);
    wire[0:0] s8559, in8559_1, in8559_2;
    wire c8559;
    assign in8559_1 = {c5452};
    assign in8559_2 = {c5453};
    Full_Adder FA_8559(s8559, c8559, in8559_1, in8559_2, c5451);
    wire[0:0] s8560, in8560_1, in8560_2;
    wire c8560;
    assign in8560_1 = {c5455};
    assign in8560_2 = {c5456};
    Full_Adder FA_8560(s8560, c8560, in8560_1, in8560_2, c5454);
    wire[0:0] s8561, in8561_1, in8561_2;
    wire c8561;
    assign in8561_1 = {c5458};
    assign in8561_2 = {c5459};
    Full_Adder FA_8561(s8561, c8561, in8561_1, in8561_2, c5457);
    wire[0:0] s8562, in8562_1, in8562_2;
    wire c8562;
    assign in8562_1 = {c5461};
    assign in8562_2 = {c5462};
    Full_Adder FA_8562(s8562, c8562, in8562_1, in8562_2, c5460);
    wire[0:0] s8563, in8563_1, in8563_2;
    wire c8563;
    assign in8563_1 = {c5464};
    assign in8563_2 = {s5465[0]};
    Full_Adder FA_8563(s8563, c8563, in8563_1, in8563_2, c5463);
    wire[0:0] s8564, in8564_1, in8564_2;
    wire c8564;
    assign in8564_1 = {s5467[0]};
    assign in8564_2 = {s5468[0]};
    Full_Adder FA_8564(s8564, c8564, in8564_1, in8564_2, s5466[0]);
    wire[0:0] s8565, in8565_1, in8565_2;
    wire c8565;
    assign in8565_1 = {s5470[0]};
    assign in8565_2 = {s5471[0]};
    Full_Adder FA_8565(s8565, c8565, in8565_1, in8565_2, s5469[0]);
    wire[0:0] s8566, in8566_1, in8566_2;
    wire c8566;
    assign in8566_1 = {s5473[0]};
    assign in8566_2 = {s5474[0]};
    Full_Adder FA_8566(s8566, c8566, in8566_1, in8566_2, s5472[0]);
    wire[0:0] s8567, in8567_1, in8567_2;
    wire c8567;
    assign in8567_1 = {s5476[0]};
    assign in8567_2 = {s5477[0]};
    Full_Adder FA_8567(s8567, c8567, in8567_1, in8567_2, s5475[0]);
    wire[0:0] s8568, in8568_1, in8568_2;
    wire c8568;
    assign in8568_1 = {s5479[0]};
    assign in8568_2 = {s5480[0]};
    Full_Adder FA_8568(s8568, c8568, in8568_1, in8568_2, s5478[0]);
    wire[0:0] s8569, in8569_1, in8569_2;
    wire c8569;
    assign in8569_1 = {s5482[0]};
    assign in8569_2 = {s5483[0]};
    Full_Adder FA_8569(s8569, c8569, in8569_1, in8569_2, s5481[0]);
    wire[0:0] s8570, in8570_1, in8570_2;
    wire c8570;
    assign in8570_1 = {c5465};
    assign in8570_2 = {c5466};
    Full_Adder FA_8570(s8570, c8570, in8570_1, in8570_2, s1977[0]);
    wire[0:0] s8571, in8571_1, in8571_2;
    wire c8571;
    assign in8571_1 = {c5468};
    assign in8571_2 = {c5469};
    Full_Adder FA_8571(s8571, c8571, in8571_1, in8571_2, c5467);
    wire[0:0] s8572, in8572_1, in8572_2;
    wire c8572;
    assign in8572_1 = {c5471};
    assign in8572_2 = {c5472};
    Full_Adder FA_8572(s8572, c8572, in8572_1, in8572_2, c5470);
    wire[0:0] s8573, in8573_1, in8573_2;
    wire c8573;
    assign in8573_1 = {c5474};
    assign in8573_2 = {c5475};
    Full_Adder FA_8573(s8573, c8573, in8573_1, in8573_2, c5473);
    wire[0:0] s8574, in8574_1, in8574_2;
    wire c8574;
    assign in8574_1 = {c5477};
    assign in8574_2 = {c5478};
    Full_Adder FA_8574(s8574, c8574, in8574_1, in8574_2, c5476);
    wire[0:0] s8575, in8575_1, in8575_2;
    wire c8575;
    assign in8575_1 = {c5480};
    assign in8575_2 = {c5481};
    Full_Adder FA_8575(s8575, c8575, in8575_1, in8575_2, c5479);
    wire[0:0] s8576, in8576_1, in8576_2;
    wire c8576;
    assign in8576_1 = {c5483};
    assign in8576_2 = {s5484[0]};
    Full_Adder FA_8576(s8576, c8576, in8576_1, in8576_2, c5482);
    wire[0:0] s8577, in8577_1, in8577_2;
    wire c8577;
    assign in8577_1 = {s5486[0]};
    assign in8577_2 = {s5487[0]};
    Full_Adder FA_8577(s8577, c8577, in8577_1, in8577_2, s5485[0]);
    wire[0:0] s8578, in8578_1, in8578_2;
    wire c8578;
    assign in8578_1 = {s5489[0]};
    assign in8578_2 = {s5490[0]};
    Full_Adder FA_8578(s8578, c8578, in8578_1, in8578_2, s5488[0]);
    wire[0:0] s8579, in8579_1, in8579_2;
    wire c8579;
    assign in8579_1 = {s5492[0]};
    assign in8579_2 = {s5493[0]};
    Full_Adder FA_8579(s8579, c8579, in8579_1, in8579_2, s5491[0]);
    wire[0:0] s8580, in8580_1, in8580_2;
    wire c8580;
    assign in8580_1 = {s5495[0]};
    assign in8580_2 = {s5496[0]};
    Full_Adder FA_8580(s8580, c8580, in8580_1, in8580_2, s5494[0]);
    wire[0:0] s8581, in8581_1, in8581_2;
    wire c8581;
    assign in8581_1 = {s5498[0]};
    assign in8581_2 = {s5499[0]};
    Full_Adder FA_8581(s8581, c8581, in8581_1, in8581_2, s5497[0]);
    wire[0:0] s8582, in8582_1, in8582_2;
    wire c8582;
    assign in8582_1 = {s5501[0]};
    assign in8582_2 = {s5502[0]};
    Full_Adder FA_8582(s8582, c8582, in8582_1, in8582_2, s5500[0]);
    wire[0:0] s8583, in8583_1, in8583_2;
    wire c8583;
    assign in8583_1 = {c5484};
    assign in8583_2 = {c5485};
    Full_Adder FA_8583(s8583, c8583, in8583_1, in8583_2, s1996[0]);
    wire[0:0] s8584, in8584_1, in8584_2;
    wire c8584;
    assign in8584_1 = {c5487};
    assign in8584_2 = {c5488};
    Full_Adder FA_8584(s8584, c8584, in8584_1, in8584_2, c5486);
    wire[0:0] s8585, in8585_1, in8585_2;
    wire c8585;
    assign in8585_1 = {c5490};
    assign in8585_2 = {c5491};
    Full_Adder FA_8585(s8585, c8585, in8585_1, in8585_2, c5489);
    wire[0:0] s8586, in8586_1, in8586_2;
    wire c8586;
    assign in8586_1 = {c5493};
    assign in8586_2 = {c5494};
    Full_Adder FA_8586(s8586, c8586, in8586_1, in8586_2, c5492);
    wire[0:0] s8587, in8587_1, in8587_2;
    wire c8587;
    assign in8587_1 = {c5496};
    assign in8587_2 = {c5497};
    Full_Adder FA_8587(s8587, c8587, in8587_1, in8587_2, c5495);
    wire[0:0] s8588, in8588_1, in8588_2;
    wire c8588;
    assign in8588_1 = {c5499};
    assign in8588_2 = {c5500};
    Full_Adder FA_8588(s8588, c8588, in8588_1, in8588_2, c5498);
    wire[0:0] s8589, in8589_1, in8589_2;
    wire c8589;
    assign in8589_1 = {c5502};
    assign in8589_2 = {s5503[0]};
    Full_Adder FA_8589(s8589, c8589, in8589_1, in8589_2, c5501);
    wire[0:0] s8590, in8590_1, in8590_2;
    wire c8590;
    assign in8590_1 = {s5505[0]};
    assign in8590_2 = {s5506[0]};
    Full_Adder FA_8590(s8590, c8590, in8590_1, in8590_2, s5504[0]);
    wire[0:0] s8591, in8591_1, in8591_2;
    wire c8591;
    assign in8591_1 = {s5508[0]};
    assign in8591_2 = {s5509[0]};
    Full_Adder FA_8591(s8591, c8591, in8591_1, in8591_2, s5507[0]);
    wire[0:0] s8592, in8592_1, in8592_2;
    wire c8592;
    assign in8592_1 = {s5511[0]};
    assign in8592_2 = {s5512[0]};
    Full_Adder FA_8592(s8592, c8592, in8592_1, in8592_2, s5510[0]);
    wire[0:0] s8593, in8593_1, in8593_2;
    wire c8593;
    assign in8593_1 = {s5514[0]};
    assign in8593_2 = {s5515[0]};
    Full_Adder FA_8593(s8593, c8593, in8593_1, in8593_2, s5513[0]);
    wire[0:0] s8594, in8594_1, in8594_2;
    wire c8594;
    assign in8594_1 = {s5517[0]};
    assign in8594_2 = {s5518[0]};
    Full_Adder FA_8594(s8594, c8594, in8594_1, in8594_2, s5516[0]);
    wire[0:0] s8595, in8595_1, in8595_2;
    wire c8595;
    assign in8595_1 = {s5520[0]};
    assign in8595_2 = {s5521[0]};
    Full_Adder FA_8595(s8595, c8595, in8595_1, in8595_2, s5519[0]);
    wire[0:0] s8596, in8596_1, in8596_2;
    wire c8596;
    assign in8596_1 = {c5503};
    assign in8596_2 = {c5504};
    Full_Adder FA_8596(s8596, c8596, in8596_1, in8596_2, s2016[0]);
    wire[0:0] s8597, in8597_1, in8597_2;
    wire c8597;
    assign in8597_1 = {c5506};
    assign in8597_2 = {c5507};
    Full_Adder FA_8597(s8597, c8597, in8597_1, in8597_2, c5505);
    wire[0:0] s8598, in8598_1, in8598_2;
    wire c8598;
    assign in8598_1 = {c5509};
    assign in8598_2 = {c5510};
    Full_Adder FA_8598(s8598, c8598, in8598_1, in8598_2, c5508);
    wire[0:0] s8599, in8599_1, in8599_2;
    wire c8599;
    assign in8599_1 = {c5512};
    assign in8599_2 = {c5513};
    Full_Adder FA_8599(s8599, c8599, in8599_1, in8599_2, c5511);
    wire[0:0] s8600, in8600_1, in8600_2;
    wire c8600;
    assign in8600_1 = {c5515};
    assign in8600_2 = {c5516};
    Full_Adder FA_8600(s8600, c8600, in8600_1, in8600_2, c5514);
    wire[0:0] s8601, in8601_1, in8601_2;
    wire c8601;
    assign in8601_1 = {c5518};
    assign in8601_2 = {c5519};
    Full_Adder FA_8601(s8601, c8601, in8601_1, in8601_2, c5517);
    wire[0:0] s8602, in8602_1, in8602_2;
    wire c8602;
    assign in8602_1 = {c5521};
    assign in8602_2 = {s5522[0]};
    Full_Adder FA_8602(s8602, c8602, in8602_1, in8602_2, c5520);
    wire[0:0] s8603, in8603_1, in8603_2;
    wire c8603;
    assign in8603_1 = {s5524[0]};
    assign in8603_2 = {s5525[0]};
    Full_Adder FA_8603(s8603, c8603, in8603_1, in8603_2, s5523[0]);
    wire[0:0] s8604, in8604_1, in8604_2;
    wire c8604;
    assign in8604_1 = {s5527[0]};
    assign in8604_2 = {s5528[0]};
    Full_Adder FA_8604(s8604, c8604, in8604_1, in8604_2, s5526[0]);
    wire[0:0] s8605, in8605_1, in8605_2;
    wire c8605;
    assign in8605_1 = {s5530[0]};
    assign in8605_2 = {s5531[0]};
    Full_Adder FA_8605(s8605, c8605, in8605_1, in8605_2, s5529[0]);
    wire[0:0] s8606, in8606_1, in8606_2;
    wire c8606;
    assign in8606_1 = {s5533[0]};
    assign in8606_2 = {s5534[0]};
    Full_Adder FA_8606(s8606, c8606, in8606_1, in8606_2, s5532[0]);
    wire[0:0] s8607, in8607_1, in8607_2;
    wire c8607;
    assign in8607_1 = {s5536[0]};
    assign in8607_2 = {s5537[0]};
    Full_Adder FA_8607(s8607, c8607, in8607_1, in8607_2, s5535[0]);
    wire[0:0] s8608, in8608_1, in8608_2;
    wire c8608;
    assign in8608_1 = {s5539[0]};
    assign in8608_2 = {s5540[0]};
    Full_Adder FA_8608(s8608, c8608, in8608_1, in8608_2, s5538[0]);
    wire[0:0] s8609, in8609_1, in8609_2;
    wire c8609;
    assign in8609_1 = {c5522};
    assign in8609_2 = {c5523};
    Full_Adder FA_8609(s8609, c8609, in8609_1, in8609_2, s2037[0]);
    wire[0:0] s8610, in8610_1, in8610_2;
    wire c8610;
    assign in8610_1 = {c5525};
    assign in8610_2 = {c5526};
    Full_Adder FA_8610(s8610, c8610, in8610_1, in8610_2, c5524);
    wire[0:0] s8611, in8611_1, in8611_2;
    wire c8611;
    assign in8611_1 = {c5528};
    assign in8611_2 = {c5529};
    Full_Adder FA_8611(s8611, c8611, in8611_1, in8611_2, c5527);
    wire[0:0] s8612, in8612_1, in8612_2;
    wire c8612;
    assign in8612_1 = {c5531};
    assign in8612_2 = {c5532};
    Full_Adder FA_8612(s8612, c8612, in8612_1, in8612_2, c5530);
    wire[0:0] s8613, in8613_1, in8613_2;
    wire c8613;
    assign in8613_1 = {c5534};
    assign in8613_2 = {c5535};
    Full_Adder FA_8613(s8613, c8613, in8613_1, in8613_2, c5533);
    wire[0:0] s8614, in8614_1, in8614_2;
    wire c8614;
    assign in8614_1 = {c5537};
    assign in8614_2 = {c5538};
    Full_Adder FA_8614(s8614, c8614, in8614_1, in8614_2, c5536);
    wire[0:0] s8615, in8615_1, in8615_2;
    wire c8615;
    assign in8615_1 = {c5540};
    assign in8615_2 = {s5541[0]};
    Full_Adder FA_8615(s8615, c8615, in8615_1, in8615_2, c5539);
    wire[0:0] s8616, in8616_1, in8616_2;
    wire c8616;
    assign in8616_1 = {s5543[0]};
    assign in8616_2 = {s5544[0]};
    Full_Adder FA_8616(s8616, c8616, in8616_1, in8616_2, s5542[0]);
    wire[0:0] s8617, in8617_1, in8617_2;
    wire c8617;
    assign in8617_1 = {s5546[0]};
    assign in8617_2 = {s5547[0]};
    Full_Adder FA_8617(s8617, c8617, in8617_1, in8617_2, s5545[0]);
    wire[0:0] s8618, in8618_1, in8618_2;
    wire c8618;
    assign in8618_1 = {s5549[0]};
    assign in8618_2 = {s5550[0]};
    Full_Adder FA_8618(s8618, c8618, in8618_1, in8618_2, s5548[0]);
    wire[0:0] s8619, in8619_1, in8619_2;
    wire c8619;
    assign in8619_1 = {s5552[0]};
    assign in8619_2 = {s5553[0]};
    Full_Adder FA_8619(s8619, c8619, in8619_1, in8619_2, s5551[0]);
    wire[0:0] s8620, in8620_1, in8620_2;
    wire c8620;
    assign in8620_1 = {s5555[0]};
    assign in8620_2 = {s5556[0]};
    Full_Adder FA_8620(s8620, c8620, in8620_1, in8620_2, s5554[0]);
    wire[0:0] s8621, in8621_1, in8621_2;
    wire c8621;
    assign in8621_1 = {s5558[0]};
    assign in8621_2 = {s5559[0]};
    Full_Adder FA_8621(s8621, c8621, in8621_1, in8621_2, s5557[0]);
    wire[0:0] s8622, in8622_1, in8622_2;
    wire c8622;
    assign in8622_1 = {c5541};
    assign in8622_2 = {c5542};
    Full_Adder FA_8622(s8622, c8622, in8622_1, in8622_2, s2059[0]);
    wire[0:0] s8623, in8623_1, in8623_2;
    wire c8623;
    assign in8623_1 = {c5544};
    assign in8623_2 = {c5545};
    Full_Adder FA_8623(s8623, c8623, in8623_1, in8623_2, c5543);
    wire[0:0] s8624, in8624_1, in8624_2;
    wire c8624;
    assign in8624_1 = {c5547};
    assign in8624_2 = {c5548};
    Full_Adder FA_8624(s8624, c8624, in8624_1, in8624_2, c5546);
    wire[0:0] s8625, in8625_1, in8625_2;
    wire c8625;
    assign in8625_1 = {c5550};
    assign in8625_2 = {c5551};
    Full_Adder FA_8625(s8625, c8625, in8625_1, in8625_2, c5549);
    wire[0:0] s8626, in8626_1, in8626_2;
    wire c8626;
    assign in8626_1 = {c5553};
    assign in8626_2 = {c5554};
    Full_Adder FA_8626(s8626, c8626, in8626_1, in8626_2, c5552);
    wire[0:0] s8627, in8627_1, in8627_2;
    wire c8627;
    assign in8627_1 = {c5556};
    assign in8627_2 = {c5557};
    Full_Adder FA_8627(s8627, c8627, in8627_1, in8627_2, c5555);
    wire[0:0] s8628, in8628_1, in8628_2;
    wire c8628;
    assign in8628_1 = {c5559};
    assign in8628_2 = {s5560[0]};
    Full_Adder FA_8628(s8628, c8628, in8628_1, in8628_2, c5558);
    wire[0:0] s8629, in8629_1, in8629_2;
    wire c8629;
    assign in8629_1 = {s5562[0]};
    assign in8629_2 = {s5563[0]};
    Full_Adder FA_8629(s8629, c8629, in8629_1, in8629_2, s5561[0]);
    wire[0:0] s8630, in8630_1, in8630_2;
    wire c8630;
    assign in8630_1 = {s5565[0]};
    assign in8630_2 = {s5566[0]};
    Full_Adder FA_8630(s8630, c8630, in8630_1, in8630_2, s5564[0]);
    wire[0:0] s8631, in8631_1, in8631_2;
    wire c8631;
    assign in8631_1 = {s5568[0]};
    assign in8631_2 = {s5569[0]};
    Full_Adder FA_8631(s8631, c8631, in8631_1, in8631_2, s5567[0]);
    wire[0:0] s8632, in8632_1, in8632_2;
    wire c8632;
    assign in8632_1 = {s5571[0]};
    assign in8632_2 = {s5572[0]};
    Full_Adder FA_8632(s8632, c8632, in8632_1, in8632_2, s5570[0]);
    wire[0:0] s8633, in8633_1, in8633_2;
    wire c8633;
    assign in8633_1 = {s5574[0]};
    assign in8633_2 = {s5575[0]};
    Full_Adder FA_8633(s8633, c8633, in8633_1, in8633_2, s5573[0]);
    wire[0:0] s8634, in8634_1, in8634_2;
    wire c8634;
    assign in8634_1 = {s5577[0]};
    assign in8634_2 = {s5578[0]};
    Full_Adder FA_8634(s8634, c8634, in8634_1, in8634_2, s5576[0]);
    wire[0:0] s8635, in8635_1, in8635_2;
    wire c8635;
    assign in8635_1 = {c5560};
    assign in8635_2 = {c5561};
    Full_Adder FA_8635(s8635, c8635, in8635_1, in8635_2, s2082[0]);
    wire[0:0] s8636, in8636_1, in8636_2;
    wire c8636;
    assign in8636_1 = {c5563};
    assign in8636_2 = {c5564};
    Full_Adder FA_8636(s8636, c8636, in8636_1, in8636_2, c5562);
    wire[0:0] s8637, in8637_1, in8637_2;
    wire c8637;
    assign in8637_1 = {c5566};
    assign in8637_2 = {c5567};
    Full_Adder FA_8637(s8637, c8637, in8637_1, in8637_2, c5565);
    wire[0:0] s8638, in8638_1, in8638_2;
    wire c8638;
    assign in8638_1 = {c5569};
    assign in8638_2 = {c5570};
    Full_Adder FA_8638(s8638, c8638, in8638_1, in8638_2, c5568);
    wire[0:0] s8639, in8639_1, in8639_2;
    wire c8639;
    assign in8639_1 = {c5572};
    assign in8639_2 = {c5573};
    Full_Adder FA_8639(s8639, c8639, in8639_1, in8639_2, c5571);
    wire[0:0] s8640, in8640_1, in8640_2;
    wire c8640;
    assign in8640_1 = {c5575};
    assign in8640_2 = {c5576};
    Full_Adder FA_8640(s8640, c8640, in8640_1, in8640_2, c5574);
    wire[0:0] s8641, in8641_1, in8641_2;
    wire c8641;
    assign in8641_1 = {c5578};
    assign in8641_2 = {s5579[0]};
    Full_Adder FA_8641(s8641, c8641, in8641_1, in8641_2, c5577);
    wire[0:0] s8642, in8642_1, in8642_2;
    wire c8642;
    assign in8642_1 = {s5581[0]};
    assign in8642_2 = {s5582[0]};
    Full_Adder FA_8642(s8642, c8642, in8642_1, in8642_2, s5580[0]);
    wire[0:0] s8643, in8643_1, in8643_2;
    wire c8643;
    assign in8643_1 = {s5584[0]};
    assign in8643_2 = {s5585[0]};
    Full_Adder FA_8643(s8643, c8643, in8643_1, in8643_2, s5583[0]);
    wire[0:0] s8644, in8644_1, in8644_2;
    wire c8644;
    assign in8644_1 = {s5587[0]};
    assign in8644_2 = {s5588[0]};
    Full_Adder FA_8644(s8644, c8644, in8644_1, in8644_2, s5586[0]);
    wire[0:0] s8645, in8645_1, in8645_2;
    wire c8645;
    assign in8645_1 = {s5590[0]};
    assign in8645_2 = {s5591[0]};
    Full_Adder FA_8645(s8645, c8645, in8645_1, in8645_2, s5589[0]);
    wire[0:0] s8646, in8646_1, in8646_2;
    wire c8646;
    assign in8646_1 = {s5593[0]};
    assign in8646_2 = {s5594[0]};
    Full_Adder FA_8646(s8646, c8646, in8646_1, in8646_2, s5592[0]);
    wire[0:0] s8647, in8647_1, in8647_2;
    wire c8647;
    assign in8647_1 = {s5596[0]};
    assign in8647_2 = {s5597[0]};
    Full_Adder FA_8647(s8647, c8647, in8647_1, in8647_2, s5595[0]);
    wire[0:0] s8648, in8648_1, in8648_2;
    wire c8648;
    assign in8648_1 = {c5579};
    assign in8648_2 = {c5580};
    Full_Adder FA_8648(s8648, c8648, in8648_1, in8648_2, s2106[0]);
    wire[0:0] s8649, in8649_1, in8649_2;
    wire c8649;
    assign in8649_1 = {c5582};
    assign in8649_2 = {c5583};
    Full_Adder FA_8649(s8649, c8649, in8649_1, in8649_2, c5581);
    wire[0:0] s8650, in8650_1, in8650_2;
    wire c8650;
    assign in8650_1 = {c5585};
    assign in8650_2 = {c5586};
    Full_Adder FA_8650(s8650, c8650, in8650_1, in8650_2, c5584);
    wire[0:0] s8651, in8651_1, in8651_2;
    wire c8651;
    assign in8651_1 = {c5588};
    assign in8651_2 = {c5589};
    Full_Adder FA_8651(s8651, c8651, in8651_1, in8651_2, c5587);
    wire[0:0] s8652, in8652_1, in8652_2;
    wire c8652;
    assign in8652_1 = {c5591};
    assign in8652_2 = {c5592};
    Full_Adder FA_8652(s8652, c8652, in8652_1, in8652_2, c5590);
    wire[0:0] s8653, in8653_1, in8653_2;
    wire c8653;
    assign in8653_1 = {c5594};
    assign in8653_2 = {c5595};
    Full_Adder FA_8653(s8653, c8653, in8653_1, in8653_2, c5593);
    wire[0:0] s8654, in8654_1, in8654_2;
    wire c8654;
    assign in8654_1 = {c5597};
    assign in8654_2 = {s5598[0]};
    Full_Adder FA_8654(s8654, c8654, in8654_1, in8654_2, c5596);
    wire[0:0] s8655, in8655_1, in8655_2;
    wire c8655;
    assign in8655_1 = {s5600[0]};
    assign in8655_2 = {s5601[0]};
    Full_Adder FA_8655(s8655, c8655, in8655_1, in8655_2, s5599[0]);
    wire[0:0] s8656, in8656_1, in8656_2;
    wire c8656;
    assign in8656_1 = {s5603[0]};
    assign in8656_2 = {s5604[0]};
    Full_Adder FA_8656(s8656, c8656, in8656_1, in8656_2, s5602[0]);
    wire[0:0] s8657, in8657_1, in8657_2;
    wire c8657;
    assign in8657_1 = {s5606[0]};
    assign in8657_2 = {s5607[0]};
    Full_Adder FA_8657(s8657, c8657, in8657_1, in8657_2, s5605[0]);
    wire[0:0] s8658, in8658_1, in8658_2;
    wire c8658;
    assign in8658_1 = {s5609[0]};
    assign in8658_2 = {s5610[0]};
    Full_Adder FA_8658(s8658, c8658, in8658_1, in8658_2, s5608[0]);
    wire[0:0] s8659, in8659_1, in8659_2;
    wire c8659;
    assign in8659_1 = {s5612[0]};
    assign in8659_2 = {s5613[0]};
    Full_Adder FA_8659(s8659, c8659, in8659_1, in8659_2, s5611[0]);
    wire[0:0] s8660, in8660_1, in8660_2;
    wire c8660;
    assign in8660_1 = {s5615[0]};
    assign in8660_2 = {s5616[0]};
    Full_Adder FA_8660(s8660, c8660, in8660_1, in8660_2, s5614[0]);
    wire[0:0] s8661, in8661_1, in8661_2;
    wire c8661;
    assign in8661_1 = {c5598};
    assign in8661_2 = {c5599};
    Full_Adder FA_8661(s8661, c8661, in8661_1, in8661_2, s2131[0]);
    wire[0:0] s8662, in8662_1, in8662_2;
    wire c8662;
    assign in8662_1 = {c5601};
    assign in8662_2 = {c5602};
    Full_Adder FA_8662(s8662, c8662, in8662_1, in8662_2, c5600);
    wire[0:0] s8663, in8663_1, in8663_2;
    wire c8663;
    assign in8663_1 = {c5604};
    assign in8663_2 = {c5605};
    Full_Adder FA_8663(s8663, c8663, in8663_1, in8663_2, c5603);
    wire[0:0] s8664, in8664_1, in8664_2;
    wire c8664;
    assign in8664_1 = {c5607};
    assign in8664_2 = {c5608};
    Full_Adder FA_8664(s8664, c8664, in8664_1, in8664_2, c5606);
    wire[0:0] s8665, in8665_1, in8665_2;
    wire c8665;
    assign in8665_1 = {c5610};
    assign in8665_2 = {c5611};
    Full_Adder FA_8665(s8665, c8665, in8665_1, in8665_2, c5609);
    wire[0:0] s8666, in8666_1, in8666_2;
    wire c8666;
    assign in8666_1 = {c5613};
    assign in8666_2 = {c5614};
    Full_Adder FA_8666(s8666, c8666, in8666_1, in8666_2, c5612);
    wire[0:0] s8667, in8667_1, in8667_2;
    wire c8667;
    assign in8667_1 = {c5616};
    assign in8667_2 = {s5617[0]};
    Full_Adder FA_8667(s8667, c8667, in8667_1, in8667_2, c5615);
    wire[0:0] s8668, in8668_1, in8668_2;
    wire c8668;
    assign in8668_1 = {s5619[0]};
    assign in8668_2 = {s5620[0]};
    Full_Adder FA_8668(s8668, c8668, in8668_1, in8668_2, s5618[0]);
    wire[0:0] s8669, in8669_1, in8669_2;
    wire c8669;
    assign in8669_1 = {s5622[0]};
    assign in8669_2 = {s5623[0]};
    Full_Adder FA_8669(s8669, c8669, in8669_1, in8669_2, s5621[0]);
    wire[0:0] s8670, in8670_1, in8670_2;
    wire c8670;
    assign in8670_1 = {s5625[0]};
    assign in8670_2 = {s5626[0]};
    Full_Adder FA_8670(s8670, c8670, in8670_1, in8670_2, s5624[0]);
    wire[0:0] s8671, in8671_1, in8671_2;
    wire c8671;
    assign in8671_1 = {s5628[0]};
    assign in8671_2 = {s5629[0]};
    Full_Adder FA_8671(s8671, c8671, in8671_1, in8671_2, s5627[0]);
    wire[0:0] s8672, in8672_1, in8672_2;
    wire c8672;
    assign in8672_1 = {s5631[0]};
    assign in8672_2 = {s5632[0]};
    Full_Adder FA_8672(s8672, c8672, in8672_1, in8672_2, s5630[0]);
    wire[0:0] s8673, in8673_1, in8673_2;
    wire c8673;
    assign in8673_1 = {s5634[0]};
    assign in8673_2 = {s5635[0]};
    Full_Adder FA_8673(s8673, c8673, in8673_1, in8673_2, s5633[0]);
    wire[0:0] s8674, in8674_1, in8674_2;
    wire c8674;
    assign in8674_1 = {c5617};
    assign in8674_2 = {c5618};
    Full_Adder FA_8674(s8674, c8674, in8674_1, in8674_2, s2157[0]);
    wire[0:0] s8675, in8675_1, in8675_2;
    wire c8675;
    assign in8675_1 = {c5620};
    assign in8675_2 = {c5621};
    Full_Adder FA_8675(s8675, c8675, in8675_1, in8675_2, c5619);
    wire[0:0] s8676, in8676_1, in8676_2;
    wire c8676;
    assign in8676_1 = {c5623};
    assign in8676_2 = {c5624};
    Full_Adder FA_8676(s8676, c8676, in8676_1, in8676_2, c5622);
    wire[0:0] s8677, in8677_1, in8677_2;
    wire c8677;
    assign in8677_1 = {c5626};
    assign in8677_2 = {c5627};
    Full_Adder FA_8677(s8677, c8677, in8677_1, in8677_2, c5625);
    wire[0:0] s8678, in8678_1, in8678_2;
    wire c8678;
    assign in8678_1 = {c5629};
    assign in8678_2 = {c5630};
    Full_Adder FA_8678(s8678, c8678, in8678_1, in8678_2, c5628);
    wire[0:0] s8679, in8679_1, in8679_2;
    wire c8679;
    assign in8679_1 = {c5632};
    assign in8679_2 = {c5633};
    Full_Adder FA_8679(s8679, c8679, in8679_1, in8679_2, c5631);
    wire[0:0] s8680, in8680_1, in8680_2;
    wire c8680;
    assign in8680_1 = {c5635};
    assign in8680_2 = {s5636[0]};
    Full_Adder FA_8680(s8680, c8680, in8680_1, in8680_2, c5634);
    wire[0:0] s8681, in8681_1, in8681_2;
    wire c8681;
    assign in8681_1 = {s5638[0]};
    assign in8681_2 = {s5639[0]};
    Full_Adder FA_8681(s8681, c8681, in8681_1, in8681_2, s5637[0]);
    wire[0:0] s8682, in8682_1, in8682_2;
    wire c8682;
    assign in8682_1 = {s5641[0]};
    assign in8682_2 = {s5642[0]};
    Full_Adder FA_8682(s8682, c8682, in8682_1, in8682_2, s5640[0]);
    wire[0:0] s8683, in8683_1, in8683_2;
    wire c8683;
    assign in8683_1 = {s5644[0]};
    assign in8683_2 = {s5645[0]};
    Full_Adder FA_8683(s8683, c8683, in8683_1, in8683_2, s5643[0]);
    wire[0:0] s8684, in8684_1, in8684_2;
    wire c8684;
    assign in8684_1 = {s5647[0]};
    assign in8684_2 = {s5648[0]};
    Full_Adder FA_8684(s8684, c8684, in8684_1, in8684_2, s5646[0]);
    wire[0:0] s8685, in8685_1, in8685_2;
    wire c8685;
    assign in8685_1 = {s5650[0]};
    assign in8685_2 = {s5651[0]};
    Full_Adder FA_8685(s8685, c8685, in8685_1, in8685_2, s5649[0]);
    wire[0:0] s8686, in8686_1, in8686_2;
    wire c8686;
    assign in8686_1 = {s5653[0]};
    assign in8686_2 = {s5654[0]};
    Full_Adder FA_8686(s8686, c8686, in8686_1, in8686_2, s5652[0]);
    wire[0:0] s8687, in8687_1, in8687_2;
    wire c8687;
    assign in8687_1 = {c5636};
    assign in8687_2 = {c5637};
    Full_Adder FA_8687(s8687, c8687, in8687_1, in8687_2, s2184[0]);
    wire[0:0] s8688, in8688_1, in8688_2;
    wire c8688;
    assign in8688_1 = {c5639};
    assign in8688_2 = {c5640};
    Full_Adder FA_8688(s8688, c8688, in8688_1, in8688_2, c5638);
    wire[0:0] s8689, in8689_1, in8689_2;
    wire c8689;
    assign in8689_1 = {c5642};
    assign in8689_2 = {c5643};
    Full_Adder FA_8689(s8689, c8689, in8689_1, in8689_2, c5641);
    wire[0:0] s8690, in8690_1, in8690_2;
    wire c8690;
    assign in8690_1 = {c5645};
    assign in8690_2 = {c5646};
    Full_Adder FA_8690(s8690, c8690, in8690_1, in8690_2, c5644);
    wire[0:0] s8691, in8691_1, in8691_2;
    wire c8691;
    assign in8691_1 = {c5648};
    assign in8691_2 = {c5649};
    Full_Adder FA_8691(s8691, c8691, in8691_1, in8691_2, c5647);
    wire[0:0] s8692, in8692_1, in8692_2;
    wire c8692;
    assign in8692_1 = {c5651};
    assign in8692_2 = {c5652};
    Full_Adder FA_8692(s8692, c8692, in8692_1, in8692_2, c5650);
    wire[0:0] s8693, in8693_1, in8693_2;
    wire c8693;
    assign in8693_1 = {c5654};
    assign in8693_2 = {s5655[0]};
    Full_Adder FA_8693(s8693, c8693, in8693_1, in8693_2, c5653);
    wire[0:0] s8694, in8694_1, in8694_2;
    wire c8694;
    assign in8694_1 = {s5657[0]};
    assign in8694_2 = {s5658[0]};
    Full_Adder FA_8694(s8694, c8694, in8694_1, in8694_2, s5656[0]);
    wire[0:0] s8695, in8695_1, in8695_2;
    wire c8695;
    assign in8695_1 = {s5660[0]};
    assign in8695_2 = {s5661[0]};
    Full_Adder FA_8695(s8695, c8695, in8695_1, in8695_2, s5659[0]);
    wire[0:0] s8696, in8696_1, in8696_2;
    wire c8696;
    assign in8696_1 = {s5663[0]};
    assign in8696_2 = {s5664[0]};
    Full_Adder FA_8696(s8696, c8696, in8696_1, in8696_2, s5662[0]);
    wire[0:0] s8697, in8697_1, in8697_2;
    wire c8697;
    assign in8697_1 = {s5666[0]};
    assign in8697_2 = {s5667[0]};
    Full_Adder FA_8697(s8697, c8697, in8697_1, in8697_2, s5665[0]);
    wire[0:0] s8698, in8698_1, in8698_2;
    wire c8698;
    assign in8698_1 = {s5669[0]};
    assign in8698_2 = {s5670[0]};
    Full_Adder FA_8698(s8698, c8698, in8698_1, in8698_2, s5668[0]);
    wire[0:0] s8699, in8699_1, in8699_2;
    wire c8699;
    assign in8699_1 = {s5672[0]};
    assign in8699_2 = {s5673[0]};
    Full_Adder FA_8699(s8699, c8699, in8699_1, in8699_2, s5671[0]);
    wire[0:0] s8700, in8700_1, in8700_2;
    wire c8700;
    assign in8700_1 = {c5655};
    assign in8700_2 = {c5656};
    Full_Adder FA_8700(s8700, c8700, in8700_1, in8700_2, s2212[0]);
    wire[0:0] s8701, in8701_1, in8701_2;
    wire c8701;
    assign in8701_1 = {c5658};
    assign in8701_2 = {c5659};
    Full_Adder FA_8701(s8701, c8701, in8701_1, in8701_2, c5657);
    wire[0:0] s8702, in8702_1, in8702_2;
    wire c8702;
    assign in8702_1 = {c5661};
    assign in8702_2 = {c5662};
    Full_Adder FA_8702(s8702, c8702, in8702_1, in8702_2, c5660);
    wire[0:0] s8703, in8703_1, in8703_2;
    wire c8703;
    assign in8703_1 = {c5664};
    assign in8703_2 = {c5665};
    Full_Adder FA_8703(s8703, c8703, in8703_1, in8703_2, c5663);
    wire[0:0] s8704, in8704_1, in8704_2;
    wire c8704;
    assign in8704_1 = {c5667};
    assign in8704_2 = {c5668};
    Full_Adder FA_8704(s8704, c8704, in8704_1, in8704_2, c5666);
    wire[0:0] s8705, in8705_1, in8705_2;
    wire c8705;
    assign in8705_1 = {c5670};
    assign in8705_2 = {c5671};
    Full_Adder FA_8705(s8705, c8705, in8705_1, in8705_2, c5669);
    wire[0:0] s8706, in8706_1, in8706_2;
    wire c8706;
    assign in8706_1 = {c5673};
    assign in8706_2 = {s5674[0]};
    Full_Adder FA_8706(s8706, c8706, in8706_1, in8706_2, c5672);
    wire[0:0] s8707, in8707_1, in8707_2;
    wire c8707;
    assign in8707_1 = {s5676[0]};
    assign in8707_2 = {s5677[0]};
    Full_Adder FA_8707(s8707, c8707, in8707_1, in8707_2, s5675[0]);
    wire[0:0] s8708, in8708_1, in8708_2;
    wire c8708;
    assign in8708_1 = {s5679[0]};
    assign in8708_2 = {s5680[0]};
    Full_Adder FA_8708(s8708, c8708, in8708_1, in8708_2, s5678[0]);
    wire[0:0] s8709, in8709_1, in8709_2;
    wire c8709;
    assign in8709_1 = {s5682[0]};
    assign in8709_2 = {s5683[0]};
    Full_Adder FA_8709(s8709, c8709, in8709_1, in8709_2, s5681[0]);
    wire[0:0] s8710, in8710_1, in8710_2;
    wire c8710;
    assign in8710_1 = {s5685[0]};
    assign in8710_2 = {s5686[0]};
    Full_Adder FA_8710(s8710, c8710, in8710_1, in8710_2, s5684[0]);
    wire[0:0] s8711, in8711_1, in8711_2;
    wire c8711;
    assign in8711_1 = {s5688[0]};
    assign in8711_2 = {s5689[0]};
    Full_Adder FA_8711(s8711, c8711, in8711_1, in8711_2, s5687[0]);
    wire[0:0] s8712, in8712_1, in8712_2;
    wire c8712;
    assign in8712_1 = {s5691[0]};
    assign in8712_2 = {s5692[0]};
    Full_Adder FA_8712(s8712, c8712, in8712_1, in8712_2, s5690[0]);
    wire[0:0] s8713, in8713_1, in8713_2;
    wire c8713;
    assign in8713_1 = {c5674};
    assign in8713_2 = {c5675};
    Full_Adder FA_8713(s8713, c8713, in8713_1, in8713_2, s2240[0]);
    wire[0:0] s8714, in8714_1, in8714_2;
    wire c8714;
    assign in8714_1 = {c5677};
    assign in8714_2 = {c5678};
    Full_Adder FA_8714(s8714, c8714, in8714_1, in8714_2, c5676);
    wire[0:0] s8715, in8715_1, in8715_2;
    wire c8715;
    assign in8715_1 = {c5680};
    assign in8715_2 = {c5681};
    Full_Adder FA_8715(s8715, c8715, in8715_1, in8715_2, c5679);
    wire[0:0] s8716, in8716_1, in8716_2;
    wire c8716;
    assign in8716_1 = {c5683};
    assign in8716_2 = {c5684};
    Full_Adder FA_8716(s8716, c8716, in8716_1, in8716_2, c5682);
    wire[0:0] s8717, in8717_1, in8717_2;
    wire c8717;
    assign in8717_1 = {c5686};
    assign in8717_2 = {c5687};
    Full_Adder FA_8717(s8717, c8717, in8717_1, in8717_2, c5685);
    wire[0:0] s8718, in8718_1, in8718_2;
    wire c8718;
    assign in8718_1 = {c5689};
    assign in8718_2 = {c5690};
    Full_Adder FA_8718(s8718, c8718, in8718_1, in8718_2, c5688);
    wire[0:0] s8719, in8719_1, in8719_2;
    wire c8719;
    assign in8719_1 = {c5692};
    assign in8719_2 = {s5693[0]};
    Full_Adder FA_8719(s8719, c8719, in8719_1, in8719_2, c5691);
    wire[0:0] s8720, in8720_1, in8720_2;
    wire c8720;
    assign in8720_1 = {s5695[0]};
    assign in8720_2 = {s5696[0]};
    Full_Adder FA_8720(s8720, c8720, in8720_1, in8720_2, s5694[0]);
    wire[0:0] s8721, in8721_1, in8721_2;
    wire c8721;
    assign in8721_1 = {s5698[0]};
    assign in8721_2 = {s5699[0]};
    Full_Adder FA_8721(s8721, c8721, in8721_1, in8721_2, s5697[0]);
    wire[0:0] s8722, in8722_1, in8722_2;
    wire c8722;
    assign in8722_1 = {s5701[0]};
    assign in8722_2 = {s5702[0]};
    Full_Adder FA_8722(s8722, c8722, in8722_1, in8722_2, s5700[0]);
    wire[0:0] s8723, in8723_1, in8723_2;
    wire c8723;
    assign in8723_1 = {s5704[0]};
    assign in8723_2 = {s5705[0]};
    Full_Adder FA_8723(s8723, c8723, in8723_1, in8723_2, s5703[0]);
    wire[0:0] s8724, in8724_1, in8724_2;
    wire c8724;
    assign in8724_1 = {s5707[0]};
    assign in8724_2 = {s5708[0]};
    Full_Adder FA_8724(s8724, c8724, in8724_1, in8724_2, s5706[0]);
    wire[0:0] s8725, in8725_1, in8725_2;
    wire c8725;
    assign in8725_1 = {s5710[0]};
    assign in8725_2 = {s5711[0]};
    Full_Adder FA_8725(s8725, c8725, in8725_1, in8725_2, s5709[0]);
    wire[0:0] s8726, in8726_1, in8726_2;
    wire c8726;
    assign in8726_1 = {c5693};
    assign in8726_2 = {c5694};
    Full_Adder FA_8726(s8726, c8726, in8726_1, in8726_2, s2268[0]);
    wire[0:0] s8727, in8727_1, in8727_2;
    wire c8727;
    assign in8727_1 = {c5696};
    assign in8727_2 = {c5697};
    Full_Adder FA_8727(s8727, c8727, in8727_1, in8727_2, c5695);
    wire[0:0] s8728, in8728_1, in8728_2;
    wire c8728;
    assign in8728_1 = {c5699};
    assign in8728_2 = {c5700};
    Full_Adder FA_8728(s8728, c8728, in8728_1, in8728_2, c5698);
    wire[0:0] s8729, in8729_1, in8729_2;
    wire c8729;
    assign in8729_1 = {c5702};
    assign in8729_2 = {c5703};
    Full_Adder FA_8729(s8729, c8729, in8729_1, in8729_2, c5701);
    wire[0:0] s8730, in8730_1, in8730_2;
    wire c8730;
    assign in8730_1 = {c5705};
    assign in8730_2 = {c5706};
    Full_Adder FA_8730(s8730, c8730, in8730_1, in8730_2, c5704);
    wire[0:0] s8731, in8731_1, in8731_2;
    wire c8731;
    assign in8731_1 = {c5708};
    assign in8731_2 = {c5709};
    Full_Adder FA_8731(s8731, c8731, in8731_1, in8731_2, c5707);
    wire[0:0] s8732, in8732_1, in8732_2;
    wire c8732;
    assign in8732_1 = {c5711};
    assign in8732_2 = {s5712[0]};
    Full_Adder FA_8732(s8732, c8732, in8732_1, in8732_2, c5710);
    wire[0:0] s8733, in8733_1, in8733_2;
    wire c8733;
    assign in8733_1 = {s5714[0]};
    assign in8733_2 = {s5715[0]};
    Full_Adder FA_8733(s8733, c8733, in8733_1, in8733_2, s5713[0]);
    wire[0:0] s8734, in8734_1, in8734_2;
    wire c8734;
    assign in8734_1 = {s5717[0]};
    assign in8734_2 = {s5718[0]};
    Full_Adder FA_8734(s8734, c8734, in8734_1, in8734_2, s5716[0]);
    wire[0:0] s8735, in8735_1, in8735_2;
    wire c8735;
    assign in8735_1 = {s5720[0]};
    assign in8735_2 = {s5721[0]};
    Full_Adder FA_8735(s8735, c8735, in8735_1, in8735_2, s5719[0]);
    wire[0:0] s8736, in8736_1, in8736_2;
    wire c8736;
    assign in8736_1 = {s5723[0]};
    assign in8736_2 = {s5724[0]};
    Full_Adder FA_8736(s8736, c8736, in8736_1, in8736_2, s5722[0]);
    wire[0:0] s8737, in8737_1, in8737_2;
    wire c8737;
    assign in8737_1 = {s5726[0]};
    assign in8737_2 = {s5727[0]};
    Full_Adder FA_8737(s8737, c8737, in8737_1, in8737_2, s5725[0]);
    wire[0:0] s8738, in8738_1, in8738_2;
    wire c8738;
    assign in8738_1 = {s5729[0]};
    assign in8738_2 = {s5730[0]};
    Full_Adder FA_8738(s8738, c8738, in8738_1, in8738_2, s5728[0]);
    wire[0:0] s8739, in8739_1, in8739_2;
    wire c8739;
    assign in8739_1 = {c5712};
    assign in8739_2 = {c5713};
    Full_Adder FA_8739(s8739, c8739, in8739_1, in8739_2, s2296[0]);
    wire[0:0] s8740, in8740_1, in8740_2;
    wire c8740;
    assign in8740_1 = {c5715};
    assign in8740_2 = {c5716};
    Full_Adder FA_8740(s8740, c8740, in8740_1, in8740_2, c5714);
    wire[0:0] s8741, in8741_1, in8741_2;
    wire c8741;
    assign in8741_1 = {c5718};
    assign in8741_2 = {c5719};
    Full_Adder FA_8741(s8741, c8741, in8741_1, in8741_2, c5717);
    wire[0:0] s8742, in8742_1, in8742_2;
    wire c8742;
    assign in8742_1 = {c5721};
    assign in8742_2 = {c5722};
    Full_Adder FA_8742(s8742, c8742, in8742_1, in8742_2, c5720);
    wire[0:0] s8743, in8743_1, in8743_2;
    wire c8743;
    assign in8743_1 = {c5724};
    assign in8743_2 = {c5725};
    Full_Adder FA_8743(s8743, c8743, in8743_1, in8743_2, c5723);
    wire[0:0] s8744, in8744_1, in8744_2;
    wire c8744;
    assign in8744_1 = {c5727};
    assign in8744_2 = {c5728};
    Full_Adder FA_8744(s8744, c8744, in8744_1, in8744_2, c5726);
    wire[0:0] s8745, in8745_1, in8745_2;
    wire c8745;
    assign in8745_1 = {c5730};
    assign in8745_2 = {s5731[0]};
    Full_Adder FA_8745(s8745, c8745, in8745_1, in8745_2, c5729);
    wire[0:0] s8746, in8746_1, in8746_2;
    wire c8746;
    assign in8746_1 = {s5733[0]};
    assign in8746_2 = {s5734[0]};
    Full_Adder FA_8746(s8746, c8746, in8746_1, in8746_2, s5732[0]);
    wire[0:0] s8747, in8747_1, in8747_2;
    wire c8747;
    assign in8747_1 = {s5736[0]};
    assign in8747_2 = {s5737[0]};
    Full_Adder FA_8747(s8747, c8747, in8747_1, in8747_2, s5735[0]);
    wire[0:0] s8748, in8748_1, in8748_2;
    wire c8748;
    assign in8748_1 = {s5739[0]};
    assign in8748_2 = {s5740[0]};
    Full_Adder FA_8748(s8748, c8748, in8748_1, in8748_2, s5738[0]);
    wire[0:0] s8749, in8749_1, in8749_2;
    wire c8749;
    assign in8749_1 = {s5742[0]};
    assign in8749_2 = {s5743[0]};
    Full_Adder FA_8749(s8749, c8749, in8749_1, in8749_2, s5741[0]);
    wire[0:0] s8750, in8750_1, in8750_2;
    wire c8750;
    assign in8750_1 = {s5745[0]};
    assign in8750_2 = {s5746[0]};
    Full_Adder FA_8750(s8750, c8750, in8750_1, in8750_2, s5744[0]);
    wire[0:0] s8751, in8751_1, in8751_2;
    wire c8751;
    assign in8751_1 = {s5748[0]};
    assign in8751_2 = {s5749[0]};
    Full_Adder FA_8751(s8751, c8751, in8751_1, in8751_2, s5747[0]);
    wire[0:0] s8752, in8752_1, in8752_2;
    wire c8752;
    assign in8752_1 = {c5731};
    assign in8752_2 = {c5732};
    Full_Adder FA_8752(s8752, c8752, in8752_1, in8752_2, s2324[0]);
    wire[0:0] s8753, in8753_1, in8753_2;
    wire c8753;
    assign in8753_1 = {c5734};
    assign in8753_2 = {c5735};
    Full_Adder FA_8753(s8753, c8753, in8753_1, in8753_2, c5733);
    wire[0:0] s8754, in8754_1, in8754_2;
    wire c8754;
    assign in8754_1 = {c5737};
    assign in8754_2 = {c5738};
    Full_Adder FA_8754(s8754, c8754, in8754_1, in8754_2, c5736);
    wire[0:0] s8755, in8755_1, in8755_2;
    wire c8755;
    assign in8755_1 = {c5740};
    assign in8755_2 = {c5741};
    Full_Adder FA_8755(s8755, c8755, in8755_1, in8755_2, c5739);
    wire[0:0] s8756, in8756_1, in8756_2;
    wire c8756;
    assign in8756_1 = {c5743};
    assign in8756_2 = {c5744};
    Full_Adder FA_8756(s8756, c8756, in8756_1, in8756_2, c5742);
    wire[0:0] s8757, in8757_1, in8757_2;
    wire c8757;
    assign in8757_1 = {c5746};
    assign in8757_2 = {c5747};
    Full_Adder FA_8757(s8757, c8757, in8757_1, in8757_2, c5745);
    wire[0:0] s8758, in8758_1, in8758_2;
    wire c8758;
    assign in8758_1 = {c5749};
    assign in8758_2 = {s5750[0]};
    Full_Adder FA_8758(s8758, c8758, in8758_1, in8758_2, c5748);
    wire[0:0] s8759, in8759_1, in8759_2;
    wire c8759;
    assign in8759_1 = {s5752[0]};
    assign in8759_2 = {s5753[0]};
    Full_Adder FA_8759(s8759, c8759, in8759_1, in8759_2, s5751[0]);
    wire[0:0] s8760, in8760_1, in8760_2;
    wire c8760;
    assign in8760_1 = {s5755[0]};
    assign in8760_2 = {s5756[0]};
    Full_Adder FA_8760(s8760, c8760, in8760_1, in8760_2, s5754[0]);
    wire[0:0] s8761, in8761_1, in8761_2;
    wire c8761;
    assign in8761_1 = {s5758[0]};
    assign in8761_2 = {s5759[0]};
    Full_Adder FA_8761(s8761, c8761, in8761_1, in8761_2, s5757[0]);
    wire[0:0] s8762, in8762_1, in8762_2;
    wire c8762;
    assign in8762_1 = {s5761[0]};
    assign in8762_2 = {s5762[0]};
    Full_Adder FA_8762(s8762, c8762, in8762_1, in8762_2, s5760[0]);
    wire[0:0] s8763, in8763_1, in8763_2;
    wire c8763;
    assign in8763_1 = {s5764[0]};
    assign in8763_2 = {s5765[0]};
    Full_Adder FA_8763(s8763, c8763, in8763_1, in8763_2, s5763[0]);
    wire[0:0] s8764, in8764_1, in8764_2;
    wire c8764;
    assign in8764_1 = {s5767[0]};
    assign in8764_2 = {s5768[0]};
    Full_Adder FA_8764(s8764, c8764, in8764_1, in8764_2, s5766[0]);
    wire[0:0] s8765, in8765_1, in8765_2;
    wire c8765;
    assign in8765_1 = {c5750};
    assign in8765_2 = {c5751};
    Full_Adder FA_8765(s8765, c8765, in8765_1, in8765_2, s2352[0]);
    wire[0:0] s8766, in8766_1, in8766_2;
    wire c8766;
    assign in8766_1 = {c5753};
    assign in8766_2 = {c5754};
    Full_Adder FA_8766(s8766, c8766, in8766_1, in8766_2, c5752);
    wire[0:0] s8767, in8767_1, in8767_2;
    wire c8767;
    assign in8767_1 = {c5756};
    assign in8767_2 = {c5757};
    Full_Adder FA_8767(s8767, c8767, in8767_1, in8767_2, c5755);
    wire[0:0] s8768, in8768_1, in8768_2;
    wire c8768;
    assign in8768_1 = {c5759};
    assign in8768_2 = {c5760};
    Full_Adder FA_8768(s8768, c8768, in8768_1, in8768_2, c5758);
    wire[0:0] s8769, in8769_1, in8769_2;
    wire c8769;
    assign in8769_1 = {c5762};
    assign in8769_2 = {c5763};
    Full_Adder FA_8769(s8769, c8769, in8769_1, in8769_2, c5761);
    wire[0:0] s8770, in8770_1, in8770_2;
    wire c8770;
    assign in8770_1 = {c5765};
    assign in8770_2 = {c5766};
    Full_Adder FA_8770(s8770, c8770, in8770_1, in8770_2, c5764);
    wire[0:0] s8771, in8771_1, in8771_2;
    wire c8771;
    assign in8771_1 = {c5768};
    assign in8771_2 = {s5769[0]};
    Full_Adder FA_8771(s8771, c8771, in8771_1, in8771_2, c5767);
    wire[0:0] s8772, in8772_1, in8772_2;
    wire c8772;
    assign in8772_1 = {s5771[0]};
    assign in8772_2 = {s5772[0]};
    Full_Adder FA_8772(s8772, c8772, in8772_1, in8772_2, s5770[0]);
    wire[0:0] s8773, in8773_1, in8773_2;
    wire c8773;
    assign in8773_1 = {s5774[0]};
    assign in8773_2 = {s5775[0]};
    Full_Adder FA_8773(s8773, c8773, in8773_1, in8773_2, s5773[0]);
    wire[0:0] s8774, in8774_1, in8774_2;
    wire c8774;
    assign in8774_1 = {s5777[0]};
    assign in8774_2 = {s5778[0]};
    Full_Adder FA_8774(s8774, c8774, in8774_1, in8774_2, s5776[0]);
    wire[0:0] s8775, in8775_1, in8775_2;
    wire c8775;
    assign in8775_1 = {s5780[0]};
    assign in8775_2 = {s5781[0]};
    Full_Adder FA_8775(s8775, c8775, in8775_1, in8775_2, s5779[0]);
    wire[0:0] s8776, in8776_1, in8776_2;
    wire c8776;
    assign in8776_1 = {s5783[0]};
    assign in8776_2 = {s5784[0]};
    Full_Adder FA_8776(s8776, c8776, in8776_1, in8776_2, s5782[0]);
    wire[0:0] s8777, in8777_1, in8777_2;
    wire c8777;
    assign in8777_1 = {s5786[0]};
    assign in8777_2 = {s5787[0]};
    Full_Adder FA_8777(s8777, c8777, in8777_1, in8777_2, s5785[0]);
    wire[0:0] s8778, in8778_1, in8778_2;
    wire c8778;
    assign in8778_1 = {c5769};
    assign in8778_2 = {c5770};
    Full_Adder FA_8778(s8778, c8778, in8778_1, in8778_2, s2380[0]);
    wire[0:0] s8779, in8779_1, in8779_2;
    wire c8779;
    assign in8779_1 = {c5772};
    assign in8779_2 = {c5773};
    Full_Adder FA_8779(s8779, c8779, in8779_1, in8779_2, c5771);
    wire[0:0] s8780, in8780_1, in8780_2;
    wire c8780;
    assign in8780_1 = {c5775};
    assign in8780_2 = {c5776};
    Full_Adder FA_8780(s8780, c8780, in8780_1, in8780_2, c5774);
    wire[0:0] s8781, in8781_1, in8781_2;
    wire c8781;
    assign in8781_1 = {c5778};
    assign in8781_2 = {c5779};
    Full_Adder FA_8781(s8781, c8781, in8781_1, in8781_2, c5777);
    wire[0:0] s8782, in8782_1, in8782_2;
    wire c8782;
    assign in8782_1 = {c5781};
    assign in8782_2 = {c5782};
    Full_Adder FA_8782(s8782, c8782, in8782_1, in8782_2, c5780);
    wire[0:0] s8783, in8783_1, in8783_2;
    wire c8783;
    assign in8783_1 = {c5784};
    assign in8783_2 = {c5785};
    Full_Adder FA_8783(s8783, c8783, in8783_1, in8783_2, c5783);
    wire[0:0] s8784, in8784_1, in8784_2;
    wire c8784;
    assign in8784_1 = {c5787};
    assign in8784_2 = {s5788[0]};
    Full_Adder FA_8784(s8784, c8784, in8784_1, in8784_2, c5786);
    wire[0:0] s8785, in8785_1, in8785_2;
    wire c8785;
    assign in8785_1 = {s5790[0]};
    assign in8785_2 = {s5791[0]};
    Full_Adder FA_8785(s8785, c8785, in8785_1, in8785_2, s5789[0]);
    wire[0:0] s8786, in8786_1, in8786_2;
    wire c8786;
    assign in8786_1 = {s5793[0]};
    assign in8786_2 = {s5794[0]};
    Full_Adder FA_8786(s8786, c8786, in8786_1, in8786_2, s5792[0]);
    wire[0:0] s8787, in8787_1, in8787_2;
    wire c8787;
    assign in8787_1 = {s5796[0]};
    assign in8787_2 = {s5797[0]};
    Full_Adder FA_8787(s8787, c8787, in8787_1, in8787_2, s5795[0]);
    wire[0:0] s8788, in8788_1, in8788_2;
    wire c8788;
    assign in8788_1 = {s5799[0]};
    assign in8788_2 = {s5800[0]};
    Full_Adder FA_8788(s8788, c8788, in8788_1, in8788_2, s5798[0]);
    wire[0:0] s8789, in8789_1, in8789_2;
    wire c8789;
    assign in8789_1 = {s5802[0]};
    assign in8789_2 = {s5803[0]};
    Full_Adder FA_8789(s8789, c8789, in8789_1, in8789_2, s5801[0]);
    wire[0:0] s8790, in8790_1, in8790_2;
    wire c8790;
    assign in8790_1 = {s5805[0]};
    assign in8790_2 = {s5806[0]};
    Full_Adder FA_8790(s8790, c8790, in8790_1, in8790_2, s5804[0]);
    wire[0:0] s8791, in8791_1, in8791_2;
    wire c8791;
    assign in8791_1 = {c5788};
    assign in8791_2 = {c5789};
    Full_Adder FA_8791(s8791, c8791, in8791_1, in8791_2, s2408[0]);
    wire[0:0] s8792, in8792_1, in8792_2;
    wire c8792;
    assign in8792_1 = {c5791};
    assign in8792_2 = {c5792};
    Full_Adder FA_8792(s8792, c8792, in8792_1, in8792_2, c5790);
    wire[0:0] s8793, in8793_1, in8793_2;
    wire c8793;
    assign in8793_1 = {c5794};
    assign in8793_2 = {c5795};
    Full_Adder FA_8793(s8793, c8793, in8793_1, in8793_2, c5793);
    wire[0:0] s8794, in8794_1, in8794_2;
    wire c8794;
    assign in8794_1 = {c5797};
    assign in8794_2 = {c5798};
    Full_Adder FA_8794(s8794, c8794, in8794_1, in8794_2, c5796);
    wire[0:0] s8795, in8795_1, in8795_2;
    wire c8795;
    assign in8795_1 = {c5800};
    assign in8795_2 = {c5801};
    Full_Adder FA_8795(s8795, c8795, in8795_1, in8795_2, c5799);
    wire[0:0] s8796, in8796_1, in8796_2;
    wire c8796;
    assign in8796_1 = {c5803};
    assign in8796_2 = {c5804};
    Full_Adder FA_8796(s8796, c8796, in8796_1, in8796_2, c5802);
    wire[0:0] s8797, in8797_1, in8797_2;
    wire c8797;
    assign in8797_1 = {c5806};
    assign in8797_2 = {s5807[0]};
    Full_Adder FA_8797(s8797, c8797, in8797_1, in8797_2, c5805);
    wire[0:0] s8798, in8798_1, in8798_2;
    wire c8798;
    assign in8798_1 = {s5809[0]};
    assign in8798_2 = {s5810[0]};
    Full_Adder FA_8798(s8798, c8798, in8798_1, in8798_2, s5808[0]);
    wire[0:0] s8799, in8799_1, in8799_2;
    wire c8799;
    assign in8799_1 = {s5812[0]};
    assign in8799_2 = {s5813[0]};
    Full_Adder FA_8799(s8799, c8799, in8799_1, in8799_2, s5811[0]);
    wire[0:0] s8800, in8800_1, in8800_2;
    wire c8800;
    assign in8800_1 = {s5815[0]};
    assign in8800_2 = {s5816[0]};
    Full_Adder FA_8800(s8800, c8800, in8800_1, in8800_2, s5814[0]);
    wire[0:0] s8801, in8801_1, in8801_2;
    wire c8801;
    assign in8801_1 = {s5818[0]};
    assign in8801_2 = {s5819[0]};
    Full_Adder FA_8801(s8801, c8801, in8801_1, in8801_2, s5817[0]);
    wire[0:0] s8802, in8802_1, in8802_2;
    wire c8802;
    assign in8802_1 = {s5821[0]};
    assign in8802_2 = {s5822[0]};
    Full_Adder FA_8802(s8802, c8802, in8802_1, in8802_2, s5820[0]);
    wire[0:0] s8803, in8803_1, in8803_2;
    wire c8803;
    assign in8803_1 = {s5824[0]};
    assign in8803_2 = {s5825[0]};
    Full_Adder FA_8803(s8803, c8803, in8803_1, in8803_2, s5823[0]);
    wire[0:0] s8804, in8804_1, in8804_2;
    wire c8804;
    assign in8804_1 = {c5807};
    assign in8804_2 = {c5808};
    Full_Adder FA_8804(s8804, c8804, in8804_1, in8804_2, s2436[0]);
    wire[0:0] s8805, in8805_1, in8805_2;
    wire c8805;
    assign in8805_1 = {c5810};
    assign in8805_2 = {c5811};
    Full_Adder FA_8805(s8805, c8805, in8805_1, in8805_2, c5809);
    wire[0:0] s8806, in8806_1, in8806_2;
    wire c8806;
    assign in8806_1 = {c5813};
    assign in8806_2 = {c5814};
    Full_Adder FA_8806(s8806, c8806, in8806_1, in8806_2, c5812);
    wire[0:0] s8807, in8807_1, in8807_2;
    wire c8807;
    assign in8807_1 = {c5816};
    assign in8807_2 = {c5817};
    Full_Adder FA_8807(s8807, c8807, in8807_1, in8807_2, c5815);
    wire[0:0] s8808, in8808_1, in8808_2;
    wire c8808;
    assign in8808_1 = {c5819};
    assign in8808_2 = {c5820};
    Full_Adder FA_8808(s8808, c8808, in8808_1, in8808_2, c5818);
    wire[0:0] s8809, in8809_1, in8809_2;
    wire c8809;
    assign in8809_1 = {c5822};
    assign in8809_2 = {c5823};
    Full_Adder FA_8809(s8809, c8809, in8809_1, in8809_2, c5821);
    wire[0:0] s8810, in8810_1, in8810_2;
    wire c8810;
    assign in8810_1 = {c5825};
    assign in8810_2 = {s5826[0]};
    Full_Adder FA_8810(s8810, c8810, in8810_1, in8810_2, c5824);
    wire[0:0] s8811, in8811_1, in8811_2;
    wire c8811;
    assign in8811_1 = {s5828[0]};
    assign in8811_2 = {s5829[0]};
    Full_Adder FA_8811(s8811, c8811, in8811_1, in8811_2, s5827[0]);
    wire[0:0] s8812, in8812_1, in8812_2;
    wire c8812;
    assign in8812_1 = {s5831[0]};
    assign in8812_2 = {s5832[0]};
    Full_Adder FA_8812(s8812, c8812, in8812_1, in8812_2, s5830[0]);
    wire[0:0] s8813, in8813_1, in8813_2;
    wire c8813;
    assign in8813_1 = {s5834[0]};
    assign in8813_2 = {s5835[0]};
    Full_Adder FA_8813(s8813, c8813, in8813_1, in8813_2, s5833[0]);
    wire[0:0] s8814, in8814_1, in8814_2;
    wire c8814;
    assign in8814_1 = {s5837[0]};
    assign in8814_2 = {s5838[0]};
    Full_Adder FA_8814(s8814, c8814, in8814_1, in8814_2, s5836[0]);
    wire[0:0] s8815, in8815_1, in8815_2;
    wire c8815;
    assign in8815_1 = {s5840[0]};
    assign in8815_2 = {s5841[0]};
    Full_Adder FA_8815(s8815, c8815, in8815_1, in8815_2, s5839[0]);
    wire[0:0] s8816, in8816_1, in8816_2;
    wire c8816;
    assign in8816_1 = {s5843[0]};
    assign in8816_2 = {s5844[0]};
    Full_Adder FA_8816(s8816, c8816, in8816_1, in8816_2, s5842[0]);
    wire[0:0] s8817, in8817_1, in8817_2;
    wire c8817;
    assign in8817_1 = {c5826};
    assign in8817_2 = {c5827};
    Full_Adder FA_8817(s8817, c8817, in8817_1, in8817_2, s2464[0]);
    wire[0:0] s8818, in8818_1, in8818_2;
    wire c8818;
    assign in8818_1 = {c5829};
    assign in8818_2 = {c5830};
    Full_Adder FA_8818(s8818, c8818, in8818_1, in8818_2, c5828);
    wire[0:0] s8819, in8819_1, in8819_2;
    wire c8819;
    assign in8819_1 = {c5832};
    assign in8819_2 = {c5833};
    Full_Adder FA_8819(s8819, c8819, in8819_1, in8819_2, c5831);
    wire[0:0] s8820, in8820_1, in8820_2;
    wire c8820;
    assign in8820_1 = {c5835};
    assign in8820_2 = {c5836};
    Full_Adder FA_8820(s8820, c8820, in8820_1, in8820_2, c5834);
    wire[0:0] s8821, in8821_1, in8821_2;
    wire c8821;
    assign in8821_1 = {c5838};
    assign in8821_2 = {c5839};
    Full_Adder FA_8821(s8821, c8821, in8821_1, in8821_2, c5837);
    wire[0:0] s8822, in8822_1, in8822_2;
    wire c8822;
    assign in8822_1 = {c5841};
    assign in8822_2 = {c5842};
    Full_Adder FA_8822(s8822, c8822, in8822_1, in8822_2, c5840);
    wire[0:0] s8823, in8823_1, in8823_2;
    wire c8823;
    assign in8823_1 = {c5844};
    assign in8823_2 = {s5845[0]};
    Full_Adder FA_8823(s8823, c8823, in8823_1, in8823_2, c5843);
    wire[0:0] s8824, in8824_1, in8824_2;
    wire c8824;
    assign in8824_1 = {s5847[0]};
    assign in8824_2 = {s5848[0]};
    Full_Adder FA_8824(s8824, c8824, in8824_1, in8824_2, s5846[0]);
    wire[0:0] s8825, in8825_1, in8825_2;
    wire c8825;
    assign in8825_1 = {s5850[0]};
    assign in8825_2 = {s5851[0]};
    Full_Adder FA_8825(s8825, c8825, in8825_1, in8825_2, s5849[0]);
    wire[0:0] s8826, in8826_1, in8826_2;
    wire c8826;
    assign in8826_1 = {s5853[0]};
    assign in8826_2 = {s5854[0]};
    Full_Adder FA_8826(s8826, c8826, in8826_1, in8826_2, s5852[0]);
    wire[0:0] s8827, in8827_1, in8827_2;
    wire c8827;
    assign in8827_1 = {s5856[0]};
    assign in8827_2 = {s5857[0]};
    Full_Adder FA_8827(s8827, c8827, in8827_1, in8827_2, s5855[0]);
    wire[0:0] s8828, in8828_1, in8828_2;
    wire c8828;
    assign in8828_1 = {s5859[0]};
    assign in8828_2 = {s5860[0]};
    Full_Adder FA_8828(s8828, c8828, in8828_1, in8828_2, s5858[0]);
    wire[0:0] s8829, in8829_1, in8829_2;
    wire c8829;
    assign in8829_1 = {s5862[0]};
    assign in8829_2 = {s5863[0]};
    Full_Adder FA_8829(s8829, c8829, in8829_1, in8829_2, s5861[0]);
    wire[0:0] s8830, in8830_1, in8830_2;
    wire c8830;
    assign in8830_1 = {c5845};
    assign in8830_2 = {c5846};
    Full_Adder FA_8830(s8830, c8830, in8830_1, in8830_2, s2492[0]);
    wire[0:0] s8831, in8831_1, in8831_2;
    wire c8831;
    assign in8831_1 = {c5848};
    assign in8831_2 = {c5849};
    Full_Adder FA_8831(s8831, c8831, in8831_1, in8831_2, c5847);
    wire[0:0] s8832, in8832_1, in8832_2;
    wire c8832;
    assign in8832_1 = {c5851};
    assign in8832_2 = {c5852};
    Full_Adder FA_8832(s8832, c8832, in8832_1, in8832_2, c5850);
    wire[0:0] s8833, in8833_1, in8833_2;
    wire c8833;
    assign in8833_1 = {c5854};
    assign in8833_2 = {c5855};
    Full_Adder FA_8833(s8833, c8833, in8833_1, in8833_2, c5853);
    wire[0:0] s8834, in8834_1, in8834_2;
    wire c8834;
    assign in8834_1 = {c5857};
    assign in8834_2 = {c5858};
    Full_Adder FA_8834(s8834, c8834, in8834_1, in8834_2, c5856);
    wire[0:0] s8835, in8835_1, in8835_2;
    wire c8835;
    assign in8835_1 = {c5860};
    assign in8835_2 = {c5861};
    Full_Adder FA_8835(s8835, c8835, in8835_1, in8835_2, c5859);
    wire[0:0] s8836, in8836_1, in8836_2;
    wire c8836;
    assign in8836_1 = {c5863};
    assign in8836_2 = {s5864[0]};
    Full_Adder FA_8836(s8836, c8836, in8836_1, in8836_2, c5862);
    wire[0:0] s8837, in8837_1, in8837_2;
    wire c8837;
    assign in8837_1 = {s5866[0]};
    assign in8837_2 = {s5867[0]};
    Full_Adder FA_8837(s8837, c8837, in8837_1, in8837_2, s5865[0]);
    wire[0:0] s8838, in8838_1, in8838_2;
    wire c8838;
    assign in8838_1 = {s5869[0]};
    assign in8838_2 = {s5870[0]};
    Full_Adder FA_8838(s8838, c8838, in8838_1, in8838_2, s5868[0]);
    wire[0:0] s8839, in8839_1, in8839_2;
    wire c8839;
    assign in8839_1 = {s5872[0]};
    assign in8839_2 = {s5873[0]};
    Full_Adder FA_8839(s8839, c8839, in8839_1, in8839_2, s5871[0]);
    wire[0:0] s8840, in8840_1, in8840_2;
    wire c8840;
    assign in8840_1 = {s5875[0]};
    assign in8840_2 = {s5876[0]};
    Full_Adder FA_8840(s8840, c8840, in8840_1, in8840_2, s5874[0]);
    wire[0:0] s8841, in8841_1, in8841_2;
    wire c8841;
    assign in8841_1 = {s5878[0]};
    assign in8841_2 = {s5879[0]};
    Full_Adder FA_8841(s8841, c8841, in8841_1, in8841_2, s5877[0]);
    wire[0:0] s8842, in8842_1, in8842_2;
    wire c8842;
    assign in8842_1 = {s5881[0]};
    assign in8842_2 = {s5882[0]};
    Full_Adder FA_8842(s8842, c8842, in8842_1, in8842_2, s5880[0]);
    wire[0:0] s8843, in8843_1, in8843_2;
    wire c8843;
    assign in8843_1 = {c5864};
    assign in8843_2 = {c5865};
    Full_Adder FA_8843(s8843, c8843, in8843_1, in8843_2, s2520[0]);
    wire[0:0] s8844, in8844_1, in8844_2;
    wire c8844;
    assign in8844_1 = {c5867};
    assign in8844_2 = {c5868};
    Full_Adder FA_8844(s8844, c8844, in8844_1, in8844_2, c5866);
    wire[0:0] s8845, in8845_1, in8845_2;
    wire c8845;
    assign in8845_1 = {c5870};
    assign in8845_2 = {c5871};
    Full_Adder FA_8845(s8845, c8845, in8845_1, in8845_2, c5869);
    wire[0:0] s8846, in8846_1, in8846_2;
    wire c8846;
    assign in8846_1 = {c5873};
    assign in8846_2 = {c5874};
    Full_Adder FA_8846(s8846, c8846, in8846_1, in8846_2, c5872);
    wire[0:0] s8847, in8847_1, in8847_2;
    wire c8847;
    assign in8847_1 = {c5876};
    assign in8847_2 = {c5877};
    Full_Adder FA_8847(s8847, c8847, in8847_1, in8847_2, c5875);
    wire[0:0] s8848, in8848_1, in8848_2;
    wire c8848;
    assign in8848_1 = {c5879};
    assign in8848_2 = {c5880};
    Full_Adder FA_8848(s8848, c8848, in8848_1, in8848_2, c5878);
    wire[0:0] s8849, in8849_1, in8849_2;
    wire c8849;
    assign in8849_1 = {c5882};
    assign in8849_2 = {s5883[0]};
    Full_Adder FA_8849(s8849, c8849, in8849_1, in8849_2, c5881);
    wire[0:0] s8850, in8850_1, in8850_2;
    wire c8850;
    assign in8850_1 = {s5885[0]};
    assign in8850_2 = {s5886[0]};
    Full_Adder FA_8850(s8850, c8850, in8850_1, in8850_2, s5884[0]);
    wire[0:0] s8851, in8851_1, in8851_2;
    wire c8851;
    assign in8851_1 = {s5888[0]};
    assign in8851_2 = {s5889[0]};
    Full_Adder FA_8851(s8851, c8851, in8851_1, in8851_2, s5887[0]);
    wire[0:0] s8852, in8852_1, in8852_2;
    wire c8852;
    assign in8852_1 = {s5891[0]};
    assign in8852_2 = {s5892[0]};
    Full_Adder FA_8852(s8852, c8852, in8852_1, in8852_2, s5890[0]);
    wire[0:0] s8853, in8853_1, in8853_2;
    wire c8853;
    assign in8853_1 = {s5894[0]};
    assign in8853_2 = {s5895[0]};
    Full_Adder FA_8853(s8853, c8853, in8853_1, in8853_2, s5893[0]);
    wire[0:0] s8854, in8854_1, in8854_2;
    wire c8854;
    assign in8854_1 = {s5897[0]};
    assign in8854_2 = {s5898[0]};
    Full_Adder FA_8854(s8854, c8854, in8854_1, in8854_2, s5896[0]);
    wire[0:0] s8855, in8855_1, in8855_2;
    wire c8855;
    assign in8855_1 = {s5900[0]};
    assign in8855_2 = {s5901[0]};
    Full_Adder FA_8855(s8855, c8855, in8855_1, in8855_2, s5899[0]);
    wire[0:0] s8856, in8856_1, in8856_2;
    wire c8856;
    assign in8856_1 = {c5883};
    assign in8856_2 = {c5884};
    Full_Adder FA_8856(s8856, c8856, in8856_1, in8856_2, s2548[0]);
    wire[0:0] s8857, in8857_1, in8857_2;
    wire c8857;
    assign in8857_1 = {c5886};
    assign in8857_2 = {c5887};
    Full_Adder FA_8857(s8857, c8857, in8857_1, in8857_2, c5885);
    wire[0:0] s8858, in8858_1, in8858_2;
    wire c8858;
    assign in8858_1 = {c5889};
    assign in8858_2 = {c5890};
    Full_Adder FA_8858(s8858, c8858, in8858_1, in8858_2, c5888);
    wire[0:0] s8859, in8859_1, in8859_2;
    wire c8859;
    assign in8859_1 = {c5892};
    assign in8859_2 = {c5893};
    Full_Adder FA_8859(s8859, c8859, in8859_1, in8859_2, c5891);
    wire[0:0] s8860, in8860_1, in8860_2;
    wire c8860;
    assign in8860_1 = {c5895};
    assign in8860_2 = {c5896};
    Full_Adder FA_8860(s8860, c8860, in8860_1, in8860_2, c5894);
    wire[0:0] s8861, in8861_1, in8861_2;
    wire c8861;
    assign in8861_1 = {c5898};
    assign in8861_2 = {c5899};
    Full_Adder FA_8861(s8861, c8861, in8861_1, in8861_2, c5897);
    wire[0:0] s8862, in8862_1, in8862_2;
    wire c8862;
    assign in8862_1 = {c5901};
    assign in8862_2 = {s5902[0]};
    Full_Adder FA_8862(s8862, c8862, in8862_1, in8862_2, c5900);
    wire[0:0] s8863, in8863_1, in8863_2;
    wire c8863;
    assign in8863_1 = {s5904[0]};
    assign in8863_2 = {s5905[0]};
    Full_Adder FA_8863(s8863, c8863, in8863_1, in8863_2, s5903[0]);
    wire[0:0] s8864, in8864_1, in8864_2;
    wire c8864;
    assign in8864_1 = {s5907[0]};
    assign in8864_2 = {s5908[0]};
    Full_Adder FA_8864(s8864, c8864, in8864_1, in8864_2, s5906[0]);
    wire[0:0] s8865, in8865_1, in8865_2;
    wire c8865;
    assign in8865_1 = {s5910[0]};
    assign in8865_2 = {s5911[0]};
    Full_Adder FA_8865(s8865, c8865, in8865_1, in8865_2, s5909[0]);
    wire[0:0] s8866, in8866_1, in8866_2;
    wire c8866;
    assign in8866_1 = {s5913[0]};
    assign in8866_2 = {s5914[0]};
    Full_Adder FA_8866(s8866, c8866, in8866_1, in8866_2, s5912[0]);
    wire[0:0] s8867, in8867_1, in8867_2;
    wire c8867;
    assign in8867_1 = {s5916[0]};
    assign in8867_2 = {s5917[0]};
    Full_Adder FA_8867(s8867, c8867, in8867_1, in8867_2, s5915[0]);
    wire[0:0] s8868, in8868_1, in8868_2;
    wire c8868;
    assign in8868_1 = {s5919[0]};
    assign in8868_2 = {s5920[0]};
    Full_Adder FA_8868(s8868, c8868, in8868_1, in8868_2, s5918[0]);
    wire[0:0] s8869, in8869_1, in8869_2;
    wire c8869;
    assign in8869_1 = {c5902};
    assign in8869_2 = {c5903};
    Full_Adder FA_8869(s8869, c8869, in8869_1, in8869_2, s2576[0]);
    wire[0:0] s8870, in8870_1, in8870_2;
    wire c8870;
    assign in8870_1 = {c5905};
    assign in8870_2 = {c5906};
    Full_Adder FA_8870(s8870, c8870, in8870_1, in8870_2, c5904);
    wire[0:0] s8871, in8871_1, in8871_2;
    wire c8871;
    assign in8871_1 = {c5908};
    assign in8871_2 = {c5909};
    Full_Adder FA_8871(s8871, c8871, in8871_1, in8871_2, c5907);
    wire[0:0] s8872, in8872_1, in8872_2;
    wire c8872;
    assign in8872_1 = {c5911};
    assign in8872_2 = {c5912};
    Full_Adder FA_8872(s8872, c8872, in8872_1, in8872_2, c5910);
    wire[0:0] s8873, in8873_1, in8873_2;
    wire c8873;
    assign in8873_1 = {c5914};
    assign in8873_2 = {c5915};
    Full_Adder FA_8873(s8873, c8873, in8873_1, in8873_2, c5913);
    wire[0:0] s8874, in8874_1, in8874_2;
    wire c8874;
    assign in8874_1 = {c5917};
    assign in8874_2 = {c5918};
    Full_Adder FA_8874(s8874, c8874, in8874_1, in8874_2, c5916);
    wire[0:0] s8875, in8875_1, in8875_2;
    wire c8875;
    assign in8875_1 = {c5920};
    assign in8875_2 = {s5921[0]};
    Full_Adder FA_8875(s8875, c8875, in8875_1, in8875_2, c5919);
    wire[0:0] s8876, in8876_1, in8876_2;
    wire c8876;
    assign in8876_1 = {s5923[0]};
    assign in8876_2 = {s5924[0]};
    Full_Adder FA_8876(s8876, c8876, in8876_1, in8876_2, s5922[0]);
    wire[0:0] s8877, in8877_1, in8877_2;
    wire c8877;
    assign in8877_1 = {s5926[0]};
    assign in8877_2 = {s5927[0]};
    Full_Adder FA_8877(s8877, c8877, in8877_1, in8877_2, s5925[0]);
    wire[0:0] s8878, in8878_1, in8878_2;
    wire c8878;
    assign in8878_1 = {s5929[0]};
    assign in8878_2 = {s5930[0]};
    Full_Adder FA_8878(s8878, c8878, in8878_1, in8878_2, s5928[0]);
    wire[0:0] s8879, in8879_1, in8879_2;
    wire c8879;
    assign in8879_1 = {s5932[0]};
    assign in8879_2 = {s5933[0]};
    Full_Adder FA_8879(s8879, c8879, in8879_1, in8879_2, s5931[0]);
    wire[0:0] s8880, in8880_1, in8880_2;
    wire c8880;
    assign in8880_1 = {s5935[0]};
    assign in8880_2 = {s5936[0]};
    Full_Adder FA_8880(s8880, c8880, in8880_1, in8880_2, s5934[0]);
    wire[0:0] s8881, in8881_1, in8881_2;
    wire c8881;
    assign in8881_1 = {s5938[0]};
    assign in8881_2 = {s5939[0]};
    Full_Adder FA_8881(s8881, c8881, in8881_1, in8881_2, s5937[0]);
    wire[0:0] s8882, in8882_1, in8882_2;
    wire c8882;
    assign in8882_1 = {c5921};
    assign in8882_2 = {c5922};
    Full_Adder FA_8882(s8882, c8882, in8882_1, in8882_2, s2604[0]);
    wire[0:0] s8883, in8883_1, in8883_2;
    wire c8883;
    assign in8883_1 = {c5924};
    assign in8883_2 = {c5925};
    Full_Adder FA_8883(s8883, c8883, in8883_1, in8883_2, c5923);
    wire[0:0] s8884, in8884_1, in8884_2;
    wire c8884;
    assign in8884_1 = {c5927};
    assign in8884_2 = {c5928};
    Full_Adder FA_8884(s8884, c8884, in8884_1, in8884_2, c5926);
    wire[0:0] s8885, in8885_1, in8885_2;
    wire c8885;
    assign in8885_1 = {c5930};
    assign in8885_2 = {c5931};
    Full_Adder FA_8885(s8885, c8885, in8885_1, in8885_2, c5929);
    wire[0:0] s8886, in8886_1, in8886_2;
    wire c8886;
    assign in8886_1 = {c5933};
    assign in8886_2 = {c5934};
    Full_Adder FA_8886(s8886, c8886, in8886_1, in8886_2, c5932);
    wire[0:0] s8887, in8887_1, in8887_2;
    wire c8887;
    assign in8887_1 = {c5936};
    assign in8887_2 = {c5937};
    Full_Adder FA_8887(s8887, c8887, in8887_1, in8887_2, c5935);
    wire[0:0] s8888, in8888_1, in8888_2;
    wire c8888;
    assign in8888_1 = {c5939};
    assign in8888_2 = {s5940[0]};
    Full_Adder FA_8888(s8888, c8888, in8888_1, in8888_2, c5938);
    wire[0:0] s8889, in8889_1, in8889_2;
    wire c8889;
    assign in8889_1 = {s5942[0]};
    assign in8889_2 = {s5943[0]};
    Full_Adder FA_8889(s8889, c8889, in8889_1, in8889_2, s5941[0]);
    wire[0:0] s8890, in8890_1, in8890_2;
    wire c8890;
    assign in8890_1 = {s5945[0]};
    assign in8890_2 = {s5946[0]};
    Full_Adder FA_8890(s8890, c8890, in8890_1, in8890_2, s5944[0]);
    wire[0:0] s8891, in8891_1, in8891_2;
    wire c8891;
    assign in8891_1 = {s5948[0]};
    assign in8891_2 = {s5949[0]};
    Full_Adder FA_8891(s8891, c8891, in8891_1, in8891_2, s5947[0]);
    wire[0:0] s8892, in8892_1, in8892_2;
    wire c8892;
    assign in8892_1 = {s5951[0]};
    assign in8892_2 = {s5952[0]};
    Full_Adder FA_8892(s8892, c8892, in8892_1, in8892_2, s5950[0]);
    wire[0:0] s8893, in8893_1, in8893_2;
    wire c8893;
    assign in8893_1 = {s5954[0]};
    assign in8893_2 = {s5955[0]};
    Full_Adder FA_8893(s8893, c8893, in8893_1, in8893_2, s5953[0]);
    wire[0:0] s8894, in8894_1, in8894_2;
    wire c8894;
    assign in8894_1 = {s5957[0]};
    assign in8894_2 = {s5958[0]};
    Full_Adder FA_8894(s8894, c8894, in8894_1, in8894_2, s5956[0]);
    wire[0:0] s8895, in8895_1, in8895_2;
    wire c8895;
    assign in8895_1 = {c5940};
    assign in8895_2 = {c5941};
    Full_Adder FA_8895(s8895, c8895, in8895_1, in8895_2, s2632[0]);
    wire[0:0] s8896, in8896_1, in8896_2;
    wire c8896;
    assign in8896_1 = {c5943};
    assign in8896_2 = {c5944};
    Full_Adder FA_8896(s8896, c8896, in8896_1, in8896_2, c5942);
    wire[0:0] s8897, in8897_1, in8897_2;
    wire c8897;
    assign in8897_1 = {c5946};
    assign in8897_2 = {c5947};
    Full_Adder FA_8897(s8897, c8897, in8897_1, in8897_2, c5945);
    wire[0:0] s8898, in8898_1, in8898_2;
    wire c8898;
    assign in8898_1 = {c5949};
    assign in8898_2 = {c5950};
    Full_Adder FA_8898(s8898, c8898, in8898_1, in8898_2, c5948);
    wire[0:0] s8899, in8899_1, in8899_2;
    wire c8899;
    assign in8899_1 = {c5952};
    assign in8899_2 = {c5953};
    Full_Adder FA_8899(s8899, c8899, in8899_1, in8899_2, c5951);
    wire[0:0] s8900, in8900_1, in8900_2;
    wire c8900;
    assign in8900_1 = {c5955};
    assign in8900_2 = {c5956};
    Full_Adder FA_8900(s8900, c8900, in8900_1, in8900_2, c5954);
    wire[0:0] s8901, in8901_1, in8901_2;
    wire c8901;
    assign in8901_1 = {c5958};
    assign in8901_2 = {s5959[0]};
    Full_Adder FA_8901(s8901, c8901, in8901_1, in8901_2, c5957);
    wire[0:0] s8902, in8902_1, in8902_2;
    wire c8902;
    assign in8902_1 = {s5961[0]};
    assign in8902_2 = {s5962[0]};
    Full_Adder FA_8902(s8902, c8902, in8902_1, in8902_2, s5960[0]);
    wire[0:0] s8903, in8903_1, in8903_2;
    wire c8903;
    assign in8903_1 = {s5964[0]};
    assign in8903_2 = {s5965[0]};
    Full_Adder FA_8903(s8903, c8903, in8903_1, in8903_2, s5963[0]);
    wire[0:0] s8904, in8904_1, in8904_2;
    wire c8904;
    assign in8904_1 = {s5967[0]};
    assign in8904_2 = {s5968[0]};
    Full_Adder FA_8904(s8904, c8904, in8904_1, in8904_2, s5966[0]);
    wire[0:0] s8905, in8905_1, in8905_2;
    wire c8905;
    assign in8905_1 = {s5970[0]};
    assign in8905_2 = {s5971[0]};
    Full_Adder FA_8905(s8905, c8905, in8905_1, in8905_2, s5969[0]);
    wire[0:0] s8906, in8906_1, in8906_2;
    wire c8906;
    assign in8906_1 = {s5973[0]};
    assign in8906_2 = {s5974[0]};
    Full_Adder FA_8906(s8906, c8906, in8906_1, in8906_2, s5972[0]);
    wire[0:0] s8907, in8907_1, in8907_2;
    wire c8907;
    assign in8907_1 = {s5976[0]};
    assign in8907_2 = {s5977[0]};
    Full_Adder FA_8907(s8907, c8907, in8907_1, in8907_2, s5975[0]);
    wire[0:0] s8908, in8908_1, in8908_2;
    wire c8908;
    assign in8908_1 = {c5959};
    assign in8908_2 = {c5960};
    Full_Adder FA_8908(s8908, c8908, in8908_1, in8908_2, s2660[0]);
    wire[0:0] s8909, in8909_1, in8909_2;
    wire c8909;
    assign in8909_1 = {c5962};
    assign in8909_2 = {c5963};
    Full_Adder FA_8909(s8909, c8909, in8909_1, in8909_2, c5961);
    wire[0:0] s8910, in8910_1, in8910_2;
    wire c8910;
    assign in8910_1 = {c5965};
    assign in8910_2 = {c5966};
    Full_Adder FA_8910(s8910, c8910, in8910_1, in8910_2, c5964);
    wire[0:0] s8911, in8911_1, in8911_2;
    wire c8911;
    assign in8911_1 = {c5968};
    assign in8911_2 = {c5969};
    Full_Adder FA_8911(s8911, c8911, in8911_1, in8911_2, c5967);
    wire[0:0] s8912, in8912_1, in8912_2;
    wire c8912;
    assign in8912_1 = {c5971};
    assign in8912_2 = {c5972};
    Full_Adder FA_8912(s8912, c8912, in8912_1, in8912_2, c5970);
    wire[0:0] s8913, in8913_1, in8913_2;
    wire c8913;
    assign in8913_1 = {c5974};
    assign in8913_2 = {c5975};
    Full_Adder FA_8913(s8913, c8913, in8913_1, in8913_2, c5973);
    wire[0:0] s8914, in8914_1, in8914_2;
    wire c8914;
    assign in8914_1 = {c5977};
    assign in8914_2 = {s5978[0]};
    Full_Adder FA_8914(s8914, c8914, in8914_1, in8914_2, c5976);
    wire[0:0] s8915, in8915_1, in8915_2;
    wire c8915;
    assign in8915_1 = {s5980[0]};
    assign in8915_2 = {s5981[0]};
    Full_Adder FA_8915(s8915, c8915, in8915_1, in8915_2, s5979[0]);
    wire[0:0] s8916, in8916_1, in8916_2;
    wire c8916;
    assign in8916_1 = {s5983[0]};
    assign in8916_2 = {s5984[0]};
    Full_Adder FA_8916(s8916, c8916, in8916_1, in8916_2, s5982[0]);
    wire[0:0] s8917, in8917_1, in8917_2;
    wire c8917;
    assign in8917_1 = {s5986[0]};
    assign in8917_2 = {s5987[0]};
    Full_Adder FA_8917(s8917, c8917, in8917_1, in8917_2, s5985[0]);
    wire[0:0] s8918, in8918_1, in8918_2;
    wire c8918;
    assign in8918_1 = {s5989[0]};
    assign in8918_2 = {s5990[0]};
    Full_Adder FA_8918(s8918, c8918, in8918_1, in8918_2, s5988[0]);
    wire[0:0] s8919, in8919_1, in8919_2;
    wire c8919;
    assign in8919_1 = {s5992[0]};
    assign in8919_2 = {s5993[0]};
    Full_Adder FA_8919(s8919, c8919, in8919_1, in8919_2, s5991[0]);
    wire[0:0] s8920, in8920_1, in8920_2;
    wire c8920;
    assign in8920_1 = {s5995[0]};
    assign in8920_2 = {s5996[0]};
    Full_Adder FA_8920(s8920, c8920, in8920_1, in8920_2, s5994[0]);
    wire[0:0] s8921, in8921_1, in8921_2;
    wire c8921;
    assign in8921_1 = {c5978};
    assign in8921_2 = {c5979};
    Full_Adder FA_8921(s8921, c8921, in8921_1, in8921_2, s2688[0]);
    wire[0:0] s8922, in8922_1, in8922_2;
    wire c8922;
    assign in8922_1 = {c5981};
    assign in8922_2 = {c5982};
    Full_Adder FA_8922(s8922, c8922, in8922_1, in8922_2, c5980);
    wire[0:0] s8923, in8923_1, in8923_2;
    wire c8923;
    assign in8923_1 = {c5984};
    assign in8923_2 = {c5985};
    Full_Adder FA_8923(s8923, c8923, in8923_1, in8923_2, c5983);
    wire[0:0] s8924, in8924_1, in8924_2;
    wire c8924;
    assign in8924_1 = {c5987};
    assign in8924_2 = {c5988};
    Full_Adder FA_8924(s8924, c8924, in8924_1, in8924_2, c5986);
    wire[0:0] s8925, in8925_1, in8925_2;
    wire c8925;
    assign in8925_1 = {c5990};
    assign in8925_2 = {c5991};
    Full_Adder FA_8925(s8925, c8925, in8925_1, in8925_2, c5989);
    wire[0:0] s8926, in8926_1, in8926_2;
    wire c8926;
    assign in8926_1 = {c5993};
    assign in8926_2 = {c5994};
    Full_Adder FA_8926(s8926, c8926, in8926_1, in8926_2, c5992);
    wire[0:0] s8927, in8927_1, in8927_2;
    wire c8927;
    assign in8927_1 = {c5996};
    assign in8927_2 = {s5997[0]};
    Full_Adder FA_8927(s8927, c8927, in8927_1, in8927_2, c5995);
    wire[0:0] s8928, in8928_1, in8928_2;
    wire c8928;
    assign in8928_1 = {s5999[0]};
    assign in8928_2 = {s6000[0]};
    Full_Adder FA_8928(s8928, c8928, in8928_1, in8928_2, s5998[0]);
    wire[0:0] s8929, in8929_1, in8929_2;
    wire c8929;
    assign in8929_1 = {s6002[0]};
    assign in8929_2 = {s6003[0]};
    Full_Adder FA_8929(s8929, c8929, in8929_1, in8929_2, s6001[0]);
    wire[0:0] s8930, in8930_1, in8930_2;
    wire c8930;
    assign in8930_1 = {s6005[0]};
    assign in8930_2 = {s6006[0]};
    Full_Adder FA_8930(s8930, c8930, in8930_1, in8930_2, s6004[0]);
    wire[0:0] s8931, in8931_1, in8931_2;
    wire c8931;
    assign in8931_1 = {s6008[0]};
    assign in8931_2 = {s6009[0]};
    Full_Adder FA_8931(s8931, c8931, in8931_1, in8931_2, s6007[0]);
    wire[0:0] s8932, in8932_1, in8932_2;
    wire c8932;
    assign in8932_1 = {s6011[0]};
    assign in8932_2 = {s6012[0]};
    Full_Adder FA_8932(s8932, c8932, in8932_1, in8932_2, s6010[0]);
    wire[0:0] s8933, in8933_1, in8933_2;
    wire c8933;
    assign in8933_1 = {s6014[0]};
    assign in8933_2 = {s6015[0]};
    Full_Adder FA_8933(s8933, c8933, in8933_1, in8933_2, s6013[0]);
    wire[0:0] s8934, in8934_1, in8934_2;
    wire c8934;
    assign in8934_1 = {c5997};
    assign in8934_2 = {c5998};
    Full_Adder FA_8934(s8934, c8934, in8934_1, in8934_2, s2716[0]);
    wire[0:0] s8935, in8935_1, in8935_2;
    wire c8935;
    assign in8935_1 = {c6000};
    assign in8935_2 = {c6001};
    Full_Adder FA_8935(s8935, c8935, in8935_1, in8935_2, c5999);
    wire[0:0] s8936, in8936_1, in8936_2;
    wire c8936;
    assign in8936_1 = {c6003};
    assign in8936_2 = {c6004};
    Full_Adder FA_8936(s8936, c8936, in8936_1, in8936_2, c6002);
    wire[0:0] s8937, in8937_1, in8937_2;
    wire c8937;
    assign in8937_1 = {c6006};
    assign in8937_2 = {c6007};
    Full_Adder FA_8937(s8937, c8937, in8937_1, in8937_2, c6005);
    wire[0:0] s8938, in8938_1, in8938_2;
    wire c8938;
    assign in8938_1 = {c6009};
    assign in8938_2 = {c6010};
    Full_Adder FA_8938(s8938, c8938, in8938_1, in8938_2, c6008);
    wire[0:0] s8939, in8939_1, in8939_2;
    wire c8939;
    assign in8939_1 = {c6012};
    assign in8939_2 = {c6013};
    Full_Adder FA_8939(s8939, c8939, in8939_1, in8939_2, c6011);
    wire[0:0] s8940, in8940_1, in8940_2;
    wire c8940;
    assign in8940_1 = {c6015};
    assign in8940_2 = {s6016[0]};
    Full_Adder FA_8940(s8940, c8940, in8940_1, in8940_2, c6014);
    wire[0:0] s8941, in8941_1, in8941_2;
    wire c8941;
    assign in8941_1 = {s6018[0]};
    assign in8941_2 = {s6019[0]};
    Full_Adder FA_8941(s8941, c8941, in8941_1, in8941_2, s6017[0]);
    wire[0:0] s8942, in8942_1, in8942_2;
    wire c8942;
    assign in8942_1 = {s6021[0]};
    assign in8942_2 = {s6022[0]};
    Full_Adder FA_8942(s8942, c8942, in8942_1, in8942_2, s6020[0]);
    wire[0:0] s8943, in8943_1, in8943_2;
    wire c8943;
    assign in8943_1 = {s6024[0]};
    assign in8943_2 = {s6025[0]};
    Full_Adder FA_8943(s8943, c8943, in8943_1, in8943_2, s6023[0]);
    wire[0:0] s8944, in8944_1, in8944_2;
    wire c8944;
    assign in8944_1 = {s6027[0]};
    assign in8944_2 = {s6028[0]};
    Full_Adder FA_8944(s8944, c8944, in8944_1, in8944_2, s6026[0]);
    wire[0:0] s8945, in8945_1, in8945_2;
    wire c8945;
    assign in8945_1 = {s6030[0]};
    assign in8945_2 = {s6031[0]};
    Full_Adder FA_8945(s8945, c8945, in8945_1, in8945_2, s6029[0]);
    wire[0:0] s8946, in8946_1, in8946_2;
    wire c8946;
    assign in8946_1 = {s6033[0]};
    assign in8946_2 = {s6034[0]};
    Full_Adder FA_8946(s8946, c8946, in8946_1, in8946_2, s6032[0]);
    wire[0:0] s8947, in8947_1, in8947_2;
    wire c8947;
    assign in8947_1 = {c6016};
    assign in8947_2 = {c6017};
    Full_Adder FA_8947(s8947, c8947, in8947_1, in8947_2, s2744[0]);
    wire[0:0] s8948, in8948_1, in8948_2;
    wire c8948;
    assign in8948_1 = {c6019};
    assign in8948_2 = {c6020};
    Full_Adder FA_8948(s8948, c8948, in8948_1, in8948_2, c6018);
    wire[0:0] s8949, in8949_1, in8949_2;
    wire c8949;
    assign in8949_1 = {c6022};
    assign in8949_2 = {c6023};
    Full_Adder FA_8949(s8949, c8949, in8949_1, in8949_2, c6021);
    wire[0:0] s8950, in8950_1, in8950_2;
    wire c8950;
    assign in8950_1 = {c6025};
    assign in8950_2 = {c6026};
    Full_Adder FA_8950(s8950, c8950, in8950_1, in8950_2, c6024);
    wire[0:0] s8951, in8951_1, in8951_2;
    wire c8951;
    assign in8951_1 = {c6028};
    assign in8951_2 = {c6029};
    Full_Adder FA_8951(s8951, c8951, in8951_1, in8951_2, c6027);
    wire[0:0] s8952, in8952_1, in8952_2;
    wire c8952;
    assign in8952_1 = {c6031};
    assign in8952_2 = {c6032};
    Full_Adder FA_8952(s8952, c8952, in8952_1, in8952_2, c6030);
    wire[0:0] s8953, in8953_1, in8953_2;
    wire c8953;
    assign in8953_1 = {c6034};
    assign in8953_2 = {s6035[0]};
    Full_Adder FA_8953(s8953, c8953, in8953_1, in8953_2, c6033);
    wire[0:0] s8954, in8954_1, in8954_2;
    wire c8954;
    assign in8954_1 = {s6037[0]};
    assign in8954_2 = {s6038[0]};
    Full_Adder FA_8954(s8954, c8954, in8954_1, in8954_2, s6036[0]);
    wire[0:0] s8955, in8955_1, in8955_2;
    wire c8955;
    assign in8955_1 = {s6040[0]};
    assign in8955_2 = {s6041[0]};
    Full_Adder FA_8955(s8955, c8955, in8955_1, in8955_2, s6039[0]);
    wire[0:0] s8956, in8956_1, in8956_2;
    wire c8956;
    assign in8956_1 = {s6043[0]};
    assign in8956_2 = {s6044[0]};
    Full_Adder FA_8956(s8956, c8956, in8956_1, in8956_2, s6042[0]);
    wire[0:0] s8957, in8957_1, in8957_2;
    wire c8957;
    assign in8957_1 = {s6046[0]};
    assign in8957_2 = {s6047[0]};
    Full_Adder FA_8957(s8957, c8957, in8957_1, in8957_2, s6045[0]);
    wire[0:0] s8958, in8958_1, in8958_2;
    wire c8958;
    assign in8958_1 = {s6049[0]};
    assign in8958_2 = {s6050[0]};
    Full_Adder FA_8958(s8958, c8958, in8958_1, in8958_2, s6048[0]);
    wire[0:0] s8959, in8959_1, in8959_2;
    wire c8959;
    assign in8959_1 = {s6052[0]};
    assign in8959_2 = {s6053[0]};
    Full_Adder FA_8959(s8959, c8959, in8959_1, in8959_2, s6051[0]);
    wire[0:0] s8960, in8960_1, in8960_2;
    wire c8960;
    assign in8960_1 = {c6035};
    assign in8960_2 = {c6036};
    Full_Adder FA_8960(s8960, c8960, in8960_1, in8960_2, s2772[0]);
    wire[0:0] s8961, in8961_1, in8961_2;
    wire c8961;
    assign in8961_1 = {c6038};
    assign in8961_2 = {c6039};
    Full_Adder FA_8961(s8961, c8961, in8961_1, in8961_2, c6037);
    wire[0:0] s8962, in8962_1, in8962_2;
    wire c8962;
    assign in8962_1 = {c6041};
    assign in8962_2 = {c6042};
    Full_Adder FA_8962(s8962, c8962, in8962_1, in8962_2, c6040);
    wire[0:0] s8963, in8963_1, in8963_2;
    wire c8963;
    assign in8963_1 = {c6044};
    assign in8963_2 = {c6045};
    Full_Adder FA_8963(s8963, c8963, in8963_1, in8963_2, c6043);
    wire[0:0] s8964, in8964_1, in8964_2;
    wire c8964;
    assign in8964_1 = {c6047};
    assign in8964_2 = {c6048};
    Full_Adder FA_8964(s8964, c8964, in8964_1, in8964_2, c6046);
    wire[0:0] s8965, in8965_1, in8965_2;
    wire c8965;
    assign in8965_1 = {c6050};
    assign in8965_2 = {c6051};
    Full_Adder FA_8965(s8965, c8965, in8965_1, in8965_2, c6049);
    wire[0:0] s8966, in8966_1, in8966_2;
    wire c8966;
    assign in8966_1 = {c6053};
    assign in8966_2 = {s6054[0]};
    Full_Adder FA_8966(s8966, c8966, in8966_1, in8966_2, c6052);
    wire[0:0] s8967, in8967_1, in8967_2;
    wire c8967;
    assign in8967_1 = {s6056[0]};
    assign in8967_2 = {s6057[0]};
    Full_Adder FA_8967(s8967, c8967, in8967_1, in8967_2, s6055[0]);
    wire[0:0] s8968, in8968_1, in8968_2;
    wire c8968;
    assign in8968_1 = {s6059[0]};
    assign in8968_2 = {s6060[0]};
    Full_Adder FA_8968(s8968, c8968, in8968_1, in8968_2, s6058[0]);
    wire[0:0] s8969, in8969_1, in8969_2;
    wire c8969;
    assign in8969_1 = {s6062[0]};
    assign in8969_2 = {s6063[0]};
    Full_Adder FA_8969(s8969, c8969, in8969_1, in8969_2, s6061[0]);
    wire[0:0] s8970, in8970_1, in8970_2;
    wire c8970;
    assign in8970_1 = {s6065[0]};
    assign in8970_2 = {s6066[0]};
    Full_Adder FA_8970(s8970, c8970, in8970_1, in8970_2, s6064[0]);
    wire[0:0] s8971, in8971_1, in8971_2;
    wire c8971;
    assign in8971_1 = {s6068[0]};
    assign in8971_2 = {s6069[0]};
    Full_Adder FA_8971(s8971, c8971, in8971_1, in8971_2, s6067[0]);
    wire[0:0] s8972, in8972_1, in8972_2;
    wire c8972;
    assign in8972_1 = {s6071[0]};
    assign in8972_2 = {s6072[0]};
    Full_Adder FA_8972(s8972, c8972, in8972_1, in8972_2, s6070[0]);
    wire[0:0] s8973, in8973_1, in8973_2;
    wire c8973;
    assign in8973_1 = {c6054};
    assign in8973_2 = {c6055};
    Full_Adder FA_8973(s8973, c8973, in8973_1, in8973_2, s2800[0]);
    wire[0:0] s8974, in8974_1, in8974_2;
    wire c8974;
    assign in8974_1 = {c6057};
    assign in8974_2 = {c6058};
    Full_Adder FA_8974(s8974, c8974, in8974_1, in8974_2, c6056);
    wire[0:0] s8975, in8975_1, in8975_2;
    wire c8975;
    assign in8975_1 = {c6060};
    assign in8975_2 = {c6061};
    Full_Adder FA_8975(s8975, c8975, in8975_1, in8975_2, c6059);
    wire[0:0] s8976, in8976_1, in8976_2;
    wire c8976;
    assign in8976_1 = {c6063};
    assign in8976_2 = {c6064};
    Full_Adder FA_8976(s8976, c8976, in8976_1, in8976_2, c6062);
    wire[0:0] s8977, in8977_1, in8977_2;
    wire c8977;
    assign in8977_1 = {c6066};
    assign in8977_2 = {c6067};
    Full_Adder FA_8977(s8977, c8977, in8977_1, in8977_2, c6065);
    wire[0:0] s8978, in8978_1, in8978_2;
    wire c8978;
    assign in8978_1 = {c6069};
    assign in8978_2 = {c6070};
    Full_Adder FA_8978(s8978, c8978, in8978_1, in8978_2, c6068);
    wire[0:0] s8979, in8979_1, in8979_2;
    wire c8979;
    assign in8979_1 = {c6072};
    assign in8979_2 = {s6073[0]};
    Full_Adder FA_8979(s8979, c8979, in8979_1, in8979_2, c6071);
    wire[0:0] s8980, in8980_1, in8980_2;
    wire c8980;
    assign in8980_1 = {s6075[0]};
    assign in8980_2 = {s6076[0]};
    Full_Adder FA_8980(s8980, c8980, in8980_1, in8980_2, s6074[0]);
    wire[0:0] s8981, in8981_1, in8981_2;
    wire c8981;
    assign in8981_1 = {s6078[0]};
    assign in8981_2 = {s6079[0]};
    Full_Adder FA_8981(s8981, c8981, in8981_1, in8981_2, s6077[0]);
    wire[0:0] s8982, in8982_1, in8982_2;
    wire c8982;
    assign in8982_1 = {s6081[0]};
    assign in8982_2 = {s6082[0]};
    Full_Adder FA_8982(s8982, c8982, in8982_1, in8982_2, s6080[0]);
    wire[0:0] s8983, in8983_1, in8983_2;
    wire c8983;
    assign in8983_1 = {s6084[0]};
    assign in8983_2 = {s6085[0]};
    Full_Adder FA_8983(s8983, c8983, in8983_1, in8983_2, s6083[0]);
    wire[0:0] s8984, in8984_1, in8984_2;
    wire c8984;
    assign in8984_1 = {s6087[0]};
    assign in8984_2 = {s6088[0]};
    Full_Adder FA_8984(s8984, c8984, in8984_1, in8984_2, s6086[0]);
    wire[0:0] s8985, in8985_1, in8985_2;
    wire c8985;
    assign in8985_1 = {s6090[0]};
    assign in8985_2 = {s6091[0]};
    Full_Adder FA_8985(s8985, c8985, in8985_1, in8985_2, s6089[0]);
    wire[0:0] s8986, in8986_1, in8986_2;
    wire c8986;
    assign in8986_1 = {c6073};
    assign in8986_2 = {c6074};
    Full_Adder FA_8986(s8986, c8986, in8986_1, in8986_2, s2828[0]);
    wire[0:0] s8987, in8987_1, in8987_2;
    wire c8987;
    assign in8987_1 = {c6076};
    assign in8987_2 = {c6077};
    Full_Adder FA_8987(s8987, c8987, in8987_1, in8987_2, c6075);
    wire[0:0] s8988, in8988_1, in8988_2;
    wire c8988;
    assign in8988_1 = {c6079};
    assign in8988_2 = {c6080};
    Full_Adder FA_8988(s8988, c8988, in8988_1, in8988_2, c6078);
    wire[0:0] s8989, in8989_1, in8989_2;
    wire c8989;
    assign in8989_1 = {c6082};
    assign in8989_2 = {c6083};
    Full_Adder FA_8989(s8989, c8989, in8989_1, in8989_2, c6081);
    wire[0:0] s8990, in8990_1, in8990_2;
    wire c8990;
    assign in8990_1 = {c6085};
    assign in8990_2 = {c6086};
    Full_Adder FA_8990(s8990, c8990, in8990_1, in8990_2, c6084);
    wire[0:0] s8991, in8991_1, in8991_2;
    wire c8991;
    assign in8991_1 = {c6088};
    assign in8991_2 = {c6089};
    Full_Adder FA_8991(s8991, c8991, in8991_1, in8991_2, c6087);
    wire[0:0] s8992, in8992_1, in8992_2;
    wire c8992;
    assign in8992_1 = {c6091};
    assign in8992_2 = {s6092[0]};
    Full_Adder FA_8992(s8992, c8992, in8992_1, in8992_2, c6090);
    wire[0:0] s8993, in8993_1, in8993_2;
    wire c8993;
    assign in8993_1 = {s6094[0]};
    assign in8993_2 = {s6095[0]};
    Full_Adder FA_8993(s8993, c8993, in8993_1, in8993_2, s6093[0]);
    wire[0:0] s8994, in8994_1, in8994_2;
    wire c8994;
    assign in8994_1 = {s6097[0]};
    assign in8994_2 = {s6098[0]};
    Full_Adder FA_8994(s8994, c8994, in8994_1, in8994_2, s6096[0]);
    wire[0:0] s8995, in8995_1, in8995_2;
    wire c8995;
    assign in8995_1 = {s6100[0]};
    assign in8995_2 = {s6101[0]};
    Full_Adder FA_8995(s8995, c8995, in8995_1, in8995_2, s6099[0]);
    wire[0:0] s8996, in8996_1, in8996_2;
    wire c8996;
    assign in8996_1 = {s6103[0]};
    assign in8996_2 = {s6104[0]};
    Full_Adder FA_8996(s8996, c8996, in8996_1, in8996_2, s6102[0]);
    wire[0:0] s8997, in8997_1, in8997_2;
    wire c8997;
    assign in8997_1 = {s6106[0]};
    assign in8997_2 = {s6107[0]};
    Full_Adder FA_8997(s8997, c8997, in8997_1, in8997_2, s6105[0]);
    wire[0:0] s8998, in8998_1, in8998_2;
    wire c8998;
    assign in8998_1 = {s6109[0]};
    assign in8998_2 = {s6110[0]};
    Full_Adder FA_8998(s8998, c8998, in8998_1, in8998_2, s6108[0]);
    wire[0:0] s8999, in8999_1, in8999_2;
    wire c8999;
    assign in8999_1 = {c6092};
    assign in8999_2 = {c6093};
    Full_Adder FA_8999(s8999, c8999, in8999_1, in8999_2, s2856[0]);
    wire[0:0] s9000, in9000_1, in9000_2;
    wire c9000;
    assign in9000_1 = {c6095};
    assign in9000_2 = {c6096};
    Full_Adder FA_9000(s9000, c9000, in9000_1, in9000_2, c6094);
    wire[0:0] s9001, in9001_1, in9001_2;
    wire c9001;
    assign in9001_1 = {c6098};
    assign in9001_2 = {c6099};
    Full_Adder FA_9001(s9001, c9001, in9001_1, in9001_2, c6097);
    wire[0:0] s9002, in9002_1, in9002_2;
    wire c9002;
    assign in9002_1 = {c6101};
    assign in9002_2 = {c6102};
    Full_Adder FA_9002(s9002, c9002, in9002_1, in9002_2, c6100);
    wire[0:0] s9003, in9003_1, in9003_2;
    wire c9003;
    assign in9003_1 = {c6104};
    assign in9003_2 = {c6105};
    Full_Adder FA_9003(s9003, c9003, in9003_1, in9003_2, c6103);
    wire[0:0] s9004, in9004_1, in9004_2;
    wire c9004;
    assign in9004_1 = {c6107};
    assign in9004_2 = {c6108};
    Full_Adder FA_9004(s9004, c9004, in9004_1, in9004_2, c6106);
    wire[0:0] s9005, in9005_1, in9005_2;
    wire c9005;
    assign in9005_1 = {c6110};
    assign in9005_2 = {s6111[0]};
    Full_Adder FA_9005(s9005, c9005, in9005_1, in9005_2, c6109);
    wire[0:0] s9006, in9006_1, in9006_2;
    wire c9006;
    assign in9006_1 = {s6113[0]};
    assign in9006_2 = {s6114[0]};
    Full_Adder FA_9006(s9006, c9006, in9006_1, in9006_2, s6112[0]);
    wire[0:0] s9007, in9007_1, in9007_2;
    wire c9007;
    assign in9007_1 = {s6116[0]};
    assign in9007_2 = {s6117[0]};
    Full_Adder FA_9007(s9007, c9007, in9007_1, in9007_2, s6115[0]);
    wire[0:0] s9008, in9008_1, in9008_2;
    wire c9008;
    assign in9008_1 = {s6119[0]};
    assign in9008_2 = {s6120[0]};
    Full_Adder FA_9008(s9008, c9008, in9008_1, in9008_2, s6118[0]);
    wire[0:0] s9009, in9009_1, in9009_2;
    wire c9009;
    assign in9009_1 = {s6122[0]};
    assign in9009_2 = {s6123[0]};
    Full_Adder FA_9009(s9009, c9009, in9009_1, in9009_2, s6121[0]);
    wire[0:0] s9010, in9010_1, in9010_2;
    wire c9010;
    assign in9010_1 = {s6125[0]};
    assign in9010_2 = {s6126[0]};
    Full_Adder FA_9010(s9010, c9010, in9010_1, in9010_2, s6124[0]);
    wire[0:0] s9011, in9011_1, in9011_2;
    wire c9011;
    assign in9011_1 = {s6128[0]};
    assign in9011_2 = {s6129[0]};
    Full_Adder FA_9011(s9011, c9011, in9011_1, in9011_2, s6127[0]);
    wire[0:0] s9012, in9012_1, in9012_2;
    wire c9012;
    assign in9012_1 = {c6111};
    assign in9012_2 = {c6112};
    Full_Adder FA_9012(s9012, c9012, in9012_1, in9012_2, s2884[0]);
    wire[0:0] s9013, in9013_1, in9013_2;
    wire c9013;
    assign in9013_1 = {c6114};
    assign in9013_2 = {c6115};
    Full_Adder FA_9013(s9013, c9013, in9013_1, in9013_2, c6113);
    wire[0:0] s9014, in9014_1, in9014_2;
    wire c9014;
    assign in9014_1 = {c6117};
    assign in9014_2 = {c6118};
    Full_Adder FA_9014(s9014, c9014, in9014_1, in9014_2, c6116);
    wire[0:0] s9015, in9015_1, in9015_2;
    wire c9015;
    assign in9015_1 = {c6120};
    assign in9015_2 = {c6121};
    Full_Adder FA_9015(s9015, c9015, in9015_1, in9015_2, c6119);
    wire[0:0] s9016, in9016_1, in9016_2;
    wire c9016;
    assign in9016_1 = {c6123};
    assign in9016_2 = {c6124};
    Full_Adder FA_9016(s9016, c9016, in9016_1, in9016_2, c6122);
    wire[0:0] s9017, in9017_1, in9017_2;
    wire c9017;
    assign in9017_1 = {c6126};
    assign in9017_2 = {c6127};
    Full_Adder FA_9017(s9017, c9017, in9017_1, in9017_2, c6125);
    wire[0:0] s9018, in9018_1, in9018_2;
    wire c9018;
    assign in9018_1 = {c6129};
    assign in9018_2 = {s6130[0]};
    Full_Adder FA_9018(s9018, c9018, in9018_1, in9018_2, c6128);
    wire[0:0] s9019, in9019_1, in9019_2;
    wire c9019;
    assign in9019_1 = {s6132[0]};
    assign in9019_2 = {s6133[0]};
    Full_Adder FA_9019(s9019, c9019, in9019_1, in9019_2, s6131[0]);
    wire[0:0] s9020, in9020_1, in9020_2;
    wire c9020;
    assign in9020_1 = {s6135[0]};
    assign in9020_2 = {s6136[0]};
    Full_Adder FA_9020(s9020, c9020, in9020_1, in9020_2, s6134[0]);
    wire[0:0] s9021, in9021_1, in9021_2;
    wire c9021;
    assign in9021_1 = {s6138[0]};
    assign in9021_2 = {s6139[0]};
    Full_Adder FA_9021(s9021, c9021, in9021_1, in9021_2, s6137[0]);
    wire[0:0] s9022, in9022_1, in9022_2;
    wire c9022;
    assign in9022_1 = {s6141[0]};
    assign in9022_2 = {s6142[0]};
    Full_Adder FA_9022(s9022, c9022, in9022_1, in9022_2, s6140[0]);
    wire[0:0] s9023, in9023_1, in9023_2;
    wire c9023;
    assign in9023_1 = {s6144[0]};
    assign in9023_2 = {s6145[0]};
    Full_Adder FA_9023(s9023, c9023, in9023_1, in9023_2, s6143[0]);
    wire[0:0] s9024, in9024_1, in9024_2;
    wire c9024;
    assign in9024_1 = {s6147[0]};
    assign in9024_2 = {s6148[0]};
    Full_Adder FA_9024(s9024, c9024, in9024_1, in9024_2, s6146[0]);
    wire[0:0] s9025, in9025_1, in9025_2;
    wire c9025;
    assign in9025_1 = {c6130};
    assign in9025_2 = {c6131};
    Full_Adder FA_9025(s9025, c9025, in9025_1, in9025_2, s2912[0]);
    wire[0:0] s9026, in9026_1, in9026_2;
    wire c9026;
    assign in9026_1 = {c6133};
    assign in9026_2 = {c6134};
    Full_Adder FA_9026(s9026, c9026, in9026_1, in9026_2, c6132);
    wire[0:0] s9027, in9027_1, in9027_2;
    wire c9027;
    assign in9027_1 = {c6136};
    assign in9027_2 = {c6137};
    Full_Adder FA_9027(s9027, c9027, in9027_1, in9027_2, c6135);
    wire[0:0] s9028, in9028_1, in9028_2;
    wire c9028;
    assign in9028_1 = {c6139};
    assign in9028_2 = {c6140};
    Full_Adder FA_9028(s9028, c9028, in9028_1, in9028_2, c6138);
    wire[0:0] s9029, in9029_1, in9029_2;
    wire c9029;
    assign in9029_1 = {c6142};
    assign in9029_2 = {c6143};
    Full_Adder FA_9029(s9029, c9029, in9029_1, in9029_2, c6141);
    wire[0:0] s9030, in9030_1, in9030_2;
    wire c9030;
    assign in9030_1 = {c6145};
    assign in9030_2 = {c6146};
    Full_Adder FA_9030(s9030, c9030, in9030_1, in9030_2, c6144);
    wire[0:0] s9031, in9031_1, in9031_2;
    wire c9031;
    assign in9031_1 = {c6148};
    assign in9031_2 = {s6149[0]};
    Full_Adder FA_9031(s9031, c9031, in9031_1, in9031_2, c6147);
    wire[0:0] s9032, in9032_1, in9032_2;
    wire c9032;
    assign in9032_1 = {s6151[0]};
    assign in9032_2 = {s6152[0]};
    Full_Adder FA_9032(s9032, c9032, in9032_1, in9032_2, s6150[0]);
    wire[0:0] s9033, in9033_1, in9033_2;
    wire c9033;
    assign in9033_1 = {s6154[0]};
    assign in9033_2 = {s6155[0]};
    Full_Adder FA_9033(s9033, c9033, in9033_1, in9033_2, s6153[0]);
    wire[0:0] s9034, in9034_1, in9034_2;
    wire c9034;
    assign in9034_1 = {s6157[0]};
    assign in9034_2 = {s6158[0]};
    Full_Adder FA_9034(s9034, c9034, in9034_1, in9034_2, s6156[0]);
    wire[0:0] s9035, in9035_1, in9035_2;
    wire c9035;
    assign in9035_1 = {s6160[0]};
    assign in9035_2 = {s6161[0]};
    Full_Adder FA_9035(s9035, c9035, in9035_1, in9035_2, s6159[0]);
    wire[0:0] s9036, in9036_1, in9036_2;
    wire c9036;
    assign in9036_1 = {s6163[0]};
    assign in9036_2 = {s6164[0]};
    Full_Adder FA_9036(s9036, c9036, in9036_1, in9036_2, s6162[0]);
    wire[0:0] s9037, in9037_1, in9037_2;
    wire c9037;
    assign in9037_1 = {s6166[0]};
    assign in9037_2 = {s6167[0]};
    Full_Adder FA_9037(s9037, c9037, in9037_1, in9037_2, s6165[0]);
    wire[0:0] s9038, in9038_1, in9038_2;
    wire c9038;
    assign in9038_1 = {c6149};
    assign in9038_2 = {c6150};
    Full_Adder FA_9038(s9038, c9038, in9038_1, in9038_2, s2940[0]);
    wire[0:0] s9039, in9039_1, in9039_2;
    wire c9039;
    assign in9039_1 = {c6152};
    assign in9039_2 = {c6153};
    Full_Adder FA_9039(s9039, c9039, in9039_1, in9039_2, c6151);
    wire[0:0] s9040, in9040_1, in9040_2;
    wire c9040;
    assign in9040_1 = {c6155};
    assign in9040_2 = {c6156};
    Full_Adder FA_9040(s9040, c9040, in9040_1, in9040_2, c6154);
    wire[0:0] s9041, in9041_1, in9041_2;
    wire c9041;
    assign in9041_1 = {c6158};
    assign in9041_2 = {c6159};
    Full_Adder FA_9041(s9041, c9041, in9041_1, in9041_2, c6157);
    wire[0:0] s9042, in9042_1, in9042_2;
    wire c9042;
    assign in9042_1 = {c6161};
    assign in9042_2 = {c6162};
    Full_Adder FA_9042(s9042, c9042, in9042_1, in9042_2, c6160);
    wire[0:0] s9043, in9043_1, in9043_2;
    wire c9043;
    assign in9043_1 = {c6164};
    assign in9043_2 = {c6165};
    Full_Adder FA_9043(s9043, c9043, in9043_1, in9043_2, c6163);
    wire[0:0] s9044, in9044_1, in9044_2;
    wire c9044;
    assign in9044_1 = {c6167};
    assign in9044_2 = {s6168[0]};
    Full_Adder FA_9044(s9044, c9044, in9044_1, in9044_2, c6166);
    wire[0:0] s9045, in9045_1, in9045_2;
    wire c9045;
    assign in9045_1 = {s6170[0]};
    assign in9045_2 = {s6171[0]};
    Full_Adder FA_9045(s9045, c9045, in9045_1, in9045_2, s6169[0]);
    wire[0:0] s9046, in9046_1, in9046_2;
    wire c9046;
    assign in9046_1 = {s6173[0]};
    assign in9046_2 = {s6174[0]};
    Full_Adder FA_9046(s9046, c9046, in9046_1, in9046_2, s6172[0]);
    wire[0:0] s9047, in9047_1, in9047_2;
    wire c9047;
    assign in9047_1 = {s6176[0]};
    assign in9047_2 = {s6177[0]};
    Full_Adder FA_9047(s9047, c9047, in9047_1, in9047_2, s6175[0]);
    wire[0:0] s9048, in9048_1, in9048_2;
    wire c9048;
    assign in9048_1 = {s6179[0]};
    assign in9048_2 = {s6180[0]};
    Full_Adder FA_9048(s9048, c9048, in9048_1, in9048_2, s6178[0]);
    wire[0:0] s9049, in9049_1, in9049_2;
    wire c9049;
    assign in9049_1 = {s6182[0]};
    assign in9049_2 = {s6183[0]};
    Full_Adder FA_9049(s9049, c9049, in9049_1, in9049_2, s6181[0]);
    wire[0:0] s9050, in9050_1, in9050_2;
    wire c9050;
    assign in9050_1 = {s6185[0]};
    assign in9050_2 = {s6186[0]};
    Full_Adder FA_9050(s9050, c9050, in9050_1, in9050_2, s6184[0]);
    wire[0:0] s9051, in9051_1, in9051_2;
    wire c9051;
    assign in9051_1 = {c6168};
    assign in9051_2 = {c6169};
    Full_Adder FA_9051(s9051, c9051, in9051_1, in9051_2, s2968[0]);
    wire[0:0] s9052, in9052_1, in9052_2;
    wire c9052;
    assign in9052_1 = {c6171};
    assign in9052_2 = {c6172};
    Full_Adder FA_9052(s9052, c9052, in9052_1, in9052_2, c6170);
    wire[0:0] s9053, in9053_1, in9053_2;
    wire c9053;
    assign in9053_1 = {c6174};
    assign in9053_2 = {c6175};
    Full_Adder FA_9053(s9053, c9053, in9053_1, in9053_2, c6173);
    wire[0:0] s9054, in9054_1, in9054_2;
    wire c9054;
    assign in9054_1 = {c6177};
    assign in9054_2 = {c6178};
    Full_Adder FA_9054(s9054, c9054, in9054_1, in9054_2, c6176);
    wire[0:0] s9055, in9055_1, in9055_2;
    wire c9055;
    assign in9055_1 = {c6180};
    assign in9055_2 = {c6181};
    Full_Adder FA_9055(s9055, c9055, in9055_1, in9055_2, c6179);
    wire[0:0] s9056, in9056_1, in9056_2;
    wire c9056;
    assign in9056_1 = {c6183};
    assign in9056_2 = {c6184};
    Full_Adder FA_9056(s9056, c9056, in9056_1, in9056_2, c6182);
    wire[0:0] s9057, in9057_1, in9057_2;
    wire c9057;
    assign in9057_1 = {c6186};
    assign in9057_2 = {s6187[0]};
    Full_Adder FA_9057(s9057, c9057, in9057_1, in9057_2, c6185);
    wire[0:0] s9058, in9058_1, in9058_2;
    wire c9058;
    assign in9058_1 = {s6189[0]};
    assign in9058_2 = {s6190[0]};
    Full_Adder FA_9058(s9058, c9058, in9058_1, in9058_2, s6188[0]);
    wire[0:0] s9059, in9059_1, in9059_2;
    wire c9059;
    assign in9059_1 = {s6192[0]};
    assign in9059_2 = {s6193[0]};
    Full_Adder FA_9059(s9059, c9059, in9059_1, in9059_2, s6191[0]);
    wire[0:0] s9060, in9060_1, in9060_2;
    wire c9060;
    assign in9060_1 = {s6195[0]};
    assign in9060_2 = {s6196[0]};
    Full_Adder FA_9060(s9060, c9060, in9060_1, in9060_2, s6194[0]);
    wire[0:0] s9061, in9061_1, in9061_2;
    wire c9061;
    assign in9061_1 = {s6198[0]};
    assign in9061_2 = {s6199[0]};
    Full_Adder FA_9061(s9061, c9061, in9061_1, in9061_2, s6197[0]);
    wire[0:0] s9062, in9062_1, in9062_2;
    wire c9062;
    assign in9062_1 = {s6201[0]};
    assign in9062_2 = {s6202[0]};
    Full_Adder FA_9062(s9062, c9062, in9062_1, in9062_2, s6200[0]);
    wire[0:0] s9063, in9063_1, in9063_2;
    wire c9063;
    assign in9063_1 = {s6204[0]};
    assign in9063_2 = {s6205[0]};
    Full_Adder FA_9063(s9063, c9063, in9063_1, in9063_2, s6203[0]);
    wire[0:0] s9064, in9064_1, in9064_2;
    wire c9064;
    assign in9064_1 = {c6187};
    assign in9064_2 = {c6188};
    Full_Adder FA_9064(s9064, c9064, in9064_1, in9064_2, s2996[0]);
    wire[0:0] s9065, in9065_1, in9065_2;
    wire c9065;
    assign in9065_1 = {c6190};
    assign in9065_2 = {c6191};
    Full_Adder FA_9065(s9065, c9065, in9065_1, in9065_2, c6189);
    wire[0:0] s9066, in9066_1, in9066_2;
    wire c9066;
    assign in9066_1 = {c6193};
    assign in9066_2 = {c6194};
    Full_Adder FA_9066(s9066, c9066, in9066_1, in9066_2, c6192);
    wire[0:0] s9067, in9067_1, in9067_2;
    wire c9067;
    assign in9067_1 = {c6196};
    assign in9067_2 = {c6197};
    Full_Adder FA_9067(s9067, c9067, in9067_1, in9067_2, c6195);
    wire[0:0] s9068, in9068_1, in9068_2;
    wire c9068;
    assign in9068_1 = {c6199};
    assign in9068_2 = {c6200};
    Full_Adder FA_9068(s9068, c9068, in9068_1, in9068_2, c6198);
    wire[0:0] s9069, in9069_1, in9069_2;
    wire c9069;
    assign in9069_1 = {c6202};
    assign in9069_2 = {c6203};
    Full_Adder FA_9069(s9069, c9069, in9069_1, in9069_2, c6201);
    wire[0:0] s9070, in9070_1, in9070_2;
    wire c9070;
    assign in9070_1 = {c6205};
    assign in9070_2 = {s6206[0]};
    Full_Adder FA_9070(s9070, c9070, in9070_1, in9070_2, c6204);
    wire[0:0] s9071, in9071_1, in9071_2;
    wire c9071;
    assign in9071_1 = {s6208[0]};
    assign in9071_2 = {s6209[0]};
    Full_Adder FA_9071(s9071, c9071, in9071_1, in9071_2, s6207[0]);
    wire[0:0] s9072, in9072_1, in9072_2;
    wire c9072;
    assign in9072_1 = {s6211[0]};
    assign in9072_2 = {s6212[0]};
    Full_Adder FA_9072(s9072, c9072, in9072_1, in9072_2, s6210[0]);
    wire[0:0] s9073, in9073_1, in9073_2;
    wire c9073;
    assign in9073_1 = {s6214[0]};
    assign in9073_2 = {s6215[0]};
    Full_Adder FA_9073(s9073, c9073, in9073_1, in9073_2, s6213[0]);
    wire[0:0] s9074, in9074_1, in9074_2;
    wire c9074;
    assign in9074_1 = {s6217[0]};
    assign in9074_2 = {s6218[0]};
    Full_Adder FA_9074(s9074, c9074, in9074_1, in9074_2, s6216[0]);
    wire[0:0] s9075, in9075_1, in9075_2;
    wire c9075;
    assign in9075_1 = {s6220[0]};
    assign in9075_2 = {s6221[0]};
    Full_Adder FA_9075(s9075, c9075, in9075_1, in9075_2, s6219[0]);
    wire[0:0] s9076, in9076_1, in9076_2;
    wire c9076;
    assign in9076_1 = {s6223[0]};
    assign in9076_2 = {s6224[0]};
    Full_Adder FA_9076(s9076, c9076, in9076_1, in9076_2, s6222[0]);
    wire[0:0] s9077, in9077_1, in9077_2;
    wire c9077;
    assign in9077_1 = {c6206};
    assign in9077_2 = {c6207};
    Full_Adder FA_9077(s9077, c9077, in9077_1, in9077_2, s3024[0]);
    wire[0:0] s9078, in9078_1, in9078_2;
    wire c9078;
    assign in9078_1 = {c6209};
    assign in9078_2 = {c6210};
    Full_Adder FA_9078(s9078, c9078, in9078_1, in9078_2, c6208);
    wire[0:0] s9079, in9079_1, in9079_2;
    wire c9079;
    assign in9079_1 = {c6212};
    assign in9079_2 = {c6213};
    Full_Adder FA_9079(s9079, c9079, in9079_1, in9079_2, c6211);
    wire[0:0] s9080, in9080_1, in9080_2;
    wire c9080;
    assign in9080_1 = {c6215};
    assign in9080_2 = {c6216};
    Full_Adder FA_9080(s9080, c9080, in9080_1, in9080_2, c6214);
    wire[0:0] s9081, in9081_1, in9081_2;
    wire c9081;
    assign in9081_1 = {c6218};
    assign in9081_2 = {c6219};
    Full_Adder FA_9081(s9081, c9081, in9081_1, in9081_2, c6217);
    wire[0:0] s9082, in9082_1, in9082_2;
    wire c9082;
    assign in9082_1 = {c6221};
    assign in9082_2 = {c6222};
    Full_Adder FA_9082(s9082, c9082, in9082_1, in9082_2, c6220);
    wire[0:0] s9083, in9083_1, in9083_2;
    wire c9083;
    assign in9083_1 = {c6224};
    assign in9083_2 = {s6225[0]};
    Full_Adder FA_9083(s9083, c9083, in9083_1, in9083_2, c6223);
    wire[0:0] s9084, in9084_1, in9084_2;
    wire c9084;
    assign in9084_1 = {s6227[0]};
    assign in9084_2 = {s6228[0]};
    Full_Adder FA_9084(s9084, c9084, in9084_1, in9084_2, s6226[0]);
    wire[0:0] s9085, in9085_1, in9085_2;
    wire c9085;
    assign in9085_1 = {s6230[0]};
    assign in9085_2 = {s6231[0]};
    Full_Adder FA_9085(s9085, c9085, in9085_1, in9085_2, s6229[0]);
    wire[0:0] s9086, in9086_1, in9086_2;
    wire c9086;
    assign in9086_1 = {s6233[0]};
    assign in9086_2 = {s6234[0]};
    Full_Adder FA_9086(s9086, c9086, in9086_1, in9086_2, s6232[0]);
    wire[0:0] s9087, in9087_1, in9087_2;
    wire c9087;
    assign in9087_1 = {s6236[0]};
    assign in9087_2 = {s6237[0]};
    Full_Adder FA_9087(s9087, c9087, in9087_1, in9087_2, s6235[0]);
    wire[0:0] s9088, in9088_1, in9088_2;
    wire c9088;
    assign in9088_1 = {s6239[0]};
    assign in9088_2 = {s6240[0]};
    Full_Adder FA_9088(s9088, c9088, in9088_1, in9088_2, s6238[0]);
    wire[0:0] s9089, in9089_1, in9089_2;
    wire c9089;
    assign in9089_1 = {s6242[0]};
    assign in9089_2 = {s6243[0]};
    Full_Adder FA_9089(s9089, c9089, in9089_1, in9089_2, s6241[0]);
    wire[0:0] s9090, in9090_1, in9090_2;
    wire c9090;
    assign in9090_1 = {c6225};
    assign in9090_2 = {c6226};
    Full_Adder FA_9090(s9090, c9090, in9090_1, in9090_2, s3052[0]);
    wire[0:0] s9091, in9091_1, in9091_2;
    wire c9091;
    assign in9091_1 = {c6228};
    assign in9091_2 = {c6229};
    Full_Adder FA_9091(s9091, c9091, in9091_1, in9091_2, c6227);
    wire[0:0] s9092, in9092_1, in9092_2;
    wire c9092;
    assign in9092_1 = {c6231};
    assign in9092_2 = {c6232};
    Full_Adder FA_9092(s9092, c9092, in9092_1, in9092_2, c6230);
    wire[0:0] s9093, in9093_1, in9093_2;
    wire c9093;
    assign in9093_1 = {c6234};
    assign in9093_2 = {c6235};
    Full_Adder FA_9093(s9093, c9093, in9093_1, in9093_2, c6233);
    wire[0:0] s9094, in9094_1, in9094_2;
    wire c9094;
    assign in9094_1 = {c6237};
    assign in9094_2 = {c6238};
    Full_Adder FA_9094(s9094, c9094, in9094_1, in9094_2, c6236);
    wire[0:0] s9095, in9095_1, in9095_2;
    wire c9095;
    assign in9095_1 = {c6240};
    assign in9095_2 = {c6241};
    Full_Adder FA_9095(s9095, c9095, in9095_1, in9095_2, c6239);
    wire[0:0] s9096, in9096_1, in9096_2;
    wire c9096;
    assign in9096_1 = {c6243};
    assign in9096_2 = {s6244[0]};
    Full_Adder FA_9096(s9096, c9096, in9096_1, in9096_2, c6242);
    wire[0:0] s9097, in9097_1, in9097_2;
    wire c9097;
    assign in9097_1 = {s6246[0]};
    assign in9097_2 = {s6247[0]};
    Full_Adder FA_9097(s9097, c9097, in9097_1, in9097_2, s6245[0]);
    wire[0:0] s9098, in9098_1, in9098_2;
    wire c9098;
    assign in9098_1 = {s6249[0]};
    assign in9098_2 = {s6250[0]};
    Full_Adder FA_9098(s9098, c9098, in9098_1, in9098_2, s6248[0]);
    wire[0:0] s9099, in9099_1, in9099_2;
    wire c9099;
    assign in9099_1 = {s6252[0]};
    assign in9099_2 = {s6253[0]};
    Full_Adder FA_9099(s9099, c9099, in9099_1, in9099_2, s6251[0]);
    wire[0:0] s9100, in9100_1, in9100_2;
    wire c9100;
    assign in9100_1 = {s6255[0]};
    assign in9100_2 = {s6256[0]};
    Full_Adder FA_9100(s9100, c9100, in9100_1, in9100_2, s6254[0]);
    wire[0:0] s9101, in9101_1, in9101_2;
    wire c9101;
    assign in9101_1 = {s6258[0]};
    assign in9101_2 = {s6259[0]};
    Full_Adder FA_9101(s9101, c9101, in9101_1, in9101_2, s6257[0]);
    wire[0:0] s9102, in9102_1, in9102_2;
    wire c9102;
    assign in9102_1 = {s6261[0]};
    assign in9102_2 = {s6262[0]};
    Full_Adder FA_9102(s9102, c9102, in9102_1, in9102_2, s6260[0]);
    wire[0:0] s9103, in9103_1, in9103_2;
    wire c9103;
    assign in9103_1 = {c6244};
    assign in9103_2 = {c6245};
    Full_Adder FA_9103(s9103, c9103, in9103_1, in9103_2, s3080[0]);
    wire[0:0] s9104, in9104_1, in9104_2;
    wire c9104;
    assign in9104_1 = {c6247};
    assign in9104_2 = {c6248};
    Full_Adder FA_9104(s9104, c9104, in9104_1, in9104_2, c6246);
    wire[0:0] s9105, in9105_1, in9105_2;
    wire c9105;
    assign in9105_1 = {c6250};
    assign in9105_2 = {c6251};
    Full_Adder FA_9105(s9105, c9105, in9105_1, in9105_2, c6249);
    wire[0:0] s9106, in9106_1, in9106_2;
    wire c9106;
    assign in9106_1 = {c6253};
    assign in9106_2 = {c6254};
    Full_Adder FA_9106(s9106, c9106, in9106_1, in9106_2, c6252);
    wire[0:0] s9107, in9107_1, in9107_2;
    wire c9107;
    assign in9107_1 = {c6256};
    assign in9107_2 = {c6257};
    Full_Adder FA_9107(s9107, c9107, in9107_1, in9107_2, c6255);
    wire[0:0] s9108, in9108_1, in9108_2;
    wire c9108;
    assign in9108_1 = {c6259};
    assign in9108_2 = {c6260};
    Full_Adder FA_9108(s9108, c9108, in9108_1, in9108_2, c6258);
    wire[0:0] s9109, in9109_1, in9109_2;
    wire c9109;
    assign in9109_1 = {c6262};
    assign in9109_2 = {s6263[0]};
    Full_Adder FA_9109(s9109, c9109, in9109_1, in9109_2, c6261);
    wire[0:0] s9110, in9110_1, in9110_2;
    wire c9110;
    assign in9110_1 = {s6265[0]};
    assign in9110_2 = {s6266[0]};
    Full_Adder FA_9110(s9110, c9110, in9110_1, in9110_2, s6264[0]);
    wire[0:0] s9111, in9111_1, in9111_2;
    wire c9111;
    assign in9111_1 = {s6268[0]};
    assign in9111_2 = {s6269[0]};
    Full_Adder FA_9111(s9111, c9111, in9111_1, in9111_2, s6267[0]);
    wire[0:0] s9112, in9112_1, in9112_2;
    wire c9112;
    assign in9112_1 = {s6271[0]};
    assign in9112_2 = {s6272[0]};
    Full_Adder FA_9112(s9112, c9112, in9112_1, in9112_2, s6270[0]);
    wire[0:0] s9113, in9113_1, in9113_2;
    wire c9113;
    assign in9113_1 = {s6274[0]};
    assign in9113_2 = {s6275[0]};
    Full_Adder FA_9113(s9113, c9113, in9113_1, in9113_2, s6273[0]);
    wire[0:0] s9114, in9114_1, in9114_2;
    wire c9114;
    assign in9114_1 = {s6277[0]};
    assign in9114_2 = {s6278[0]};
    Full_Adder FA_9114(s9114, c9114, in9114_1, in9114_2, s6276[0]);
    wire[0:0] s9115, in9115_1, in9115_2;
    wire c9115;
    assign in9115_1 = {s6280[0]};
    assign in9115_2 = {s6281[0]};
    Full_Adder FA_9115(s9115, c9115, in9115_1, in9115_2, s6279[0]);
    wire[0:0] s9116, in9116_1, in9116_2;
    wire c9116;
    assign in9116_1 = {c6263};
    assign in9116_2 = {c6264};
    Full_Adder FA_9116(s9116, c9116, in9116_1, in9116_2, s3108[0]);
    wire[0:0] s9117, in9117_1, in9117_2;
    wire c9117;
    assign in9117_1 = {c6266};
    assign in9117_2 = {c6267};
    Full_Adder FA_9117(s9117, c9117, in9117_1, in9117_2, c6265);
    wire[0:0] s9118, in9118_1, in9118_2;
    wire c9118;
    assign in9118_1 = {c6269};
    assign in9118_2 = {c6270};
    Full_Adder FA_9118(s9118, c9118, in9118_1, in9118_2, c6268);
    wire[0:0] s9119, in9119_1, in9119_2;
    wire c9119;
    assign in9119_1 = {c6272};
    assign in9119_2 = {c6273};
    Full_Adder FA_9119(s9119, c9119, in9119_1, in9119_2, c6271);
    wire[0:0] s9120, in9120_1, in9120_2;
    wire c9120;
    assign in9120_1 = {c6275};
    assign in9120_2 = {c6276};
    Full_Adder FA_9120(s9120, c9120, in9120_1, in9120_2, c6274);
    wire[0:0] s9121, in9121_1, in9121_2;
    wire c9121;
    assign in9121_1 = {c6278};
    assign in9121_2 = {c6279};
    Full_Adder FA_9121(s9121, c9121, in9121_1, in9121_2, c6277);
    wire[0:0] s9122, in9122_1, in9122_2;
    wire c9122;
    assign in9122_1 = {c6281};
    assign in9122_2 = {s6282[0]};
    Full_Adder FA_9122(s9122, c9122, in9122_1, in9122_2, c6280);
    wire[0:0] s9123, in9123_1, in9123_2;
    wire c9123;
    assign in9123_1 = {s6284[0]};
    assign in9123_2 = {s6285[0]};
    Full_Adder FA_9123(s9123, c9123, in9123_1, in9123_2, s6283[0]);
    wire[0:0] s9124, in9124_1, in9124_2;
    wire c9124;
    assign in9124_1 = {s6287[0]};
    assign in9124_2 = {s6288[0]};
    Full_Adder FA_9124(s9124, c9124, in9124_1, in9124_2, s6286[0]);
    wire[0:0] s9125, in9125_1, in9125_2;
    wire c9125;
    assign in9125_1 = {s6290[0]};
    assign in9125_2 = {s6291[0]};
    Full_Adder FA_9125(s9125, c9125, in9125_1, in9125_2, s6289[0]);
    wire[0:0] s9126, in9126_1, in9126_2;
    wire c9126;
    assign in9126_1 = {s6293[0]};
    assign in9126_2 = {s6294[0]};
    Full_Adder FA_9126(s9126, c9126, in9126_1, in9126_2, s6292[0]);
    wire[0:0] s9127, in9127_1, in9127_2;
    wire c9127;
    assign in9127_1 = {s6296[0]};
    assign in9127_2 = {s6297[0]};
    Full_Adder FA_9127(s9127, c9127, in9127_1, in9127_2, s6295[0]);
    wire[0:0] s9128, in9128_1, in9128_2;
    wire c9128;
    assign in9128_1 = {s6299[0]};
    assign in9128_2 = {s6300[0]};
    Full_Adder FA_9128(s9128, c9128, in9128_1, in9128_2, s6298[0]);
    wire[0:0] s9129, in9129_1, in9129_2;
    wire c9129;
    assign in9129_1 = {c6282};
    assign in9129_2 = {c6283};
    Full_Adder FA_9129(s9129, c9129, in9129_1, in9129_2, s3136[0]);
    wire[0:0] s9130, in9130_1, in9130_2;
    wire c9130;
    assign in9130_1 = {c6285};
    assign in9130_2 = {c6286};
    Full_Adder FA_9130(s9130, c9130, in9130_1, in9130_2, c6284);
    wire[0:0] s9131, in9131_1, in9131_2;
    wire c9131;
    assign in9131_1 = {c6288};
    assign in9131_2 = {c6289};
    Full_Adder FA_9131(s9131, c9131, in9131_1, in9131_2, c6287);
    wire[0:0] s9132, in9132_1, in9132_2;
    wire c9132;
    assign in9132_1 = {c6291};
    assign in9132_2 = {c6292};
    Full_Adder FA_9132(s9132, c9132, in9132_1, in9132_2, c6290);
    wire[0:0] s9133, in9133_1, in9133_2;
    wire c9133;
    assign in9133_1 = {c6294};
    assign in9133_2 = {c6295};
    Full_Adder FA_9133(s9133, c9133, in9133_1, in9133_2, c6293);
    wire[0:0] s9134, in9134_1, in9134_2;
    wire c9134;
    assign in9134_1 = {c6297};
    assign in9134_2 = {c6298};
    Full_Adder FA_9134(s9134, c9134, in9134_1, in9134_2, c6296);
    wire[0:0] s9135, in9135_1, in9135_2;
    wire c9135;
    assign in9135_1 = {c6300};
    assign in9135_2 = {s6301[0]};
    Full_Adder FA_9135(s9135, c9135, in9135_1, in9135_2, c6299);
    wire[0:0] s9136, in9136_1, in9136_2;
    wire c9136;
    assign in9136_1 = {s6303[0]};
    assign in9136_2 = {s6304[0]};
    Full_Adder FA_9136(s9136, c9136, in9136_1, in9136_2, s6302[0]);
    wire[0:0] s9137, in9137_1, in9137_2;
    wire c9137;
    assign in9137_1 = {s6306[0]};
    assign in9137_2 = {s6307[0]};
    Full_Adder FA_9137(s9137, c9137, in9137_1, in9137_2, s6305[0]);
    wire[0:0] s9138, in9138_1, in9138_2;
    wire c9138;
    assign in9138_1 = {s6309[0]};
    assign in9138_2 = {s6310[0]};
    Full_Adder FA_9138(s9138, c9138, in9138_1, in9138_2, s6308[0]);
    wire[0:0] s9139, in9139_1, in9139_2;
    wire c9139;
    assign in9139_1 = {s6312[0]};
    assign in9139_2 = {s6313[0]};
    Full_Adder FA_9139(s9139, c9139, in9139_1, in9139_2, s6311[0]);
    wire[0:0] s9140, in9140_1, in9140_2;
    wire c9140;
    assign in9140_1 = {s6315[0]};
    assign in9140_2 = {s6316[0]};
    Full_Adder FA_9140(s9140, c9140, in9140_1, in9140_2, s6314[0]);
    wire[0:0] s9141, in9141_1, in9141_2;
    wire c9141;
    assign in9141_1 = {s6318[0]};
    assign in9141_2 = {s6319[0]};
    Full_Adder FA_9141(s9141, c9141, in9141_1, in9141_2, s6317[0]);
    wire[0:0] s9142, in9142_1, in9142_2;
    wire c9142;
    assign in9142_1 = {c6301};
    assign in9142_2 = {c6302};
    Full_Adder FA_9142(s9142, c9142, in9142_1, in9142_2, s3164[0]);
    wire[0:0] s9143, in9143_1, in9143_2;
    wire c9143;
    assign in9143_1 = {c6304};
    assign in9143_2 = {c6305};
    Full_Adder FA_9143(s9143, c9143, in9143_1, in9143_2, c6303);
    wire[0:0] s9144, in9144_1, in9144_2;
    wire c9144;
    assign in9144_1 = {c6307};
    assign in9144_2 = {c6308};
    Full_Adder FA_9144(s9144, c9144, in9144_1, in9144_2, c6306);
    wire[0:0] s9145, in9145_1, in9145_2;
    wire c9145;
    assign in9145_1 = {c6310};
    assign in9145_2 = {c6311};
    Full_Adder FA_9145(s9145, c9145, in9145_1, in9145_2, c6309);
    wire[0:0] s9146, in9146_1, in9146_2;
    wire c9146;
    assign in9146_1 = {c6313};
    assign in9146_2 = {c6314};
    Full_Adder FA_9146(s9146, c9146, in9146_1, in9146_2, c6312);
    wire[0:0] s9147, in9147_1, in9147_2;
    wire c9147;
    assign in9147_1 = {c6316};
    assign in9147_2 = {c6317};
    Full_Adder FA_9147(s9147, c9147, in9147_1, in9147_2, c6315);
    wire[0:0] s9148, in9148_1, in9148_2;
    wire c9148;
    assign in9148_1 = {c6319};
    assign in9148_2 = {s6320[0]};
    Full_Adder FA_9148(s9148, c9148, in9148_1, in9148_2, c6318);
    wire[0:0] s9149, in9149_1, in9149_2;
    wire c9149;
    assign in9149_1 = {s6322[0]};
    assign in9149_2 = {s6323[0]};
    Full_Adder FA_9149(s9149, c9149, in9149_1, in9149_2, s6321[0]);
    wire[0:0] s9150, in9150_1, in9150_2;
    wire c9150;
    assign in9150_1 = {s6325[0]};
    assign in9150_2 = {s6326[0]};
    Full_Adder FA_9150(s9150, c9150, in9150_1, in9150_2, s6324[0]);
    wire[0:0] s9151, in9151_1, in9151_2;
    wire c9151;
    assign in9151_1 = {s6328[0]};
    assign in9151_2 = {s6329[0]};
    Full_Adder FA_9151(s9151, c9151, in9151_1, in9151_2, s6327[0]);
    wire[0:0] s9152, in9152_1, in9152_2;
    wire c9152;
    assign in9152_1 = {s6331[0]};
    assign in9152_2 = {s6332[0]};
    Full_Adder FA_9152(s9152, c9152, in9152_1, in9152_2, s6330[0]);
    wire[0:0] s9153, in9153_1, in9153_2;
    wire c9153;
    assign in9153_1 = {s6334[0]};
    assign in9153_2 = {s6335[0]};
    Full_Adder FA_9153(s9153, c9153, in9153_1, in9153_2, s6333[0]);
    wire[0:0] s9154, in9154_1, in9154_2;
    wire c9154;
    assign in9154_1 = {s6337[0]};
    assign in9154_2 = {s6338[0]};
    Full_Adder FA_9154(s9154, c9154, in9154_1, in9154_2, s6336[0]);
    wire[0:0] s9155, in9155_1, in9155_2;
    wire c9155;
    assign in9155_1 = {c6320};
    assign in9155_2 = {c6321};
    Full_Adder FA_9155(s9155, c9155, in9155_1, in9155_2, s3192[0]);
    wire[0:0] s9156, in9156_1, in9156_2;
    wire c9156;
    assign in9156_1 = {c6323};
    assign in9156_2 = {c6324};
    Full_Adder FA_9156(s9156, c9156, in9156_1, in9156_2, c6322);
    wire[0:0] s9157, in9157_1, in9157_2;
    wire c9157;
    assign in9157_1 = {c6326};
    assign in9157_2 = {c6327};
    Full_Adder FA_9157(s9157, c9157, in9157_1, in9157_2, c6325);
    wire[0:0] s9158, in9158_1, in9158_2;
    wire c9158;
    assign in9158_1 = {c6329};
    assign in9158_2 = {c6330};
    Full_Adder FA_9158(s9158, c9158, in9158_1, in9158_2, c6328);
    wire[0:0] s9159, in9159_1, in9159_2;
    wire c9159;
    assign in9159_1 = {c6332};
    assign in9159_2 = {c6333};
    Full_Adder FA_9159(s9159, c9159, in9159_1, in9159_2, c6331);
    wire[0:0] s9160, in9160_1, in9160_2;
    wire c9160;
    assign in9160_1 = {c6335};
    assign in9160_2 = {c6336};
    Full_Adder FA_9160(s9160, c9160, in9160_1, in9160_2, c6334);
    wire[0:0] s9161, in9161_1, in9161_2;
    wire c9161;
    assign in9161_1 = {c6338};
    assign in9161_2 = {s6339[0]};
    Full_Adder FA_9161(s9161, c9161, in9161_1, in9161_2, c6337);
    wire[0:0] s9162, in9162_1, in9162_2;
    wire c9162;
    assign in9162_1 = {s6341[0]};
    assign in9162_2 = {s6342[0]};
    Full_Adder FA_9162(s9162, c9162, in9162_1, in9162_2, s6340[0]);
    wire[0:0] s9163, in9163_1, in9163_2;
    wire c9163;
    assign in9163_1 = {s6344[0]};
    assign in9163_2 = {s6345[0]};
    Full_Adder FA_9163(s9163, c9163, in9163_1, in9163_2, s6343[0]);
    wire[0:0] s9164, in9164_1, in9164_2;
    wire c9164;
    assign in9164_1 = {s6347[0]};
    assign in9164_2 = {s6348[0]};
    Full_Adder FA_9164(s9164, c9164, in9164_1, in9164_2, s6346[0]);
    wire[0:0] s9165, in9165_1, in9165_2;
    wire c9165;
    assign in9165_1 = {s6350[0]};
    assign in9165_2 = {s6351[0]};
    Full_Adder FA_9165(s9165, c9165, in9165_1, in9165_2, s6349[0]);
    wire[0:0] s9166, in9166_1, in9166_2;
    wire c9166;
    assign in9166_1 = {s6353[0]};
    assign in9166_2 = {s6354[0]};
    Full_Adder FA_9166(s9166, c9166, in9166_1, in9166_2, s6352[0]);
    wire[0:0] s9167, in9167_1, in9167_2;
    wire c9167;
    assign in9167_1 = {s6356[0]};
    assign in9167_2 = {s6357[0]};
    Full_Adder FA_9167(s9167, c9167, in9167_1, in9167_2, s6355[0]);
    wire[0:0] s9168, in9168_1, in9168_2;
    wire c9168;
    assign in9168_1 = {c6339};
    assign in9168_2 = {c6340};
    Full_Adder FA_9168(s9168, c9168, in9168_1, in9168_2, s3220[0]);
    wire[0:0] s9169, in9169_1, in9169_2;
    wire c9169;
    assign in9169_1 = {c6342};
    assign in9169_2 = {c6343};
    Full_Adder FA_9169(s9169, c9169, in9169_1, in9169_2, c6341);
    wire[0:0] s9170, in9170_1, in9170_2;
    wire c9170;
    assign in9170_1 = {c6345};
    assign in9170_2 = {c6346};
    Full_Adder FA_9170(s9170, c9170, in9170_1, in9170_2, c6344);
    wire[0:0] s9171, in9171_1, in9171_2;
    wire c9171;
    assign in9171_1 = {c6348};
    assign in9171_2 = {c6349};
    Full_Adder FA_9171(s9171, c9171, in9171_1, in9171_2, c6347);
    wire[0:0] s9172, in9172_1, in9172_2;
    wire c9172;
    assign in9172_1 = {c6351};
    assign in9172_2 = {c6352};
    Full_Adder FA_9172(s9172, c9172, in9172_1, in9172_2, c6350);
    wire[0:0] s9173, in9173_1, in9173_2;
    wire c9173;
    assign in9173_1 = {c6354};
    assign in9173_2 = {c6355};
    Full_Adder FA_9173(s9173, c9173, in9173_1, in9173_2, c6353);
    wire[0:0] s9174, in9174_1, in9174_2;
    wire c9174;
    assign in9174_1 = {c6357};
    assign in9174_2 = {s6358[0]};
    Full_Adder FA_9174(s9174, c9174, in9174_1, in9174_2, c6356);
    wire[0:0] s9175, in9175_1, in9175_2;
    wire c9175;
    assign in9175_1 = {s6360[0]};
    assign in9175_2 = {s6361[0]};
    Full_Adder FA_9175(s9175, c9175, in9175_1, in9175_2, s6359[0]);
    wire[0:0] s9176, in9176_1, in9176_2;
    wire c9176;
    assign in9176_1 = {s6363[0]};
    assign in9176_2 = {s6364[0]};
    Full_Adder FA_9176(s9176, c9176, in9176_1, in9176_2, s6362[0]);
    wire[0:0] s9177, in9177_1, in9177_2;
    wire c9177;
    assign in9177_1 = {s6366[0]};
    assign in9177_2 = {s6367[0]};
    Full_Adder FA_9177(s9177, c9177, in9177_1, in9177_2, s6365[0]);
    wire[0:0] s9178, in9178_1, in9178_2;
    wire c9178;
    assign in9178_1 = {s6369[0]};
    assign in9178_2 = {s6370[0]};
    Full_Adder FA_9178(s9178, c9178, in9178_1, in9178_2, s6368[0]);
    wire[0:0] s9179, in9179_1, in9179_2;
    wire c9179;
    assign in9179_1 = {s6372[0]};
    assign in9179_2 = {s6373[0]};
    Full_Adder FA_9179(s9179, c9179, in9179_1, in9179_2, s6371[0]);
    wire[0:0] s9180, in9180_1, in9180_2;
    wire c9180;
    assign in9180_1 = {s6375[0]};
    assign in9180_2 = {s6376[0]};
    Full_Adder FA_9180(s9180, c9180, in9180_1, in9180_2, s6374[0]);
    wire[0:0] s9181, in9181_1, in9181_2;
    wire c9181;
    assign in9181_1 = {c6358};
    assign in9181_2 = {c6359};
    Full_Adder FA_9181(s9181, c9181, in9181_1, in9181_2, s3248[0]);
    wire[0:0] s9182, in9182_1, in9182_2;
    wire c9182;
    assign in9182_1 = {c6361};
    assign in9182_2 = {c6362};
    Full_Adder FA_9182(s9182, c9182, in9182_1, in9182_2, c6360);
    wire[0:0] s9183, in9183_1, in9183_2;
    wire c9183;
    assign in9183_1 = {c6364};
    assign in9183_2 = {c6365};
    Full_Adder FA_9183(s9183, c9183, in9183_1, in9183_2, c6363);
    wire[0:0] s9184, in9184_1, in9184_2;
    wire c9184;
    assign in9184_1 = {c6367};
    assign in9184_2 = {c6368};
    Full_Adder FA_9184(s9184, c9184, in9184_1, in9184_2, c6366);
    wire[0:0] s9185, in9185_1, in9185_2;
    wire c9185;
    assign in9185_1 = {c6370};
    assign in9185_2 = {c6371};
    Full_Adder FA_9185(s9185, c9185, in9185_1, in9185_2, c6369);
    wire[0:0] s9186, in9186_1, in9186_2;
    wire c9186;
    assign in9186_1 = {c6373};
    assign in9186_2 = {c6374};
    Full_Adder FA_9186(s9186, c9186, in9186_1, in9186_2, c6372);
    wire[0:0] s9187, in9187_1, in9187_2;
    wire c9187;
    assign in9187_1 = {c6376};
    assign in9187_2 = {s6377[0]};
    Full_Adder FA_9187(s9187, c9187, in9187_1, in9187_2, c6375);
    wire[0:0] s9188, in9188_1, in9188_2;
    wire c9188;
    assign in9188_1 = {s6379[0]};
    assign in9188_2 = {s6380[0]};
    Full_Adder FA_9188(s9188, c9188, in9188_1, in9188_2, s6378[0]);
    wire[0:0] s9189, in9189_1, in9189_2;
    wire c9189;
    assign in9189_1 = {s6382[0]};
    assign in9189_2 = {s6383[0]};
    Full_Adder FA_9189(s9189, c9189, in9189_1, in9189_2, s6381[0]);
    wire[0:0] s9190, in9190_1, in9190_2;
    wire c9190;
    assign in9190_1 = {s6385[0]};
    assign in9190_2 = {s6386[0]};
    Full_Adder FA_9190(s9190, c9190, in9190_1, in9190_2, s6384[0]);
    wire[0:0] s9191, in9191_1, in9191_2;
    wire c9191;
    assign in9191_1 = {s6388[0]};
    assign in9191_2 = {s6389[0]};
    Full_Adder FA_9191(s9191, c9191, in9191_1, in9191_2, s6387[0]);
    wire[0:0] s9192, in9192_1, in9192_2;
    wire c9192;
    assign in9192_1 = {s6391[0]};
    assign in9192_2 = {s6392[0]};
    Full_Adder FA_9192(s9192, c9192, in9192_1, in9192_2, s6390[0]);
    wire[0:0] s9193, in9193_1, in9193_2;
    wire c9193;
    assign in9193_1 = {s6394[0]};
    assign in9193_2 = {s6395[0]};
    Full_Adder FA_9193(s9193, c9193, in9193_1, in9193_2, s6393[0]);
    wire[0:0] s9194, in9194_1, in9194_2;
    wire c9194;
    assign in9194_1 = {c6377};
    assign in9194_2 = {c6378};
    Full_Adder FA_9194(s9194, c9194, in9194_1, in9194_2, s3276[0]);
    wire[0:0] s9195, in9195_1, in9195_2;
    wire c9195;
    assign in9195_1 = {c6380};
    assign in9195_2 = {c6381};
    Full_Adder FA_9195(s9195, c9195, in9195_1, in9195_2, c6379);
    wire[0:0] s9196, in9196_1, in9196_2;
    wire c9196;
    assign in9196_1 = {c6383};
    assign in9196_2 = {c6384};
    Full_Adder FA_9196(s9196, c9196, in9196_1, in9196_2, c6382);
    wire[0:0] s9197, in9197_1, in9197_2;
    wire c9197;
    assign in9197_1 = {c6386};
    assign in9197_2 = {c6387};
    Full_Adder FA_9197(s9197, c9197, in9197_1, in9197_2, c6385);
    wire[0:0] s9198, in9198_1, in9198_2;
    wire c9198;
    assign in9198_1 = {c6389};
    assign in9198_2 = {c6390};
    Full_Adder FA_9198(s9198, c9198, in9198_1, in9198_2, c6388);
    wire[0:0] s9199, in9199_1, in9199_2;
    wire c9199;
    assign in9199_1 = {c6392};
    assign in9199_2 = {c6393};
    Full_Adder FA_9199(s9199, c9199, in9199_1, in9199_2, c6391);
    wire[0:0] s9200, in9200_1, in9200_2;
    wire c9200;
    assign in9200_1 = {c6395};
    assign in9200_2 = {s6396[0]};
    Full_Adder FA_9200(s9200, c9200, in9200_1, in9200_2, c6394);
    wire[0:0] s9201, in9201_1, in9201_2;
    wire c9201;
    assign in9201_1 = {s6398[0]};
    assign in9201_2 = {s6399[0]};
    Full_Adder FA_9201(s9201, c9201, in9201_1, in9201_2, s6397[0]);
    wire[0:0] s9202, in9202_1, in9202_2;
    wire c9202;
    assign in9202_1 = {s6401[0]};
    assign in9202_2 = {s6402[0]};
    Full_Adder FA_9202(s9202, c9202, in9202_1, in9202_2, s6400[0]);
    wire[0:0] s9203, in9203_1, in9203_2;
    wire c9203;
    assign in9203_1 = {s6404[0]};
    assign in9203_2 = {s6405[0]};
    Full_Adder FA_9203(s9203, c9203, in9203_1, in9203_2, s6403[0]);
    wire[0:0] s9204, in9204_1, in9204_2;
    wire c9204;
    assign in9204_1 = {s6407[0]};
    assign in9204_2 = {s6408[0]};
    Full_Adder FA_9204(s9204, c9204, in9204_1, in9204_2, s6406[0]);
    wire[0:0] s9205, in9205_1, in9205_2;
    wire c9205;
    assign in9205_1 = {s6410[0]};
    assign in9205_2 = {s6411[0]};
    Full_Adder FA_9205(s9205, c9205, in9205_1, in9205_2, s6409[0]);
    wire[0:0] s9206, in9206_1, in9206_2;
    wire c9206;
    assign in9206_1 = {s6413[0]};
    assign in9206_2 = {s6414[0]};
    Full_Adder FA_9206(s9206, c9206, in9206_1, in9206_2, s6412[0]);
    wire[0:0] s9207, in9207_1, in9207_2;
    wire c9207;
    assign in9207_1 = {c6396};
    assign in9207_2 = {c6397};
    Full_Adder FA_9207(s9207, c9207, in9207_1, in9207_2, s3304[0]);
    wire[0:0] s9208, in9208_1, in9208_2;
    wire c9208;
    assign in9208_1 = {c6399};
    assign in9208_2 = {c6400};
    Full_Adder FA_9208(s9208, c9208, in9208_1, in9208_2, c6398);
    wire[0:0] s9209, in9209_1, in9209_2;
    wire c9209;
    assign in9209_1 = {c6402};
    assign in9209_2 = {c6403};
    Full_Adder FA_9209(s9209, c9209, in9209_1, in9209_2, c6401);
    wire[0:0] s9210, in9210_1, in9210_2;
    wire c9210;
    assign in9210_1 = {c6405};
    assign in9210_2 = {c6406};
    Full_Adder FA_9210(s9210, c9210, in9210_1, in9210_2, c6404);
    wire[0:0] s9211, in9211_1, in9211_2;
    wire c9211;
    assign in9211_1 = {c6408};
    assign in9211_2 = {c6409};
    Full_Adder FA_9211(s9211, c9211, in9211_1, in9211_2, c6407);
    wire[0:0] s9212, in9212_1, in9212_2;
    wire c9212;
    assign in9212_1 = {c6411};
    assign in9212_2 = {c6412};
    Full_Adder FA_9212(s9212, c9212, in9212_1, in9212_2, c6410);
    wire[0:0] s9213, in9213_1, in9213_2;
    wire c9213;
    assign in9213_1 = {c6414};
    assign in9213_2 = {s6415[0]};
    Full_Adder FA_9213(s9213, c9213, in9213_1, in9213_2, c6413);
    wire[0:0] s9214, in9214_1, in9214_2;
    wire c9214;
    assign in9214_1 = {s6417[0]};
    assign in9214_2 = {s6418[0]};
    Full_Adder FA_9214(s9214, c9214, in9214_1, in9214_2, s6416[0]);
    wire[0:0] s9215, in9215_1, in9215_2;
    wire c9215;
    assign in9215_1 = {s6420[0]};
    assign in9215_2 = {s6421[0]};
    Full_Adder FA_9215(s9215, c9215, in9215_1, in9215_2, s6419[0]);
    wire[0:0] s9216, in9216_1, in9216_2;
    wire c9216;
    assign in9216_1 = {s6423[0]};
    assign in9216_2 = {s6424[0]};
    Full_Adder FA_9216(s9216, c9216, in9216_1, in9216_2, s6422[0]);
    wire[0:0] s9217, in9217_1, in9217_2;
    wire c9217;
    assign in9217_1 = {s6426[0]};
    assign in9217_2 = {s6427[0]};
    Full_Adder FA_9217(s9217, c9217, in9217_1, in9217_2, s6425[0]);
    wire[0:0] s9218, in9218_1, in9218_2;
    wire c9218;
    assign in9218_1 = {s6429[0]};
    assign in9218_2 = {s6430[0]};
    Full_Adder FA_9218(s9218, c9218, in9218_1, in9218_2, s6428[0]);
    wire[0:0] s9219, in9219_1, in9219_2;
    wire c9219;
    assign in9219_1 = {s6432[0]};
    assign in9219_2 = {s6433[0]};
    Full_Adder FA_9219(s9219, c9219, in9219_1, in9219_2, s6431[0]);
    wire[0:0] s9220, in9220_1, in9220_2;
    wire c9220;
    assign in9220_1 = {c6415};
    assign in9220_2 = {c6416};
    Full_Adder FA_9220(s9220, c9220, in9220_1, in9220_2, s3332[0]);
    wire[0:0] s9221, in9221_1, in9221_2;
    wire c9221;
    assign in9221_1 = {c6418};
    assign in9221_2 = {c6419};
    Full_Adder FA_9221(s9221, c9221, in9221_1, in9221_2, c6417);
    wire[0:0] s9222, in9222_1, in9222_2;
    wire c9222;
    assign in9222_1 = {c6421};
    assign in9222_2 = {c6422};
    Full_Adder FA_9222(s9222, c9222, in9222_1, in9222_2, c6420);
    wire[0:0] s9223, in9223_1, in9223_2;
    wire c9223;
    assign in9223_1 = {c6424};
    assign in9223_2 = {c6425};
    Full_Adder FA_9223(s9223, c9223, in9223_1, in9223_2, c6423);
    wire[0:0] s9224, in9224_1, in9224_2;
    wire c9224;
    assign in9224_1 = {c6427};
    assign in9224_2 = {c6428};
    Full_Adder FA_9224(s9224, c9224, in9224_1, in9224_2, c6426);
    wire[0:0] s9225, in9225_1, in9225_2;
    wire c9225;
    assign in9225_1 = {c6430};
    assign in9225_2 = {c6431};
    Full_Adder FA_9225(s9225, c9225, in9225_1, in9225_2, c6429);
    wire[0:0] s9226, in9226_1, in9226_2;
    wire c9226;
    assign in9226_1 = {c6433};
    assign in9226_2 = {s6434[0]};
    Full_Adder FA_9226(s9226, c9226, in9226_1, in9226_2, c6432);
    wire[0:0] s9227, in9227_1, in9227_2;
    wire c9227;
    assign in9227_1 = {s6436[0]};
    assign in9227_2 = {s6437[0]};
    Full_Adder FA_9227(s9227, c9227, in9227_1, in9227_2, s6435[0]);
    wire[0:0] s9228, in9228_1, in9228_2;
    wire c9228;
    assign in9228_1 = {s6439[0]};
    assign in9228_2 = {s6440[0]};
    Full_Adder FA_9228(s9228, c9228, in9228_1, in9228_2, s6438[0]);
    wire[0:0] s9229, in9229_1, in9229_2;
    wire c9229;
    assign in9229_1 = {s6442[0]};
    assign in9229_2 = {s6443[0]};
    Full_Adder FA_9229(s9229, c9229, in9229_1, in9229_2, s6441[0]);
    wire[0:0] s9230, in9230_1, in9230_2;
    wire c9230;
    assign in9230_1 = {s6445[0]};
    assign in9230_2 = {s6446[0]};
    Full_Adder FA_9230(s9230, c9230, in9230_1, in9230_2, s6444[0]);
    wire[0:0] s9231, in9231_1, in9231_2;
    wire c9231;
    assign in9231_1 = {s6448[0]};
    assign in9231_2 = {s6449[0]};
    Full_Adder FA_9231(s9231, c9231, in9231_1, in9231_2, s6447[0]);
    wire[0:0] s9232, in9232_1, in9232_2;
    wire c9232;
    assign in9232_1 = {s6451[0]};
    assign in9232_2 = {s6452[0]};
    Full_Adder FA_9232(s9232, c9232, in9232_1, in9232_2, s6450[0]);
    wire[0:0] s9233, in9233_1, in9233_2;
    wire c9233;
    assign in9233_1 = {c6434};
    assign in9233_2 = {c6435};
    Full_Adder FA_9233(s9233, c9233, in9233_1, in9233_2, s3360[0]);
    wire[0:0] s9234, in9234_1, in9234_2;
    wire c9234;
    assign in9234_1 = {c6437};
    assign in9234_2 = {c6438};
    Full_Adder FA_9234(s9234, c9234, in9234_1, in9234_2, c6436);
    wire[0:0] s9235, in9235_1, in9235_2;
    wire c9235;
    assign in9235_1 = {c6440};
    assign in9235_2 = {c6441};
    Full_Adder FA_9235(s9235, c9235, in9235_1, in9235_2, c6439);
    wire[0:0] s9236, in9236_1, in9236_2;
    wire c9236;
    assign in9236_1 = {c6443};
    assign in9236_2 = {c6444};
    Full_Adder FA_9236(s9236, c9236, in9236_1, in9236_2, c6442);
    wire[0:0] s9237, in9237_1, in9237_2;
    wire c9237;
    assign in9237_1 = {c6446};
    assign in9237_2 = {c6447};
    Full_Adder FA_9237(s9237, c9237, in9237_1, in9237_2, c6445);
    wire[0:0] s9238, in9238_1, in9238_2;
    wire c9238;
    assign in9238_1 = {c6449};
    assign in9238_2 = {c6450};
    Full_Adder FA_9238(s9238, c9238, in9238_1, in9238_2, c6448);
    wire[0:0] s9239, in9239_1, in9239_2;
    wire c9239;
    assign in9239_1 = {c6452};
    assign in9239_2 = {s6453[0]};
    Full_Adder FA_9239(s9239, c9239, in9239_1, in9239_2, c6451);
    wire[0:0] s9240, in9240_1, in9240_2;
    wire c9240;
    assign in9240_1 = {s6455[0]};
    assign in9240_2 = {s6456[0]};
    Full_Adder FA_9240(s9240, c9240, in9240_1, in9240_2, s6454[0]);
    wire[0:0] s9241, in9241_1, in9241_2;
    wire c9241;
    assign in9241_1 = {s6458[0]};
    assign in9241_2 = {s6459[0]};
    Full_Adder FA_9241(s9241, c9241, in9241_1, in9241_2, s6457[0]);
    wire[0:0] s9242, in9242_1, in9242_2;
    wire c9242;
    assign in9242_1 = {s6461[0]};
    assign in9242_2 = {s6462[0]};
    Full_Adder FA_9242(s9242, c9242, in9242_1, in9242_2, s6460[0]);
    wire[0:0] s9243, in9243_1, in9243_2;
    wire c9243;
    assign in9243_1 = {s6464[0]};
    assign in9243_2 = {s6465[0]};
    Full_Adder FA_9243(s9243, c9243, in9243_1, in9243_2, s6463[0]);
    wire[0:0] s9244, in9244_1, in9244_2;
    wire c9244;
    assign in9244_1 = {s6467[0]};
    assign in9244_2 = {s6468[0]};
    Full_Adder FA_9244(s9244, c9244, in9244_1, in9244_2, s6466[0]);
    wire[0:0] s9245, in9245_1, in9245_2;
    wire c9245;
    assign in9245_1 = {s6470[0]};
    assign in9245_2 = {s6471[0]};
    Full_Adder FA_9245(s9245, c9245, in9245_1, in9245_2, s6469[0]);
    wire[0:0] s9246, in9246_1, in9246_2;
    wire c9246;
    assign in9246_1 = {c6453};
    assign in9246_2 = {c6454};
    Full_Adder FA_9246(s9246, c9246, in9246_1, in9246_2, s3388[0]);
    wire[0:0] s9247, in9247_1, in9247_2;
    wire c9247;
    assign in9247_1 = {c6456};
    assign in9247_2 = {c6457};
    Full_Adder FA_9247(s9247, c9247, in9247_1, in9247_2, c6455);
    wire[0:0] s9248, in9248_1, in9248_2;
    wire c9248;
    assign in9248_1 = {c6459};
    assign in9248_2 = {c6460};
    Full_Adder FA_9248(s9248, c9248, in9248_1, in9248_2, c6458);
    wire[0:0] s9249, in9249_1, in9249_2;
    wire c9249;
    assign in9249_1 = {c6462};
    assign in9249_2 = {c6463};
    Full_Adder FA_9249(s9249, c9249, in9249_1, in9249_2, c6461);
    wire[0:0] s9250, in9250_1, in9250_2;
    wire c9250;
    assign in9250_1 = {c6465};
    assign in9250_2 = {c6466};
    Full_Adder FA_9250(s9250, c9250, in9250_1, in9250_2, c6464);
    wire[0:0] s9251, in9251_1, in9251_2;
    wire c9251;
    assign in9251_1 = {c6468};
    assign in9251_2 = {c6469};
    Full_Adder FA_9251(s9251, c9251, in9251_1, in9251_2, c6467);
    wire[0:0] s9252, in9252_1, in9252_2;
    wire c9252;
    assign in9252_1 = {c6471};
    assign in9252_2 = {s6472[0]};
    Full_Adder FA_9252(s9252, c9252, in9252_1, in9252_2, c6470);
    wire[0:0] s9253, in9253_1, in9253_2;
    wire c9253;
    assign in9253_1 = {s6474[0]};
    assign in9253_2 = {s6475[0]};
    Full_Adder FA_9253(s9253, c9253, in9253_1, in9253_2, s6473[0]);
    wire[0:0] s9254, in9254_1, in9254_2;
    wire c9254;
    assign in9254_1 = {s6477[0]};
    assign in9254_2 = {s6478[0]};
    Full_Adder FA_9254(s9254, c9254, in9254_1, in9254_2, s6476[0]);
    wire[0:0] s9255, in9255_1, in9255_2;
    wire c9255;
    assign in9255_1 = {s6480[0]};
    assign in9255_2 = {s6481[0]};
    Full_Adder FA_9255(s9255, c9255, in9255_1, in9255_2, s6479[0]);
    wire[0:0] s9256, in9256_1, in9256_2;
    wire c9256;
    assign in9256_1 = {s6483[0]};
    assign in9256_2 = {s6484[0]};
    Full_Adder FA_9256(s9256, c9256, in9256_1, in9256_2, s6482[0]);
    wire[0:0] s9257, in9257_1, in9257_2;
    wire c9257;
    assign in9257_1 = {s6486[0]};
    assign in9257_2 = {s6487[0]};
    Full_Adder FA_9257(s9257, c9257, in9257_1, in9257_2, s6485[0]);
    wire[0:0] s9258, in9258_1, in9258_2;
    wire c9258;
    assign in9258_1 = {s6489[0]};
    assign in9258_2 = {s6490[0]};
    Full_Adder FA_9258(s9258, c9258, in9258_1, in9258_2, s6488[0]);
    wire[0:0] s9259, in9259_1, in9259_2;
    wire c9259;
    assign in9259_1 = {c6472};
    assign in9259_2 = {c6473};
    Full_Adder FA_9259(s9259, c9259, in9259_1, in9259_2, s3416[0]);
    wire[0:0] s9260, in9260_1, in9260_2;
    wire c9260;
    assign in9260_1 = {c6475};
    assign in9260_2 = {c6476};
    Full_Adder FA_9260(s9260, c9260, in9260_1, in9260_2, c6474);
    wire[0:0] s9261, in9261_1, in9261_2;
    wire c9261;
    assign in9261_1 = {c6478};
    assign in9261_2 = {c6479};
    Full_Adder FA_9261(s9261, c9261, in9261_1, in9261_2, c6477);
    wire[0:0] s9262, in9262_1, in9262_2;
    wire c9262;
    assign in9262_1 = {c6481};
    assign in9262_2 = {c6482};
    Full_Adder FA_9262(s9262, c9262, in9262_1, in9262_2, c6480);
    wire[0:0] s9263, in9263_1, in9263_2;
    wire c9263;
    assign in9263_1 = {c6484};
    assign in9263_2 = {c6485};
    Full_Adder FA_9263(s9263, c9263, in9263_1, in9263_2, c6483);
    wire[0:0] s9264, in9264_1, in9264_2;
    wire c9264;
    assign in9264_1 = {c6487};
    assign in9264_2 = {c6488};
    Full_Adder FA_9264(s9264, c9264, in9264_1, in9264_2, c6486);
    wire[0:0] s9265, in9265_1, in9265_2;
    wire c9265;
    assign in9265_1 = {c6490};
    assign in9265_2 = {s6491[0]};
    Full_Adder FA_9265(s9265, c9265, in9265_1, in9265_2, c6489);
    wire[0:0] s9266, in9266_1, in9266_2;
    wire c9266;
    assign in9266_1 = {s6493[0]};
    assign in9266_2 = {s6494[0]};
    Full_Adder FA_9266(s9266, c9266, in9266_1, in9266_2, s6492[0]);
    wire[0:0] s9267, in9267_1, in9267_2;
    wire c9267;
    assign in9267_1 = {s6496[0]};
    assign in9267_2 = {s6497[0]};
    Full_Adder FA_9267(s9267, c9267, in9267_1, in9267_2, s6495[0]);
    wire[0:0] s9268, in9268_1, in9268_2;
    wire c9268;
    assign in9268_1 = {s6499[0]};
    assign in9268_2 = {s6500[0]};
    Full_Adder FA_9268(s9268, c9268, in9268_1, in9268_2, s6498[0]);
    wire[0:0] s9269, in9269_1, in9269_2;
    wire c9269;
    assign in9269_1 = {s6502[0]};
    assign in9269_2 = {s6503[0]};
    Full_Adder FA_9269(s9269, c9269, in9269_1, in9269_2, s6501[0]);
    wire[0:0] s9270, in9270_1, in9270_2;
    wire c9270;
    assign in9270_1 = {s6505[0]};
    assign in9270_2 = {s6506[0]};
    Full_Adder FA_9270(s9270, c9270, in9270_1, in9270_2, s6504[0]);
    wire[0:0] s9271, in9271_1, in9271_2;
    wire c9271;
    assign in9271_1 = {s6508[0]};
    assign in9271_2 = {s6509[0]};
    Full_Adder FA_9271(s9271, c9271, in9271_1, in9271_2, s6507[0]);
    wire[0:0] s9272, in9272_1, in9272_2;
    wire c9272;
    assign in9272_1 = {c6491};
    assign in9272_2 = {c6492};
    Full_Adder FA_9272(s9272, c9272, in9272_1, in9272_2, s3444[0]);
    wire[0:0] s9273, in9273_1, in9273_2;
    wire c9273;
    assign in9273_1 = {c6494};
    assign in9273_2 = {c6495};
    Full_Adder FA_9273(s9273, c9273, in9273_1, in9273_2, c6493);
    wire[0:0] s9274, in9274_1, in9274_2;
    wire c9274;
    assign in9274_1 = {c6497};
    assign in9274_2 = {c6498};
    Full_Adder FA_9274(s9274, c9274, in9274_1, in9274_2, c6496);
    wire[0:0] s9275, in9275_1, in9275_2;
    wire c9275;
    assign in9275_1 = {c6500};
    assign in9275_2 = {c6501};
    Full_Adder FA_9275(s9275, c9275, in9275_1, in9275_2, c6499);
    wire[0:0] s9276, in9276_1, in9276_2;
    wire c9276;
    assign in9276_1 = {c6503};
    assign in9276_2 = {c6504};
    Full_Adder FA_9276(s9276, c9276, in9276_1, in9276_2, c6502);
    wire[0:0] s9277, in9277_1, in9277_2;
    wire c9277;
    assign in9277_1 = {c6506};
    assign in9277_2 = {c6507};
    Full_Adder FA_9277(s9277, c9277, in9277_1, in9277_2, c6505);
    wire[0:0] s9278, in9278_1, in9278_2;
    wire c9278;
    assign in9278_1 = {c6509};
    assign in9278_2 = {s6510[0]};
    Full_Adder FA_9278(s9278, c9278, in9278_1, in9278_2, c6508);
    wire[0:0] s9279, in9279_1, in9279_2;
    wire c9279;
    assign in9279_1 = {s6512[0]};
    assign in9279_2 = {s6513[0]};
    Full_Adder FA_9279(s9279, c9279, in9279_1, in9279_2, s6511[0]);
    wire[0:0] s9280, in9280_1, in9280_2;
    wire c9280;
    assign in9280_1 = {s6515[0]};
    assign in9280_2 = {s6516[0]};
    Full_Adder FA_9280(s9280, c9280, in9280_1, in9280_2, s6514[0]);
    wire[0:0] s9281, in9281_1, in9281_2;
    wire c9281;
    assign in9281_1 = {s6518[0]};
    assign in9281_2 = {s6519[0]};
    Full_Adder FA_9281(s9281, c9281, in9281_1, in9281_2, s6517[0]);
    wire[0:0] s9282, in9282_1, in9282_2;
    wire c9282;
    assign in9282_1 = {s6521[0]};
    assign in9282_2 = {s6522[0]};
    Full_Adder FA_9282(s9282, c9282, in9282_1, in9282_2, s6520[0]);
    wire[0:0] s9283, in9283_1, in9283_2;
    wire c9283;
    assign in9283_1 = {s6524[0]};
    assign in9283_2 = {s6525[0]};
    Full_Adder FA_9283(s9283, c9283, in9283_1, in9283_2, s6523[0]);
    wire[0:0] s9284, in9284_1, in9284_2;
    wire c9284;
    assign in9284_1 = {s6527[0]};
    assign in9284_2 = {s6528[0]};
    Full_Adder FA_9284(s9284, c9284, in9284_1, in9284_2, s6526[0]);
    wire[0:0] s9285, in9285_1, in9285_2;
    wire c9285;
    assign in9285_1 = {c6510};
    assign in9285_2 = {c6511};
    Full_Adder FA_9285(s9285, c9285, in9285_1, in9285_2, s3472[0]);
    wire[0:0] s9286, in9286_1, in9286_2;
    wire c9286;
    assign in9286_1 = {c6513};
    assign in9286_2 = {c6514};
    Full_Adder FA_9286(s9286, c9286, in9286_1, in9286_2, c6512);
    wire[0:0] s9287, in9287_1, in9287_2;
    wire c9287;
    assign in9287_1 = {c6516};
    assign in9287_2 = {c6517};
    Full_Adder FA_9287(s9287, c9287, in9287_1, in9287_2, c6515);
    wire[0:0] s9288, in9288_1, in9288_2;
    wire c9288;
    assign in9288_1 = {c6519};
    assign in9288_2 = {c6520};
    Full_Adder FA_9288(s9288, c9288, in9288_1, in9288_2, c6518);
    wire[0:0] s9289, in9289_1, in9289_2;
    wire c9289;
    assign in9289_1 = {c6522};
    assign in9289_2 = {c6523};
    Full_Adder FA_9289(s9289, c9289, in9289_1, in9289_2, c6521);
    wire[0:0] s9290, in9290_1, in9290_2;
    wire c9290;
    assign in9290_1 = {c6525};
    assign in9290_2 = {c6526};
    Full_Adder FA_9290(s9290, c9290, in9290_1, in9290_2, c6524);
    wire[0:0] s9291, in9291_1, in9291_2;
    wire c9291;
    assign in9291_1 = {c6528};
    assign in9291_2 = {s6529[0]};
    Full_Adder FA_9291(s9291, c9291, in9291_1, in9291_2, c6527);
    wire[0:0] s9292, in9292_1, in9292_2;
    wire c9292;
    assign in9292_1 = {s6531[0]};
    assign in9292_2 = {s6532[0]};
    Full_Adder FA_9292(s9292, c9292, in9292_1, in9292_2, s6530[0]);
    wire[0:0] s9293, in9293_1, in9293_2;
    wire c9293;
    assign in9293_1 = {s6534[0]};
    assign in9293_2 = {s6535[0]};
    Full_Adder FA_9293(s9293, c9293, in9293_1, in9293_2, s6533[0]);
    wire[0:0] s9294, in9294_1, in9294_2;
    wire c9294;
    assign in9294_1 = {s6537[0]};
    assign in9294_2 = {s6538[0]};
    Full_Adder FA_9294(s9294, c9294, in9294_1, in9294_2, s6536[0]);
    wire[0:0] s9295, in9295_1, in9295_2;
    wire c9295;
    assign in9295_1 = {s6540[0]};
    assign in9295_2 = {s6541[0]};
    Full_Adder FA_9295(s9295, c9295, in9295_1, in9295_2, s6539[0]);
    wire[0:0] s9296, in9296_1, in9296_2;
    wire c9296;
    assign in9296_1 = {s6543[0]};
    assign in9296_2 = {s6544[0]};
    Full_Adder FA_9296(s9296, c9296, in9296_1, in9296_2, s6542[0]);
    wire[0:0] s9297, in9297_1, in9297_2;
    wire c9297;
    assign in9297_1 = {s6546[0]};
    assign in9297_2 = {s6547[0]};
    Full_Adder FA_9297(s9297, c9297, in9297_1, in9297_2, s6545[0]);
    wire[0:0] s9298, in9298_1, in9298_2;
    wire c9298;
    assign in9298_1 = {c6529};
    assign in9298_2 = {c6530};
    Full_Adder FA_9298(s9298, c9298, in9298_1, in9298_2, s3500[0]);
    wire[0:0] s9299, in9299_1, in9299_2;
    wire c9299;
    assign in9299_1 = {c6532};
    assign in9299_2 = {c6533};
    Full_Adder FA_9299(s9299, c9299, in9299_1, in9299_2, c6531);
    wire[0:0] s9300, in9300_1, in9300_2;
    wire c9300;
    assign in9300_1 = {c6535};
    assign in9300_2 = {c6536};
    Full_Adder FA_9300(s9300, c9300, in9300_1, in9300_2, c6534);
    wire[0:0] s9301, in9301_1, in9301_2;
    wire c9301;
    assign in9301_1 = {c6538};
    assign in9301_2 = {c6539};
    Full_Adder FA_9301(s9301, c9301, in9301_1, in9301_2, c6537);
    wire[0:0] s9302, in9302_1, in9302_2;
    wire c9302;
    assign in9302_1 = {c6541};
    assign in9302_2 = {c6542};
    Full_Adder FA_9302(s9302, c9302, in9302_1, in9302_2, c6540);
    wire[0:0] s9303, in9303_1, in9303_2;
    wire c9303;
    assign in9303_1 = {c6544};
    assign in9303_2 = {c6545};
    Full_Adder FA_9303(s9303, c9303, in9303_1, in9303_2, c6543);
    wire[0:0] s9304, in9304_1, in9304_2;
    wire c9304;
    assign in9304_1 = {c6547};
    assign in9304_2 = {s6548[0]};
    Full_Adder FA_9304(s9304, c9304, in9304_1, in9304_2, c6546);
    wire[0:0] s9305, in9305_1, in9305_2;
    wire c9305;
    assign in9305_1 = {s6550[0]};
    assign in9305_2 = {s6551[0]};
    Full_Adder FA_9305(s9305, c9305, in9305_1, in9305_2, s6549[0]);
    wire[0:0] s9306, in9306_1, in9306_2;
    wire c9306;
    assign in9306_1 = {s6553[0]};
    assign in9306_2 = {s6554[0]};
    Full_Adder FA_9306(s9306, c9306, in9306_1, in9306_2, s6552[0]);
    wire[0:0] s9307, in9307_1, in9307_2;
    wire c9307;
    assign in9307_1 = {s6556[0]};
    assign in9307_2 = {s6557[0]};
    Full_Adder FA_9307(s9307, c9307, in9307_1, in9307_2, s6555[0]);
    wire[0:0] s9308, in9308_1, in9308_2;
    wire c9308;
    assign in9308_1 = {s6559[0]};
    assign in9308_2 = {s6560[0]};
    Full_Adder FA_9308(s9308, c9308, in9308_1, in9308_2, s6558[0]);
    wire[0:0] s9309, in9309_1, in9309_2;
    wire c9309;
    assign in9309_1 = {s6562[0]};
    assign in9309_2 = {s6563[0]};
    Full_Adder FA_9309(s9309, c9309, in9309_1, in9309_2, s6561[0]);
    wire[0:0] s9310, in9310_1, in9310_2;
    wire c9310;
    assign in9310_1 = {s6565[0]};
    assign in9310_2 = {s6566[0]};
    Full_Adder FA_9310(s9310, c9310, in9310_1, in9310_2, s6564[0]);
    wire[0:0] s9311, in9311_1, in9311_2;
    wire c9311;
    assign in9311_1 = {c6548};
    assign in9311_2 = {c6549};
    Full_Adder FA_9311(s9311, c9311, in9311_1, in9311_2, s3528[0]);
    wire[0:0] s9312, in9312_1, in9312_2;
    wire c9312;
    assign in9312_1 = {c6551};
    assign in9312_2 = {c6552};
    Full_Adder FA_9312(s9312, c9312, in9312_1, in9312_2, c6550);
    wire[0:0] s9313, in9313_1, in9313_2;
    wire c9313;
    assign in9313_1 = {c6554};
    assign in9313_2 = {c6555};
    Full_Adder FA_9313(s9313, c9313, in9313_1, in9313_2, c6553);
    wire[0:0] s9314, in9314_1, in9314_2;
    wire c9314;
    assign in9314_1 = {c6557};
    assign in9314_2 = {c6558};
    Full_Adder FA_9314(s9314, c9314, in9314_1, in9314_2, c6556);
    wire[0:0] s9315, in9315_1, in9315_2;
    wire c9315;
    assign in9315_1 = {c6560};
    assign in9315_2 = {c6561};
    Full_Adder FA_9315(s9315, c9315, in9315_1, in9315_2, c6559);
    wire[0:0] s9316, in9316_1, in9316_2;
    wire c9316;
    assign in9316_1 = {c6563};
    assign in9316_2 = {c6564};
    Full_Adder FA_9316(s9316, c9316, in9316_1, in9316_2, c6562);
    wire[0:0] s9317, in9317_1, in9317_2;
    wire c9317;
    assign in9317_1 = {c6566};
    assign in9317_2 = {s6567[0]};
    Full_Adder FA_9317(s9317, c9317, in9317_1, in9317_2, c6565);
    wire[0:0] s9318, in9318_1, in9318_2;
    wire c9318;
    assign in9318_1 = {s6569[0]};
    assign in9318_2 = {s6570[0]};
    Full_Adder FA_9318(s9318, c9318, in9318_1, in9318_2, s6568[0]);
    wire[0:0] s9319, in9319_1, in9319_2;
    wire c9319;
    assign in9319_1 = {s6572[0]};
    assign in9319_2 = {s6573[0]};
    Full_Adder FA_9319(s9319, c9319, in9319_1, in9319_2, s6571[0]);
    wire[0:0] s9320, in9320_1, in9320_2;
    wire c9320;
    assign in9320_1 = {s6575[0]};
    assign in9320_2 = {s6576[0]};
    Full_Adder FA_9320(s9320, c9320, in9320_1, in9320_2, s6574[0]);
    wire[0:0] s9321, in9321_1, in9321_2;
    wire c9321;
    assign in9321_1 = {s6578[0]};
    assign in9321_2 = {s6579[0]};
    Full_Adder FA_9321(s9321, c9321, in9321_1, in9321_2, s6577[0]);
    wire[0:0] s9322, in9322_1, in9322_2;
    wire c9322;
    assign in9322_1 = {s6581[0]};
    assign in9322_2 = {s6582[0]};
    Full_Adder FA_9322(s9322, c9322, in9322_1, in9322_2, s6580[0]);
    wire[0:0] s9323, in9323_1, in9323_2;
    wire c9323;
    assign in9323_1 = {s6584[0]};
    assign in9323_2 = {s6585[0]};
    Full_Adder FA_9323(s9323, c9323, in9323_1, in9323_2, s6583[0]);
    wire[0:0] s9324, in9324_1, in9324_2;
    wire c9324;
    assign in9324_1 = {c6567};
    assign in9324_2 = {c6568};
    Full_Adder FA_9324(s9324, c9324, in9324_1, in9324_2, s3556[0]);
    wire[0:0] s9325, in9325_1, in9325_2;
    wire c9325;
    assign in9325_1 = {c6570};
    assign in9325_2 = {c6571};
    Full_Adder FA_9325(s9325, c9325, in9325_1, in9325_2, c6569);
    wire[0:0] s9326, in9326_1, in9326_2;
    wire c9326;
    assign in9326_1 = {c6573};
    assign in9326_2 = {c6574};
    Full_Adder FA_9326(s9326, c9326, in9326_1, in9326_2, c6572);
    wire[0:0] s9327, in9327_1, in9327_2;
    wire c9327;
    assign in9327_1 = {c6576};
    assign in9327_2 = {c6577};
    Full_Adder FA_9327(s9327, c9327, in9327_1, in9327_2, c6575);
    wire[0:0] s9328, in9328_1, in9328_2;
    wire c9328;
    assign in9328_1 = {c6579};
    assign in9328_2 = {c6580};
    Full_Adder FA_9328(s9328, c9328, in9328_1, in9328_2, c6578);
    wire[0:0] s9329, in9329_1, in9329_2;
    wire c9329;
    assign in9329_1 = {c6582};
    assign in9329_2 = {c6583};
    Full_Adder FA_9329(s9329, c9329, in9329_1, in9329_2, c6581);
    wire[0:0] s9330, in9330_1, in9330_2;
    wire c9330;
    assign in9330_1 = {c6585};
    assign in9330_2 = {s6586[0]};
    Full_Adder FA_9330(s9330, c9330, in9330_1, in9330_2, c6584);
    wire[0:0] s9331, in9331_1, in9331_2;
    wire c9331;
    assign in9331_1 = {s6588[0]};
    assign in9331_2 = {s6589[0]};
    Full_Adder FA_9331(s9331, c9331, in9331_1, in9331_2, s6587[0]);
    wire[0:0] s9332, in9332_1, in9332_2;
    wire c9332;
    assign in9332_1 = {s6591[0]};
    assign in9332_2 = {s6592[0]};
    Full_Adder FA_9332(s9332, c9332, in9332_1, in9332_2, s6590[0]);
    wire[0:0] s9333, in9333_1, in9333_2;
    wire c9333;
    assign in9333_1 = {s6594[0]};
    assign in9333_2 = {s6595[0]};
    Full_Adder FA_9333(s9333, c9333, in9333_1, in9333_2, s6593[0]);
    wire[0:0] s9334, in9334_1, in9334_2;
    wire c9334;
    assign in9334_1 = {s6597[0]};
    assign in9334_2 = {s6598[0]};
    Full_Adder FA_9334(s9334, c9334, in9334_1, in9334_2, s6596[0]);
    wire[0:0] s9335, in9335_1, in9335_2;
    wire c9335;
    assign in9335_1 = {s6600[0]};
    assign in9335_2 = {s6601[0]};
    Full_Adder FA_9335(s9335, c9335, in9335_1, in9335_2, s6599[0]);
    wire[0:0] s9336, in9336_1, in9336_2;
    wire c9336;
    assign in9336_1 = {s6603[0]};
    assign in9336_2 = {s6604[0]};
    Full_Adder FA_9336(s9336, c9336, in9336_1, in9336_2, s6602[0]);
    wire[0:0] s9337, in9337_1, in9337_2;
    wire c9337;
    assign in9337_1 = {c6586};
    assign in9337_2 = {c6587};
    Full_Adder FA_9337(s9337, c9337, in9337_1, in9337_2, s3584[0]);
    wire[0:0] s9338, in9338_1, in9338_2;
    wire c9338;
    assign in9338_1 = {c6589};
    assign in9338_2 = {c6590};
    Full_Adder FA_9338(s9338, c9338, in9338_1, in9338_2, c6588);
    wire[0:0] s9339, in9339_1, in9339_2;
    wire c9339;
    assign in9339_1 = {c6592};
    assign in9339_2 = {c6593};
    Full_Adder FA_9339(s9339, c9339, in9339_1, in9339_2, c6591);
    wire[0:0] s9340, in9340_1, in9340_2;
    wire c9340;
    assign in9340_1 = {c6595};
    assign in9340_2 = {c6596};
    Full_Adder FA_9340(s9340, c9340, in9340_1, in9340_2, c6594);
    wire[0:0] s9341, in9341_1, in9341_2;
    wire c9341;
    assign in9341_1 = {c6598};
    assign in9341_2 = {c6599};
    Full_Adder FA_9341(s9341, c9341, in9341_1, in9341_2, c6597);
    wire[0:0] s9342, in9342_1, in9342_2;
    wire c9342;
    assign in9342_1 = {c6601};
    assign in9342_2 = {c6602};
    Full_Adder FA_9342(s9342, c9342, in9342_1, in9342_2, c6600);
    wire[0:0] s9343, in9343_1, in9343_2;
    wire c9343;
    assign in9343_1 = {c6604};
    assign in9343_2 = {s6605[0]};
    Full_Adder FA_9343(s9343, c9343, in9343_1, in9343_2, c6603);
    wire[0:0] s9344, in9344_1, in9344_2;
    wire c9344;
    assign in9344_1 = {s6607[0]};
    assign in9344_2 = {s6608[0]};
    Full_Adder FA_9344(s9344, c9344, in9344_1, in9344_2, s6606[0]);
    wire[0:0] s9345, in9345_1, in9345_2;
    wire c9345;
    assign in9345_1 = {s6610[0]};
    assign in9345_2 = {s6611[0]};
    Full_Adder FA_9345(s9345, c9345, in9345_1, in9345_2, s6609[0]);
    wire[0:0] s9346, in9346_1, in9346_2;
    wire c9346;
    assign in9346_1 = {s6613[0]};
    assign in9346_2 = {s6614[0]};
    Full_Adder FA_9346(s9346, c9346, in9346_1, in9346_2, s6612[0]);
    wire[0:0] s9347, in9347_1, in9347_2;
    wire c9347;
    assign in9347_1 = {s6616[0]};
    assign in9347_2 = {s6617[0]};
    Full_Adder FA_9347(s9347, c9347, in9347_1, in9347_2, s6615[0]);
    wire[0:0] s9348, in9348_1, in9348_2;
    wire c9348;
    assign in9348_1 = {s6619[0]};
    assign in9348_2 = {s6620[0]};
    Full_Adder FA_9348(s9348, c9348, in9348_1, in9348_2, s6618[0]);
    wire[0:0] s9349, in9349_1, in9349_2;
    wire c9349;
    assign in9349_1 = {s6622[0]};
    assign in9349_2 = {s6623[0]};
    Full_Adder FA_9349(s9349, c9349, in9349_1, in9349_2, s6621[0]);
    wire[0:0] s9350, in9350_1, in9350_2;
    wire c9350;
    assign in9350_1 = {c6605};
    assign in9350_2 = {c6606};
    Full_Adder FA_9350(s9350, c9350, in9350_1, in9350_2, s3612[0]);
    wire[0:0] s9351, in9351_1, in9351_2;
    wire c9351;
    assign in9351_1 = {c6608};
    assign in9351_2 = {c6609};
    Full_Adder FA_9351(s9351, c9351, in9351_1, in9351_2, c6607);
    wire[0:0] s9352, in9352_1, in9352_2;
    wire c9352;
    assign in9352_1 = {c6611};
    assign in9352_2 = {c6612};
    Full_Adder FA_9352(s9352, c9352, in9352_1, in9352_2, c6610);
    wire[0:0] s9353, in9353_1, in9353_2;
    wire c9353;
    assign in9353_1 = {c6614};
    assign in9353_2 = {c6615};
    Full_Adder FA_9353(s9353, c9353, in9353_1, in9353_2, c6613);
    wire[0:0] s9354, in9354_1, in9354_2;
    wire c9354;
    assign in9354_1 = {c6617};
    assign in9354_2 = {c6618};
    Full_Adder FA_9354(s9354, c9354, in9354_1, in9354_2, c6616);
    wire[0:0] s9355, in9355_1, in9355_2;
    wire c9355;
    assign in9355_1 = {c6620};
    assign in9355_2 = {c6621};
    Full_Adder FA_9355(s9355, c9355, in9355_1, in9355_2, c6619);
    wire[0:0] s9356, in9356_1, in9356_2;
    wire c9356;
    assign in9356_1 = {c6623};
    assign in9356_2 = {s6624[0]};
    Full_Adder FA_9356(s9356, c9356, in9356_1, in9356_2, c6622);
    wire[0:0] s9357, in9357_1, in9357_2;
    wire c9357;
    assign in9357_1 = {s6626[0]};
    assign in9357_2 = {s6627[0]};
    Full_Adder FA_9357(s9357, c9357, in9357_1, in9357_2, s6625[0]);
    wire[0:0] s9358, in9358_1, in9358_2;
    wire c9358;
    assign in9358_1 = {s6629[0]};
    assign in9358_2 = {s6630[0]};
    Full_Adder FA_9358(s9358, c9358, in9358_1, in9358_2, s6628[0]);
    wire[0:0] s9359, in9359_1, in9359_2;
    wire c9359;
    assign in9359_1 = {s6632[0]};
    assign in9359_2 = {s6633[0]};
    Full_Adder FA_9359(s9359, c9359, in9359_1, in9359_2, s6631[0]);
    wire[0:0] s9360, in9360_1, in9360_2;
    wire c9360;
    assign in9360_1 = {s6635[0]};
    assign in9360_2 = {s6636[0]};
    Full_Adder FA_9360(s9360, c9360, in9360_1, in9360_2, s6634[0]);
    wire[0:0] s9361, in9361_1, in9361_2;
    wire c9361;
    assign in9361_1 = {s6638[0]};
    assign in9361_2 = {s6639[0]};
    Full_Adder FA_9361(s9361, c9361, in9361_1, in9361_2, s6637[0]);
    wire[0:0] s9362, in9362_1, in9362_2;
    wire c9362;
    assign in9362_1 = {s6641[0]};
    assign in9362_2 = {s6642[0]};
    Full_Adder FA_9362(s9362, c9362, in9362_1, in9362_2, s6640[0]);
    wire[0:0] s9363, in9363_1, in9363_2;
    wire c9363;
    assign in9363_1 = {c6624};
    assign in9363_2 = {c6625};
    Full_Adder FA_9363(s9363, c9363, in9363_1, in9363_2, s3640[0]);
    wire[0:0] s9364, in9364_1, in9364_2;
    wire c9364;
    assign in9364_1 = {c6627};
    assign in9364_2 = {c6628};
    Full_Adder FA_9364(s9364, c9364, in9364_1, in9364_2, c6626);
    wire[0:0] s9365, in9365_1, in9365_2;
    wire c9365;
    assign in9365_1 = {c6630};
    assign in9365_2 = {c6631};
    Full_Adder FA_9365(s9365, c9365, in9365_1, in9365_2, c6629);
    wire[0:0] s9366, in9366_1, in9366_2;
    wire c9366;
    assign in9366_1 = {c6633};
    assign in9366_2 = {c6634};
    Full_Adder FA_9366(s9366, c9366, in9366_1, in9366_2, c6632);
    wire[0:0] s9367, in9367_1, in9367_2;
    wire c9367;
    assign in9367_1 = {c6636};
    assign in9367_2 = {c6637};
    Full_Adder FA_9367(s9367, c9367, in9367_1, in9367_2, c6635);
    wire[0:0] s9368, in9368_1, in9368_2;
    wire c9368;
    assign in9368_1 = {c6639};
    assign in9368_2 = {c6640};
    Full_Adder FA_9368(s9368, c9368, in9368_1, in9368_2, c6638);
    wire[0:0] s9369, in9369_1, in9369_2;
    wire c9369;
    assign in9369_1 = {c6642};
    assign in9369_2 = {s6643[0]};
    Full_Adder FA_9369(s9369, c9369, in9369_1, in9369_2, c6641);
    wire[0:0] s9370, in9370_1, in9370_2;
    wire c9370;
    assign in9370_1 = {s6645[0]};
    assign in9370_2 = {s6646[0]};
    Full_Adder FA_9370(s9370, c9370, in9370_1, in9370_2, s6644[0]);
    wire[0:0] s9371, in9371_1, in9371_2;
    wire c9371;
    assign in9371_1 = {s6648[0]};
    assign in9371_2 = {s6649[0]};
    Full_Adder FA_9371(s9371, c9371, in9371_1, in9371_2, s6647[0]);
    wire[0:0] s9372, in9372_1, in9372_2;
    wire c9372;
    assign in9372_1 = {s6651[0]};
    assign in9372_2 = {s6652[0]};
    Full_Adder FA_9372(s9372, c9372, in9372_1, in9372_2, s6650[0]);
    wire[0:0] s9373, in9373_1, in9373_2;
    wire c9373;
    assign in9373_1 = {s6654[0]};
    assign in9373_2 = {s6655[0]};
    Full_Adder FA_9373(s9373, c9373, in9373_1, in9373_2, s6653[0]);
    wire[0:0] s9374, in9374_1, in9374_2;
    wire c9374;
    assign in9374_1 = {s6657[0]};
    assign in9374_2 = {s6658[0]};
    Full_Adder FA_9374(s9374, c9374, in9374_1, in9374_2, s6656[0]);
    wire[0:0] s9375, in9375_1, in9375_2;
    wire c9375;
    assign in9375_1 = {s6660[0]};
    assign in9375_2 = {s6661[0]};
    Full_Adder FA_9375(s9375, c9375, in9375_1, in9375_2, s6659[0]);
    wire[0:0] s9376, in9376_1, in9376_2;
    wire c9376;
    assign in9376_1 = {c6643};
    assign in9376_2 = {c6644};
    Full_Adder FA_9376(s9376, c9376, in9376_1, in9376_2, s3668[0]);
    wire[0:0] s9377, in9377_1, in9377_2;
    wire c9377;
    assign in9377_1 = {c6646};
    assign in9377_2 = {c6647};
    Full_Adder FA_9377(s9377, c9377, in9377_1, in9377_2, c6645);
    wire[0:0] s9378, in9378_1, in9378_2;
    wire c9378;
    assign in9378_1 = {c6649};
    assign in9378_2 = {c6650};
    Full_Adder FA_9378(s9378, c9378, in9378_1, in9378_2, c6648);
    wire[0:0] s9379, in9379_1, in9379_2;
    wire c9379;
    assign in9379_1 = {c6652};
    assign in9379_2 = {c6653};
    Full_Adder FA_9379(s9379, c9379, in9379_1, in9379_2, c6651);
    wire[0:0] s9380, in9380_1, in9380_2;
    wire c9380;
    assign in9380_1 = {c6655};
    assign in9380_2 = {c6656};
    Full_Adder FA_9380(s9380, c9380, in9380_1, in9380_2, c6654);
    wire[0:0] s9381, in9381_1, in9381_2;
    wire c9381;
    assign in9381_1 = {c6658};
    assign in9381_2 = {c6659};
    Full_Adder FA_9381(s9381, c9381, in9381_1, in9381_2, c6657);
    wire[0:0] s9382, in9382_1, in9382_2;
    wire c9382;
    assign in9382_1 = {c6661};
    assign in9382_2 = {s6662[0]};
    Full_Adder FA_9382(s9382, c9382, in9382_1, in9382_2, c6660);
    wire[0:0] s9383, in9383_1, in9383_2;
    wire c9383;
    assign in9383_1 = {s6664[0]};
    assign in9383_2 = {s6665[0]};
    Full_Adder FA_9383(s9383, c9383, in9383_1, in9383_2, s6663[0]);
    wire[0:0] s9384, in9384_1, in9384_2;
    wire c9384;
    assign in9384_1 = {s6667[0]};
    assign in9384_2 = {s6668[0]};
    Full_Adder FA_9384(s9384, c9384, in9384_1, in9384_2, s6666[0]);
    wire[0:0] s9385, in9385_1, in9385_2;
    wire c9385;
    assign in9385_1 = {s6670[0]};
    assign in9385_2 = {s6671[0]};
    Full_Adder FA_9385(s9385, c9385, in9385_1, in9385_2, s6669[0]);
    wire[0:0] s9386, in9386_1, in9386_2;
    wire c9386;
    assign in9386_1 = {s6673[0]};
    assign in9386_2 = {s6674[0]};
    Full_Adder FA_9386(s9386, c9386, in9386_1, in9386_2, s6672[0]);
    wire[0:0] s9387, in9387_1, in9387_2;
    wire c9387;
    assign in9387_1 = {s6676[0]};
    assign in9387_2 = {s6677[0]};
    Full_Adder FA_9387(s9387, c9387, in9387_1, in9387_2, s6675[0]);
    wire[0:0] s9388, in9388_1, in9388_2;
    wire c9388;
    assign in9388_1 = {s6679[0]};
    assign in9388_2 = {s6680[0]};
    Full_Adder FA_9388(s9388, c9388, in9388_1, in9388_2, s6678[0]);
    wire[0:0] s9389, in9389_1, in9389_2;
    wire c9389;
    assign in9389_1 = {c6662};
    assign in9389_2 = {c6663};
    Full_Adder FA_9389(s9389, c9389, in9389_1, in9389_2, s3696[0]);
    wire[0:0] s9390, in9390_1, in9390_2;
    wire c9390;
    assign in9390_1 = {c6665};
    assign in9390_2 = {c6666};
    Full_Adder FA_9390(s9390, c9390, in9390_1, in9390_2, c6664);
    wire[0:0] s9391, in9391_1, in9391_2;
    wire c9391;
    assign in9391_1 = {c6668};
    assign in9391_2 = {c6669};
    Full_Adder FA_9391(s9391, c9391, in9391_1, in9391_2, c6667);
    wire[0:0] s9392, in9392_1, in9392_2;
    wire c9392;
    assign in9392_1 = {c6671};
    assign in9392_2 = {c6672};
    Full_Adder FA_9392(s9392, c9392, in9392_1, in9392_2, c6670);
    wire[0:0] s9393, in9393_1, in9393_2;
    wire c9393;
    assign in9393_1 = {c6674};
    assign in9393_2 = {c6675};
    Full_Adder FA_9393(s9393, c9393, in9393_1, in9393_2, c6673);
    wire[0:0] s9394, in9394_1, in9394_2;
    wire c9394;
    assign in9394_1 = {c6677};
    assign in9394_2 = {c6678};
    Full_Adder FA_9394(s9394, c9394, in9394_1, in9394_2, c6676);
    wire[0:0] s9395, in9395_1, in9395_2;
    wire c9395;
    assign in9395_1 = {c6680};
    assign in9395_2 = {s6681[0]};
    Full_Adder FA_9395(s9395, c9395, in9395_1, in9395_2, c6679);
    wire[0:0] s9396, in9396_1, in9396_2;
    wire c9396;
    assign in9396_1 = {s6683[0]};
    assign in9396_2 = {s6684[0]};
    Full_Adder FA_9396(s9396, c9396, in9396_1, in9396_2, s6682[0]);
    wire[0:0] s9397, in9397_1, in9397_2;
    wire c9397;
    assign in9397_1 = {s6686[0]};
    assign in9397_2 = {s6687[0]};
    Full_Adder FA_9397(s9397, c9397, in9397_1, in9397_2, s6685[0]);
    wire[0:0] s9398, in9398_1, in9398_2;
    wire c9398;
    assign in9398_1 = {s6689[0]};
    assign in9398_2 = {s6690[0]};
    Full_Adder FA_9398(s9398, c9398, in9398_1, in9398_2, s6688[0]);
    wire[0:0] s9399, in9399_1, in9399_2;
    wire c9399;
    assign in9399_1 = {s6692[0]};
    assign in9399_2 = {s6693[0]};
    Full_Adder FA_9399(s9399, c9399, in9399_1, in9399_2, s6691[0]);
    wire[0:0] s9400, in9400_1, in9400_2;
    wire c9400;
    assign in9400_1 = {s6695[0]};
    assign in9400_2 = {s6696[0]};
    Full_Adder FA_9400(s9400, c9400, in9400_1, in9400_2, s6694[0]);
    wire[0:0] s9401, in9401_1, in9401_2;
    wire c9401;
    assign in9401_1 = {s6698[0]};
    assign in9401_2 = {s6699[0]};
    Full_Adder FA_9401(s9401, c9401, in9401_1, in9401_2, s6697[0]);
    wire[0:0] s9402, in9402_1, in9402_2;
    wire c9402;
    assign in9402_1 = {c6681};
    assign in9402_2 = {c6682};
    Full_Adder FA_9402(s9402, c9402, in9402_1, in9402_2, s3724[0]);
    wire[0:0] s9403, in9403_1, in9403_2;
    wire c9403;
    assign in9403_1 = {c6684};
    assign in9403_2 = {c6685};
    Full_Adder FA_9403(s9403, c9403, in9403_1, in9403_2, c6683);
    wire[0:0] s9404, in9404_1, in9404_2;
    wire c9404;
    assign in9404_1 = {c6687};
    assign in9404_2 = {c6688};
    Full_Adder FA_9404(s9404, c9404, in9404_1, in9404_2, c6686);
    wire[0:0] s9405, in9405_1, in9405_2;
    wire c9405;
    assign in9405_1 = {c6690};
    assign in9405_2 = {c6691};
    Full_Adder FA_9405(s9405, c9405, in9405_1, in9405_2, c6689);
    wire[0:0] s9406, in9406_1, in9406_2;
    wire c9406;
    assign in9406_1 = {c6693};
    assign in9406_2 = {c6694};
    Full_Adder FA_9406(s9406, c9406, in9406_1, in9406_2, c6692);
    wire[0:0] s9407, in9407_1, in9407_2;
    wire c9407;
    assign in9407_1 = {c6696};
    assign in9407_2 = {c6697};
    Full_Adder FA_9407(s9407, c9407, in9407_1, in9407_2, c6695);
    wire[0:0] s9408, in9408_1, in9408_2;
    wire c9408;
    assign in9408_1 = {c6699};
    assign in9408_2 = {s6700[0]};
    Full_Adder FA_9408(s9408, c9408, in9408_1, in9408_2, c6698);
    wire[0:0] s9409, in9409_1, in9409_2;
    wire c9409;
    assign in9409_1 = {s6702[0]};
    assign in9409_2 = {s6703[0]};
    Full_Adder FA_9409(s9409, c9409, in9409_1, in9409_2, s6701[0]);
    wire[0:0] s9410, in9410_1, in9410_2;
    wire c9410;
    assign in9410_1 = {s6705[0]};
    assign in9410_2 = {s6706[0]};
    Full_Adder FA_9410(s9410, c9410, in9410_1, in9410_2, s6704[0]);
    wire[0:0] s9411, in9411_1, in9411_2;
    wire c9411;
    assign in9411_1 = {s6708[0]};
    assign in9411_2 = {s6709[0]};
    Full_Adder FA_9411(s9411, c9411, in9411_1, in9411_2, s6707[0]);
    wire[0:0] s9412, in9412_1, in9412_2;
    wire c9412;
    assign in9412_1 = {s6711[0]};
    assign in9412_2 = {s6712[0]};
    Full_Adder FA_9412(s9412, c9412, in9412_1, in9412_2, s6710[0]);
    wire[0:0] s9413, in9413_1, in9413_2;
    wire c9413;
    assign in9413_1 = {s6714[0]};
    assign in9413_2 = {s6715[0]};
    Full_Adder FA_9413(s9413, c9413, in9413_1, in9413_2, s6713[0]);
    wire[0:0] s9414, in9414_1, in9414_2;
    wire c9414;
    assign in9414_1 = {s6717[0]};
    assign in9414_2 = {s6718[0]};
    Full_Adder FA_9414(s9414, c9414, in9414_1, in9414_2, s6716[0]);
    wire[0:0] s9415, in9415_1, in9415_2;
    wire c9415;
    assign in9415_1 = {c6700};
    assign in9415_2 = {c6701};
    Full_Adder FA_9415(s9415, c9415, in9415_1, in9415_2, s3752[0]);
    wire[0:0] s9416, in9416_1, in9416_2;
    wire c9416;
    assign in9416_1 = {c6703};
    assign in9416_2 = {c6704};
    Full_Adder FA_9416(s9416, c9416, in9416_1, in9416_2, c6702);
    wire[0:0] s9417, in9417_1, in9417_2;
    wire c9417;
    assign in9417_1 = {c6706};
    assign in9417_2 = {c6707};
    Full_Adder FA_9417(s9417, c9417, in9417_1, in9417_2, c6705);
    wire[0:0] s9418, in9418_1, in9418_2;
    wire c9418;
    assign in9418_1 = {c6709};
    assign in9418_2 = {c6710};
    Full_Adder FA_9418(s9418, c9418, in9418_1, in9418_2, c6708);
    wire[0:0] s9419, in9419_1, in9419_2;
    wire c9419;
    assign in9419_1 = {c6712};
    assign in9419_2 = {c6713};
    Full_Adder FA_9419(s9419, c9419, in9419_1, in9419_2, c6711);
    wire[0:0] s9420, in9420_1, in9420_2;
    wire c9420;
    assign in9420_1 = {c6715};
    assign in9420_2 = {c6716};
    Full_Adder FA_9420(s9420, c9420, in9420_1, in9420_2, c6714);
    wire[0:0] s9421, in9421_1, in9421_2;
    wire c9421;
    assign in9421_1 = {c6718};
    assign in9421_2 = {s6719[0]};
    Full_Adder FA_9421(s9421, c9421, in9421_1, in9421_2, c6717);
    wire[0:0] s9422, in9422_1, in9422_2;
    wire c9422;
    assign in9422_1 = {s6721[0]};
    assign in9422_2 = {s6722[0]};
    Full_Adder FA_9422(s9422, c9422, in9422_1, in9422_2, s6720[0]);
    wire[0:0] s9423, in9423_1, in9423_2;
    wire c9423;
    assign in9423_1 = {s6724[0]};
    assign in9423_2 = {s6725[0]};
    Full_Adder FA_9423(s9423, c9423, in9423_1, in9423_2, s6723[0]);
    wire[0:0] s9424, in9424_1, in9424_2;
    wire c9424;
    assign in9424_1 = {s6727[0]};
    assign in9424_2 = {s6728[0]};
    Full_Adder FA_9424(s9424, c9424, in9424_1, in9424_2, s6726[0]);
    wire[0:0] s9425, in9425_1, in9425_2;
    wire c9425;
    assign in9425_1 = {s6730[0]};
    assign in9425_2 = {s6731[0]};
    Full_Adder FA_9425(s9425, c9425, in9425_1, in9425_2, s6729[0]);
    wire[0:0] s9426, in9426_1, in9426_2;
    wire c9426;
    assign in9426_1 = {s6733[0]};
    assign in9426_2 = {s6734[0]};
    Full_Adder FA_9426(s9426, c9426, in9426_1, in9426_2, s6732[0]);
    wire[0:0] s9427, in9427_1, in9427_2;
    wire c9427;
    assign in9427_1 = {s6736[0]};
    assign in9427_2 = {s6737[0]};
    Full_Adder FA_9427(s9427, c9427, in9427_1, in9427_2, s6735[0]);
    wire[0:0] s9428, in9428_1, in9428_2;
    wire c9428;
    assign in9428_1 = {c6719};
    assign in9428_2 = {c6720};
    Full_Adder FA_9428(s9428, c9428, in9428_1, in9428_2, s3780[0]);
    wire[0:0] s9429, in9429_1, in9429_2;
    wire c9429;
    assign in9429_1 = {c6722};
    assign in9429_2 = {c6723};
    Full_Adder FA_9429(s9429, c9429, in9429_1, in9429_2, c6721);
    wire[0:0] s9430, in9430_1, in9430_2;
    wire c9430;
    assign in9430_1 = {c6725};
    assign in9430_2 = {c6726};
    Full_Adder FA_9430(s9430, c9430, in9430_1, in9430_2, c6724);
    wire[0:0] s9431, in9431_1, in9431_2;
    wire c9431;
    assign in9431_1 = {c6728};
    assign in9431_2 = {c6729};
    Full_Adder FA_9431(s9431, c9431, in9431_1, in9431_2, c6727);
    wire[0:0] s9432, in9432_1, in9432_2;
    wire c9432;
    assign in9432_1 = {c6731};
    assign in9432_2 = {c6732};
    Full_Adder FA_9432(s9432, c9432, in9432_1, in9432_2, c6730);
    wire[0:0] s9433, in9433_1, in9433_2;
    wire c9433;
    assign in9433_1 = {c6734};
    assign in9433_2 = {c6735};
    Full_Adder FA_9433(s9433, c9433, in9433_1, in9433_2, c6733);
    wire[0:0] s9434, in9434_1, in9434_2;
    wire c9434;
    assign in9434_1 = {c6737};
    assign in9434_2 = {s6738[0]};
    Full_Adder FA_9434(s9434, c9434, in9434_1, in9434_2, c6736);
    wire[0:0] s9435, in9435_1, in9435_2;
    wire c9435;
    assign in9435_1 = {s6740[0]};
    assign in9435_2 = {s6741[0]};
    Full_Adder FA_9435(s9435, c9435, in9435_1, in9435_2, s6739[0]);
    wire[0:0] s9436, in9436_1, in9436_2;
    wire c9436;
    assign in9436_1 = {s6743[0]};
    assign in9436_2 = {s6744[0]};
    Full_Adder FA_9436(s9436, c9436, in9436_1, in9436_2, s6742[0]);
    wire[0:0] s9437, in9437_1, in9437_2;
    wire c9437;
    assign in9437_1 = {s6746[0]};
    assign in9437_2 = {s6747[0]};
    Full_Adder FA_9437(s9437, c9437, in9437_1, in9437_2, s6745[0]);
    wire[0:0] s9438, in9438_1, in9438_2;
    wire c9438;
    assign in9438_1 = {s6749[0]};
    assign in9438_2 = {s6750[0]};
    Full_Adder FA_9438(s9438, c9438, in9438_1, in9438_2, s6748[0]);
    wire[0:0] s9439, in9439_1, in9439_2;
    wire c9439;
    assign in9439_1 = {s6752[0]};
    assign in9439_2 = {s6753[0]};
    Full_Adder FA_9439(s9439, c9439, in9439_1, in9439_2, s6751[0]);
    wire[0:0] s9440, in9440_1, in9440_2;
    wire c9440;
    assign in9440_1 = {s6755[0]};
    assign in9440_2 = {s6756[0]};
    Full_Adder FA_9440(s9440, c9440, in9440_1, in9440_2, s6754[0]);
    wire[0:0] s9441, in9441_1, in9441_2;
    wire c9441;
    assign in9441_1 = {c6738};
    assign in9441_2 = {c6739};
    Full_Adder FA_9441(s9441, c9441, in9441_1, in9441_2, s3808[0]);
    wire[0:0] s9442, in9442_1, in9442_2;
    wire c9442;
    assign in9442_1 = {c6741};
    assign in9442_2 = {c6742};
    Full_Adder FA_9442(s9442, c9442, in9442_1, in9442_2, c6740);
    wire[0:0] s9443, in9443_1, in9443_2;
    wire c9443;
    assign in9443_1 = {c6744};
    assign in9443_2 = {c6745};
    Full_Adder FA_9443(s9443, c9443, in9443_1, in9443_2, c6743);
    wire[0:0] s9444, in9444_1, in9444_2;
    wire c9444;
    assign in9444_1 = {c6747};
    assign in9444_2 = {c6748};
    Full_Adder FA_9444(s9444, c9444, in9444_1, in9444_2, c6746);
    wire[0:0] s9445, in9445_1, in9445_2;
    wire c9445;
    assign in9445_1 = {c6750};
    assign in9445_2 = {c6751};
    Full_Adder FA_9445(s9445, c9445, in9445_1, in9445_2, c6749);
    wire[0:0] s9446, in9446_1, in9446_2;
    wire c9446;
    assign in9446_1 = {c6753};
    assign in9446_2 = {c6754};
    Full_Adder FA_9446(s9446, c9446, in9446_1, in9446_2, c6752);
    wire[0:0] s9447, in9447_1, in9447_2;
    wire c9447;
    assign in9447_1 = {c6756};
    assign in9447_2 = {s6757[0]};
    Full_Adder FA_9447(s9447, c9447, in9447_1, in9447_2, c6755);
    wire[0:0] s9448, in9448_1, in9448_2;
    wire c9448;
    assign in9448_1 = {s6759[0]};
    assign in9448_2 = {s6760[0]};
    Full_Adder FA_9448(s9448, c9448, in9448_1, in9448_2, s6758[0]);
    wire[0:0] s9449, in9449_1, in9449_2;
    wire c9449;
    assign in9449_1 = {s6762[0]};
    assign in9449_2 = {s6763[0]};
    Full_Adder FA_9449(s9449, c9449, in9449_1, in9449_2, s6761[0]);
    wire[0:0] s9450, in9450_1, in9450_2;
    wire c9450;
    assign in9450_1 = {s6765[0]};
    assign in9450_2 = {s6766[0]};
    Full_Adder FA_9450(s9450, c9450, in9450_1, in9450_2, s6764[0]);
    wire[0:0] s9451, in9451_1, in9451_2;
    wire c9451;
    assign in9451_1 = {s6768[0]};
    assign in9451_2 = {s6769[0]};
    Full_Adder FA_9451(s9451, c9451, in9451_1, in9451_2, s6767[0]);
    wire[0:0] s9452, in9452_1, in9452_2;
    wire c9452;
    assign in9452_1 = {s6771[0]};
    assign in9452_2 = {s6772[0]};
    Full_Adder FA_9452(s9452, c9452, in9452_1, in9452_2, s6770[0]);
    wire[0:0] s9453, in9453_1, in9453_2;
    wire c9453;
    assign in9453_1 = {s6774[0]};
    assign in9453_2 = {s6775[0]};
    Full_Adder FA_9453(s9453, c9453, in9453_1, in9453_2, s6773[0]);
    wire[0:0] s9454, in9454_1, in9454_2;
    wire c9454;
    assign in9454_1 = {c6757};
    assign in9454_2 = {c6758};
    Full_Adder FA_9454(s9454, c9454, in9454_1, in9454_2, s3836[0]);
    wire[0:0] s9455, in9455_1, in9455_2;
    wire c9455;
    assign in9455_1 = {c6760};
    assign in9455_2 = {c6761};
    Full_Adder FA_9455(s9455, c9455, in9455_1, in9455_2, c6759);
    wire[0:0] s9456, in9456_1, in9456_2;
    wire c9456;
    assign in9456_1 = {c6763};
    assign in9456_2 = {c6764};
    Full_Adder FA_9456(s9456, c9456, in9456_1, in9456_2, c6762);
    wire[0:0] s9457, in9457_1, in9457_2;
    wire c9457;
    assign in9457_1 = {c6766};
    assign in9457_2 = {c6767};
    Full_Adder FA_9457(s9457, c9457, in9457_1, in9457_2, c6765);
    wire[0:0] s9458, in9458_1, in9458_2;
    wire c9458;
    assign in9458_1 = {c6769};
    assign in9458_2 = {c6770};
    Full_Adder FA_9458(s9458, c9458, in9458_1, in9458_2, c6768);
    wire[0:0] s9459, in9459_1, in9459_2;
    wire c9459;
    assign in9459_1 = {c6772};
    assign in9459_2 = {c6773};
    Full_Adder FA_9459(s9459, c9459, in9459_1, in9459_2, c6771);
    wire[0:0] s9460, in9460_1, in9460_2;
    wire c9460;
    assign in9460_1 = {c6775};
    assign in9460_2 = {s6776[0]};
    Full_Adder FA_9460(s9460, c9460, in9460_1, in9460_2, c6774);
    wire[0:0] s9461, in9461_1, in9461_2;
    wire c9461;
    assign in9461_1 = {s6778[0]};
    assign in9461_2 = {s6779[0]};
    Full_Adder FA_9461(s9461, c9461, in9461_1, in9461_2, s6777[0]);
    wire[0:0] s9462, in9462_1, in9462_2;
    wire c9462;
    assign in9462_1 = {s6781[0]};
    assign in9462_2 = {s6782[0]};
    Full_Adder FA_9462(s9462, c9462, in9462_1, in9462_2, s6780[0]);
    wire[0:0] s9463, in9463_1, in9463_2;
    wire c9463;
    assign in9463_1 = {s6784[0]};
    assign in9463_2 = {s6785[0]};
    Full_Adder FA_9463(s9463, c9463, in9463_1, in9463_2, s6783[0]);
    wire[0:0] s9464, in9464_1, in9464_2;
    wire c9464;
    assign in9464_1 = {s6787[0]};
    assign in9464_2 = {s6788[0]};
    Full_Adder FA_9464(s9464, c9464, in9464_1, in9464_2, s6786[0]);
    wire[0:0] s9465, in9465_1, in9465_2;
    wire c9465;
    assign in9465_1 = {s6790[0]};
    assign in9465_2 = {s6791[0]};
    Full_Adder FA_9465(s9465, c9465, in9465_1, in9465_2, s6789[0]);
    wire[0:0] s9466, in9466_1, in9466_2;
    wire c9466;
    assign in9466_1 = {s6793[0]};
    assign in9466_2 = {s6794[0]};
    Full_Adder FA_9466(s9466, c9466, in9466_1, in9466_2, s6792[0]);
    wire[0:0] s9467, in9467_1, in9467_2;
    wire c9467;
    assign in9467_1 = {c6776};
    assign in9467_2 = {c6777};
    Full_Adder FA_9467(s9467, c9467, in9467_1, in9467_2, s3864[0]);
    wire[0:0] s9468, in9468_1, in9468_2;
    wire c9468;
    assign in9468_1 = {c6779};
    assign in9468_2 = {c6780};
    Full_Adder FA_9468(s9468, c9468, in9468_1, in9468_2, c6778);
    wire[0:0] s9469, in9469_1, in9469_2;
    wire c9469;
    assign in9469_1 = {c6782};
    assign in9469_2 = {c6783};
    Full_Adder FA_9469(s9469, c9469, in9469_1, in9469_2, c6781);
    wire[0:0] s9470, in9470_1, in9470_2;
    wire c9470;
    assign in9470_1 = {c6785};
    assign in9470_2 = {c6786};
    Full_Adder FA_9470(s9470, c9470, in9470_1, in9470_2, c6784);
    wire[0:0] s9471, in9471_1, in9471_2;
    wire c9471;
    assign in9471_1 = {c6788};
    assign in9471_2 = {c6789};
    Full_Adder FA_9471(s9471, c9471, in9471_1, in9471_2, c6787);
    wire[0:0] s9472, in9472_1, in9472_2;
    wire c9472;
    assign in9472_1 = {c6791};
    assign in9472_2 = {c6792};
    Full_Adder FA_9472(s9472, c9472, in9472_1, in9472_2, c6790);
    wire[0:0] s9473, in9473_1, in9473_2;
    wire c9473;
    assign in9473_1 = {c6794};
    assign in9473_2 = {s6795[0]};
    Full_Adder FA_9473(s9473, c9473, in9473_1, in9473_2, c6793);
    wire[0:0] s9474, in9474_1, in9474_2;
    wire c9474;
    assign in9474_1 = {s6797[0]};
    assign in9474_2 = {s6798[0]};
    Full_Adder FA_9474(s9474, c9474, in9474_1, in9474_2, s6796[0]);
    wire[0:0] s9475, in9475_1, in9475_2;
    wire c9475;
    assign in9475_1 = {s6800[0]};
    assign in9475_2 = {s6801[0]};
    Full_Adder FA_9475(s9475, c9475, in9475_1, in9475_2, s6799[0]);
    wire[0:0] s9476, in9476_1, in9476_2;
    wire c9476;
    assign in9476_1 = {s6803[0]};
    assign in9476_2 = {s6804[0]};
    Full_Adder FA_9476(s9476, c9476, in9476_1, in9476_2, s6802[0]);
    wire[0:0] s9477, in9477_1, in9477_2;
    wire c9477;
    assign in9477_1 = {s6806[0]};
    assign in9477_2 = {s6807[0]};
    Full_Adder FA_9477(s9477, c9477, in9477_1, in9477_2, s6805[0]);
    wire[0:0] s9478, in9478_1, in9478_2;
    wire c9478;
    assign in9478_1 = {s6809[0]};
    assign in9478_2 = {s6810[0]};
    Full_Adder FA_9478(s9478, c9478, in9478_1, in9478_2, s6808[0]);
    wire[0:0] s9479, in9479_1, in9479_2;
    wire c9479;
    assign in9479_1 = {s6812[0]};
    assign in9479_2 = {s6813[0]};
    Full_Adder FA_9479(s9479, c9479, in9479_1, in9479_2, s6811[0]);
    wire[0:0] s9480, in9480_1, in9480_2;
    wire c9480;
    assign in9480_1 = {c6795};
    assign in9480_2 = {c6796};
    Full_Adder FA_9480(s9480, c9480, in9480_1, in9480_2, s3892[0]);
    wire[0:0] s9481, in9481_1, in9481_2;
    wire c9481;
    assign in9481_1 = {c6798};
    assign in9481_2 = {c6799};
    Full_Adder FA_9481(s9481, c9481, in9481_1, in9481_2, c6797);
    wire[0:0] s9482, in9482_1, in9482_2;
    wire c9482;
    assign in9482_1 = {c6801};
    assign in9482_2 = {c6802};
    Full_Adder FA_9482(s9482, c9482, in9482_1, in9482_2, c6800);
    wire[0:0] s9483, in9483_1, in9483_2;
    wire c9483;
    assign in9483_1 = {c6804};
    assign in9483_2 = {c6805};
    Full_Adder FA_9483(s9483, c9483, in9483_1, in9483_2, c6803);
    wire[0:0] s9484, in9484_1, in9484_2;
    wire c9484;
    assign in9484_1 = {c6807};
    assign in9484_2 = {c6808};
    Full_Adder FA_9484(s9484, c9484, in9484_1, in9484_2, c6806);
    wire[0:0] s9485, in9485_1, in9485_2;
    wire c9485;
    assign in9485_1 = {c6810};
    assign in9485_2 = {c6811};
    Full_Adder FA_9485(s9485, c9485, in9485_1, in9485_2, c6809);
    wire[0:0] s9486, in9486_1, in9486_2;
    wire c9486;
    assign in9486_1 = {c6813};
    assign in9486_2 = {s6814[0]};
    Full_Adder FA_9486(s9486, c9486, in9486_1, in9486_2, c6812);
    wire[0:0] s9487, in9487_1, in9487_2;
    wire c9487;
    assign in9487_1 = {s6816[0]};
    assign in9487_2 = {s6817[0]};
    Full_Adder FA_9487(s9487, c9487, in9487_1, in9487_2, s6815[0]);
    wire[0:0] s9488, in9488_1, in9488_2;
    wire c9488;
    assign in9488_1 = {s6819[0]};
    assign in9488_2 = {s6820[0]};
    Full_Adder FA_9488(s9488, c9488, in9488_1, in9488_2, s6818[0]);
    wire[0:0] s9489, in9489_1, in9489_2;
    wire c9489;
    assign in9489_1 = {s6822[0]};
    assign in9489_2 = {s6823[0]};
    Full_Adder FA_9489(s9489, c9489, in9489_1, in9489_2, s6821[0]);
    wire[0:0] s9490, in9490_1, in9490_2;
    wire c9490;
    assign in9490_1 = {s6825[0]};
    assign in9490_2 = {s6826[0]};
    Full_Adder FA_9490(s9490, c9490, in9490_1, in9490_2, s6824[0]);
    wire[0:0] s9491, in9491_1, in9491_2;
    wire c9491;
    assign in9491_1 = {s6828[0]};
    assign in9491_2 = {s6829[0]};
    Full_Adder FA_9491(s9491, c9491, in9491_1, in9491_2, s6827[0]);
    wire[0:0] s9492, in9492_1, in9492_2;
    wire c9492;
    assign in9492_1 = {s6831[0]};
    assign in9492_2 = {s6832[0]};
    Full_Adder FA_9492(s9492, c9492, in9492_1, in9492_2, s6830[0]);
    wire[0:0] s9493, in9493_1, in9493_2;
    wire c9493;
    assign in9493_1 = {c6814};
    assign in9493_2 = {c6815};
    Full_Adder FA_9493(s9493, c9493, in9493_1, in9493_2, s3920[0]);
    wire[0:0] s9494, in9494_1, in9494_2;
    wire c9494;
    assign in9494_1 = {c6817};
    assign in9494_2 = {c6818};
    Full_Adder FA_9494(s9494, c9494, in9494_1, in9494_2, c6816);
    wire[0:0] s9495, in9495_1, in9495_2;
    wire c9495;
    assign in9495_1 = {c6820};
    assign in9495_2 = {c6821};
    Full_Adder FA_9495(s9495, c9495, in9495_1, in9495_2, c6819);
    wire[0:0] s9496, in9496_1, in9496_2;
    wire c9496;
    assign in9496_1 = {c6823};
    assign in9496_2 = {c6824};
    Full_Adder FA_9496(s9496, c9496, in9496_1, in9496_2, c6822);
    wire[0:0] s9497, in9497_1, in9497_2;
    wire c9497;
    assign in9497_1 = {c6826};
    assign in9497_2 = {c6827};
    Full_Adder FA_9497(s9497, c9497, in9497_1, in9497_2, c6825);
    wire[0:0] s9498, in9498_1, in9498_2;
    wire c9498;
    assign in9498_1 = {c6829};
    assign in9498_2 = {c6830};
    Full_Adder FA_9498(s9498, c9498, in9498_1, in9498_2, c6828);
    wire[0:0] s9499, in9499_1, in9499_2;
    wire c9499;
    assign in9499_1 = {c6832};
    assign in9499_2 = {s6833[0]};
    Full_Adder FA_9499(s9499, c9499, in9499_1, in9499_2, c6831);
    wire[0:0] s9500, in9500_1, in9500_2;
    wire c9500;
    assign in9500_1 = {s6835[0]};
    assign in9500_2 = {s6836[0]};
    Full_Adder FA_9500(s9500, c9500, in9500_1, in9500_2, s6834[0]);
    wire[0:0] s9501, in9501_1, in9501_2;
    wire c9501;
    assign in9501_1 = {s6838[0]};
    assign in9501_2 = {s6839[0]};
    Full_Adder FA_9501(s9501, c9501, in9501_1, in9501_2, s6837[0]);
    wire[0:0] s9502, in9502_1, in9502_2;
    wire c9502;
    assign in9502_1 = {s6841[0]};
    assign in9502_2 = {s6842[0]};
    Full_Adder FA_9502(s9502, c9502, in9502_1, in9502_2, s6840[0]);
    wire[0:0] s9503, in9503_1, in9503_2;
    wire c9503;
    assign in9503_1 = {s6844[0]};
    assign in9503_2 = {s6845[0]};
    Full_Adder FA_9503(s9503, c9503, in9503_1, in9503_2, s6843[0]);
    wire[0:0] s9504, in9504_1, in9504_2;
    wire c9504;
    assign in9504_1 = {s6847[0]};
    assign in9504_2 = {s6848[0]};
    Full_Adder FA_9504(s9504, c9504, in9504_1, in9504_2, s6846[0]);
    wire[0:0] s9505, in9505_1, in9505_2;
    wire c9505;
    assign in9505_1 = {s6850[0]};
    assign in9505_2 = {s6851[0]};
    Full_Adder FA_9505(s9505, c9505, in9505_1, in9505_2, s6849[0]);
    wire[0:0] s9506, in9506_1, in9506_2;
    wire c9506;
    assign in9506_1 = {c6833};
    assign in9506_2 = {c6834};
    Full_Adder FA_9506(s9506, c9506, in9506_1, in9506_2, s3948[0]);
    wire[0:0] s9507, in9507_1, in9507_2;
    wire c9507;
    assign in9507_1 = {c6836};
    assign in9507_2 = {c6837};
    Full_Adder FA_9507(s9507, c9507, in9507_1, in9507_2, c6835);
    wire[0:0] s9508, in9508_1, in9508_2;
    wire c9508;
    assign in9508_1 = {c6839};
    assign in9508_2 = {c6840};
    Full_Adder FA_9508(s9508, c9508, in9508_1, in9508_2, c6838);
    wire[0:0] s9509, in9509_1, in9509_2;
    wire c9509;
    assign in9509_1 = {c6842};
    assign in9509_2 = {c6843};
    Full_Adder FA_9509(s9509, c9509, in9509_1, in9509_2, c6841);
    wire[0:0] s9510, in9510_1, in9510_2;
    wire c9510;
    assign in9510_1 = {c6845};
    assign in9510_2 = {c6846};
    Full_Adder FA_9510(s9510, c9510, in9510_1, in9510_2, c6844);
    wire[0:0] s9511, in9511_1, in9511_2;
    wire c9511;
    assign in9511_1 = {c6848};
    assign in9511_2 = {c6849};
    Full_Adder FA_9511(s9511, c9511, in9511_1, in9511_2, c6847);
    wire[0:0] s9512, in9512_1, in9512_2;
    wire c9512;
    assign in9512_1 = {c6851};
    assign in9512_2 = {s6852[0]};
    Full_Adder FA_9512(s9512, c9512, in9512_1, in9512_2, c6850);
    wire[0:0] s9513, in9513_1, in9513_2;
    wire c9513;
    assign in9513_1 = {s6854[0]};
    assign in9513_2 = {s6855[0]};
    Full_Adder FA_9513(s9513, c9513, in9513_1, in9513_2, s6853[0]);
    wire[0:0] s9514, in9514_1, in9514_2;
    wire c9514;
    assign in9514_1 = {s6857[0]};
    assign in9514_2 = {s6858[0]};
    Full_Adder FA_9514(s9514, c9514, in9514_1, in9514_2, s6856[0]);
    wire[0:0] s9515, in9515_1, in9515_2;
    wire c9515;
    assign in9515_1 = {s6860[0]};
    assign in9515_2 = {s6861[0]};
    Full_Adder FA_9515(s9515, c9515, in9515_1, in9515_2, s6859[0]);
    wire[0:0] s9516, in9516_1, in9516_2;
    wire c9516;
    assign in9516_1 = {s6863[0]};
    assign in9516_2 = {s6864[0]};
    Full_Adder FA_9516(s9516, c9516, in9516_1, in9516_2, s6862[0]);
    wire[0:0] s9517, in9517_1, in9517_2;
    wire c9517;
    assign in9517_1 = {s6866[0]};
    assign in9517_2 = {s6867[0]};
    Full_Adder FA_9517(s9517, c9517, in9517_1, in9517_2, s6865[0]);
    wire[0:0] s9518, in9518_1, in9518_2;
    wire c9518;
    assign in9518_1 = {s6869[0]};
    assign in9518_2 = {s6870[0]};
    Full_Adder FA_9518(s9518, c9518, in9518_1, in9518_2, s6868[0]);
    wire[0:0] s9519, in9519_1, in9519_2;
    wire c9519;
    assign in9519_1 = {c6852};
    assign in9519_2 = {c6853};
    Full_Adder FA_9519(s9519, c9519, in9519_1, in9519_2, s3976[0]);
    wire[0:0] s9520, in9520_1, in9520_2;
    wire c9520;
    assign in9520_1 = {c6855};
    assign in9520_2 = {c6856};
    Full_Adder FA_9520(s9520, c9520, in9520_1, in9520_2, c6854);
    wire[0:0] s9521, in9521_1, in9521_2;
    wire c9521;
    assign in9521_1 = {c6858};
    assign in9521_2 = {c6859};
    Full_Adder FA_9521(s9521, c9521, in9521_1, in9521_2, c6857);
    wire[0:0] s9522, in9522_1, in9522_2;
    wire c9522;
    assign in9522_1 = {c6861};
    assign in9522_2 = {c6862};
    Full_Adder FA_9522(s9522, c9522, in9522_1, in9522_2, c6860);
    wire[0:0] s9523, in9523_1, in9523_2;
    wire c9523;
    assign in9523_1 = {c6864};
    assign in9523_2 = {c6865};
    Full_Adder FA_9523(s9523, c9523, in9523_1, in9523_2, c6863);
    wire[0:0] s9524, in9524_1, in9524_2;
    wire c9524;
    assign in9524_1 = {c6867};
    assign in9524_2 = {c6868};
    Full_Adder FA_9524(s9524, c9524, in9524_1, in9524_2, c6866);
    wire[0:0] s9525, in9525_1, in9525_2;
    wire c9525;
    assign in9525_1 = {c6870};
    assign in9525_2 = {s6871[0]};
    Full_Adder FA_9525(s9525, c9525, in9525_1, in9525_2, c6869);
    wire[0:0] s9526, in9526_1, in9526_2;
    wire c9526;
    assign in9526_1 = {s6873[0]};
    assign in9526_2 = {s6874[0]};
    Full_Adder FA_9526(s9526, c9526, in9526_1, in9526_2, s6872[0]);
    wire[0:0] s9527, in9527_1, in9527_2;
    wire c9527;
    assign in9527_1 = {s6876[0]};
    assign in9527_2 = {s6877[0]};
    Full_Adder FA_9527(s9527, c9527, in9527_1, in9527_2, s6875[0]);
    wire[0:0] s9528, in9528_1, in9528_2;
    wire c9528;
    assign in9528_1 = {s6879[0]};
    assign in9528_2 = {s6880[0]};
    Full_Adder FA_9528(s9528, c9528, in9528_1, in9528_2, s6878[0]);
    wire[0:0] s9529, in9529_1, in9529_2;
    wire c9529;
    assign in9529_1 = {s6882[0]};
    assign in9529_2 = {s6883[0]};
    Full_Adder FA_9529(s9529, c9529, in9529_1, in9529_2, s6881[0]);
    wire[0:0] s9530, in9530_1, in9530_2;
    wire c9530;
    assign in9530_1 = {s6885[0]};
    assign in9530_2 = {s6886[0]};
    Full_Adder FA_9530(s9530, c9530, in9530_1, in9530_2, s6884[0]);
    wire[0:0] s9531, in9531_1, in9531_2;
    wire c9531;
    assign in9531_1 = {s6888[0]};
    assign in9531_2 = {s6889[0]};
    Full_Adder FA_9531(s9531, c9531, in9531_1, in9531_2, s6887[0]);
    wire[0:0] s9532, in9532_1, in9532_2;
    wire c9532;
    assign in9532_1 = {c6871};
    assign in9532_2 = {c6872};
    Full_Adder FA_9532(s9532, c9532, in9532_1, in9532_2, s4004[0]);
    wire[0:0] s9533, in9533_1, in9533_2;
    wire c9533;
    assign in9533_1 = {c6874};
    assign in9533_2 = {c6875};
    Full_Adder FA_9533(s9533, c9533, in9533_1, in9533_2, c6873);
    wire[0:0] s9534, in9534_1, in9534_2;
    wire c9534;
    assign in9534_1 = {c6877};
    assign in9534_2 = {c6878};
    Full_Adder FA_9534(s9534, c9534, in9534_1, in9534_2, c6876);
    wire[0:0] s9535, in9535_1, in9535_2;
    wire c9535;
    assign in9535_1 = {c6880};
    assign in9535_2 = {c6881};
    Full_Adder FA_9535(s9535, c9535, in9535_1, in9535_2, c6879);
    wire[0:0] s9536, in9536_1, in9536_2;
    wire c9536;
    assign in9536_1 = {c6883};
    assign in9536_2 = {c6884};
    Full_Adder FA_9536(s9536, c9536, in9536_1, in9536_2, c6882);
    wire[0:0] s9537, in9537_1, in9537_2;
    wire c9537;
    assign in9537_1 = {c6886};
    assign in9537_2 = {c6887};
    Full_Adder FA_9537(s9537, c9537, in9537_1, in9537_2, c6885);
    wire[0:0] s9538, in9538_1, in9538_2;
    wire c9538;
    assign in9538_1 = {c6889};
    assign in9538_2 = {s6890[0]};
    Full_Adder FA_9538(s9538, c9538, in9538_1, in9538_2, c6888);
    wire[0:0] s9539, in9539_1, in9539_2;
    wire c9539;
    assign in9539_1 = {s6892[0]};
    assign in9539_2 = {s6893[0]};
    Full_Adder FA_9539(s9539, c9539, in9539_1, in9539_2, s6891[0]);
    wire[0:0] s9540, in9540_1, in9540_2;
    wire c9540;
    assign in9540_1 = {s6895[0]};
    assign in9540_2 = {s6896[0]};
    Full_Adder FA_9540(s9540, c9540, in9540_1, in9540_2, s6894[0]);
    wire[0:0] s9541, in9541_1, in9541_2;
    wire c9541;
    assign in9541_1 = {s6898[0]};
    assign in9541_2 = {s6899[0]};
    Full_Adder FA_9541(s9541, c9541, in9541_1, in9541_2, s6897[0]);
    wire[0:0] s9542, in9542_1, in9542_2;
    wire c9542;
    assign in9542_1 = {s6901[0]};
    assign in9542_2 = {s6902[0]};
    Full_Adder FA_9542(s9542, c9542, in9542_1, in9542_2, s6900[0]);
    wire[0:0] s9543, in9543_1, in9543_2;
    wire c9543;
    assign in9543_1 = {s6904[0]};
    assign in9543_2 = {s6905[0]};
    Full_Adder FA_9543(s9543, c9543, in9543_1, in9543_2, s6903[0]);
    wire[0:0] s9544, in9544_1, in9544_2;
    wire c9544;
    assign in9544_1 = {s6907[0]};
    assign in9544_2 = {s6908[0]};
    Full_Adder FA_9544(s9544, c9544, in9544_1, in9544_2, s6906[0]);
    wire[0:0] s9545, in9545_1, in9545_2;
    wire c9545;
    assign in9545_1 = {c6890};
    assign in9545_2 = {c6891};
    Full_Adder FA_9545(s9545, c9545, in9545_1, in9545_2, s4032[0]);
    wire[0:0] s9546, in9546_1, in9546_2;
    wire c9546;
    assign in9546_1 = {c6893};
    assign in9546_2 = {c6894};
    Full_Adder FA_9546(s9546, c9546, in9546_1, in9546_2, c6892);
    wire[0:0] s9547, in9547_1, in9547_2;
    wire c9547;
    assign in9547_1 = {c6896};
    assign in9547_2 = {c6897};
    Full_Adder FA_9547(s9547, c9547, in9547_1, in9547_2, c6895);
    wire[0:0] s9548, in9548_1, in9548_2;
    wire c9548;
    assign in9548_1 = {c6899};
    assign in9548_2 = {c6900};
    Full_Adder FA_9548(s9548, c9548, in9548_1, in9548_2, c6898);
    wire[0:0] s9549, in9549_1, in9549_2;
    wire c9549;
    assign in9549_1 = {c6902};
    assign in9549_2 = {c6903};
    Full_Adder FA_9549(s9549, c9549, in9549_1, in9549_2, c6901);
    wire[0:0] s9550, in9550_1, in9550_2;
    wire c9550;
    assign in9550_1 = {c6905};
    assign in9550_2 = {c6906};
    Full_Adder FA_9550(s9550, c9550, in9550_1, in9550_2, c6904);
    wire[0:0] s9551, in9551_1, in9551_2;
    wire c9551;
    assign in9551_1 = {c6908};
    assign in9551_2 = {s6909[0]};
    Full_Adder FA_9551(s9551, c9551, in9551_1, in9551_2, c6907);
    wire[0:0] s9552, in9552_1, in9552_2;
    wire c9552;
    assign in9552_1 = {s6911[0]};
    assign in9552_2 = {s6912[0]};
    Full_Adder FA_9552(s9552, c9552, in9552_1, in9552_2, s6910[0]);
    wire[0:0] s9553, in9553_1, in9553_2;
    wire c9553;
    assign in9553_1 = {s6914[0]};
    assign in9553_2 = {s6915[0]};
    Full_Adder FA_9553(s9553, c9553, in9553_1, in9553_2, s6913[0]);
    wire[0:0] s9554, in9554_1, in9554_2;
    wire c9554;
    assign in9554_1 = {s6917[0]};
    assign in9554_2 = {s6918[0]};
    Full_Adder FA_9554(s9554, c9554, in9554_1, in9554_2, s6916[0]);
    wire[0:0] s9555, in9555_1, in9555_2;
    wire c9555;
    assign in9555_1 = {s6920[0]};
    assign in9555_2 = {s6921[0]};
    Full_Adder FA_9555(s9555, c9555, in9555_1, in9555_2, s6919[0]);
    wire[0:0] s9556, in9556_1, in9556_2;
    wire c9556;
    assign in9556_1 = {s6923[0]};
    assign in9556_2 = {s6924[0]};
    Full_Adder FA_9556(s9556, c9556, in9556_1, in9556_2, s6922[0]);
    wire[0:0] s9557, in9557_1, in9557_2;
    wire c9557;
    assign in9557_1 = {s6926[0]};
    assign in9557_2 = {s6927[0]};
    Full_Adder FA_9557(s9557, c9557, in9557_1, in9557_2, s6925[0]);
    wire[0:0] s9558, in9558_1, in9558_2;
    wire c9558;
    assign in9558_1 = {c6909};
    assign in9558_2 = {c6910};
    Full_Adder FA_9558(s9558, c9558, in9558_1, in9558_2, s4060[0]);
    wire[0:0] s9559, in9559_1, in9559_2;
    wire c9559;
    assign in9559_1 = {c6912};
    assign in9559_2 = {c6913};
    Full_Adder FA_9559(s9559, c9559, in9559_1, in9559_2, c6911);
    wire[0:0] s9560, in9560_1, in9560_2;
    wire c9560;
    assign in9560_1 = {c6915};
    assign in9560_2 = {c6916};
    Full_Adder FA_9560(s9560, c9560, in9560_1, in9560_2, c6914);
    wire[0:0] s9561, in9561_1, in9561_2;
    wire c9561;
    assign in9561_1 = {c6918};
    assign in9561_2 = {c6919};
    Full_Adder FA_9561(s9561, c9561, in9561_1, in9561_2, c6917);
    wire[0:0] s9562, in9562_1, in9562_2;
    wire c9562;
    assign in9562_1 = {c6921};
    assign in9562_2 = {c6922};
    Full_Adder FA_9562(s9562, c9562, in9562_1, in9562_2, c6920);
    wire[0:0] s9563, in9563_1, in9563_2;
    wire c9563;
    assign in9563_1 = {c6924};
    assign in9563_2 = {c6925};
    Full_Adder FA_9563(s9563, c9563, in9563_1, in9563_2, c6923);
    wire[0:0] s9564, in9564_1, in9564_2;
    wire c9564;
    assign in9564_1 = {c6927};
    assign in9564_2 = {s6928[0]};
    Full_Adder FA_9564(s9564, c9564, in9564_1, in9564_2, c6926);
    wire[0:0] s9565, in9565_1, in9565_2;
    wire c9565;
    assign in9565_1 = {s6930[0]};
    assign in9565_2 = {s6931[0]};
    Full_Adder FA_9565(s9565, c9565, in9565_1, in9565_2, s6929[0]);
    wire[0:0] s9566, in9566_1, in9566_2;
    wire c9566;
    assign in9566_1 = {s6933[0]};
    assign in9566_2 = {s6934[0]};
    Full_Adder FA_9566(s9566, c9566, in9566_1, in9566_2, s6932[0]);
    wire[0:0] s9567, in9567_1, in9567_2;
    wire c9567;
    assign in9567_1 = {s6936[0]};
    assign in9567_2 = {s6937[0]};
    Full_Adder FA_9567(s9567, c9567, in9567_1, in9567_2, s6935[0]);
    wire[0:0] s9568, in9568_1, in9568_2;
    wire c9568;
    assign in9568_1 = {s6939[0]};
    assign in9568_2 = {s6940[0]};
    Full_Adder FA_9568(s9568, c9568, in9568_1, in9568_2, s6938[0]);
    wire[0:0] s9569, in9569_1, in9569_2;
    wire c9569;
    assign in9569_1 = {s6942[0]};
    assign in9569_2 = {s6943[0]};
    Full_Adder FA_9569(s9569, c9569, in9569_1, in9569_2, s6941[0]);
    wire[0:0] s9570, in9570_1, in9570_2;
    wire c9570;
    assign in9570_1 = {s6945[0]};
    assign in9570_2 = {s6946[0]};
    Full_Adder FA_9570(s9570, c9570, in9570_1, in9570_2, s6944[0]);
    wire[0:0] s9571, in9571_1, in9571_2;
    wire c9571;
    assign in9571_1 = {c6928};
    assign in9571_2 = {c6929};
    Full_Adder FA_9571(s9571, c9571, in9571_1, in9571_2, s4088[0]);
    wire[0:0] s9572, in9572_1, in9572_2;
    wire c9572;
    assign in9572_1 = {c6931};
    assign in9572_2 = {c6932};
    Full_Adder FA_9572(s9572, c9572, in9572_1, in9572_2, c6930);
    wire[0:0] s9573, in9573_1, in9573_2;
    wire c9573;
    assign in9573_1 = {c6934};
    assign in9573_2 = {c6935};
    Full_Adder FA_9573(s9573, c9573, in9573_1, in9573_2, c6933);
    wire[0:0] s9574, in9574_1, in9574_2;
    wire c9574;
    assign in9574_1 = {c6937};
    assign in9574_2 = {c6938};
    Full_Adder FA_9574(s9574, c9574, in9574_1, in9574_2, c6936);
    wire[0:0] s9575, in9575_1, in9575_2;
    wire c9575;
    assign in9575_1 = {c6940};
    assign in9575_2 = {c6941};
    Full_Adder FA_9575(s9575, c9575, in9575_1, in9575_2, c6939);
    wire[0:0] s9576, in9576_1, in9576_2;
    wire c9576;
    assign in9576_1 = {c6943};
    assign in9576_2 = {c6944};
    Full_Adder FA_9576(s9576, c9576, in9576_1, in9576_2, c6942);
    wire[0:0] s9577, in9577_1, in9577_2;
    wire c9577;
    assign in9577_1 = {c6946};
    assign in9577_2 = {s6947[0]};
    Full_Adder FA_9577(s9577, c9577, in9577_1, in9577_2, c6945);
    wire[0:0] s9578, in9578_1, in9578_2;
    wire c9578;
    assign in9578_1 = {s6949[0]};
    assign in9578_2 = {s6950[0]};
    Full_Adder FA_9578(s9578, c9578, in9578_1, in9578_2, s6948[0]);
    wire[0:0] s9579, in9579_1, in9579_2;
    wire c9579;
    assign in9579_1 = {s6952[0]};
    assign in9579_2 = {s6953[0]};
    Full_Adder FA_9579(s9579, c9579, in9579_1, in9579_2, s6951[0]);
    wire[0:0] s9580, in9580_1, in9580_2;
    wire c9580;
    assign in9580_1 = {s6955[0]};
    assign in9580_2 = {s6956[0]};
    Full_Adder FA_9580(s9580, c9580, in9580_1, in9580_2, s6954[0]);
    wire[0:0] s9581, in9581_1, in9581_2;
    wire c9581;
    assign in9581_1 = {s6958[0]};
    assign in9581_2 = {s6959[0]};
    Full_Adder FA_9581(s9581, c9581, in9581_1, in9581_2, s6957[0]);
    wire[0:0] s9582, in9582_1, in9582_2;
    wire c9582;
    assign in9582_1 = {s6961[0]};
    assign in9582_2 = {s6962[0]};
    Full_Adder FA_9582(s9582, c9582, in9582_1, in9582_2, s6960[0]);
    wire[0:0] s9583, in9583_1, in9583_2;
    wire c9583;
    assign in9583_1 = {s6964[0]};
    assign in9583_2 = {s6965[0]};
    Full_Adder FA_9583(s9583, c9583, in9583_1, in9583_2, s6963[0]);
    wire[0:0] s9584, in9584_1, in9584_2;
    wire c9584;
    assign in9584_1 = {c6947};
    assign in9584_2 = {c6948};
    Full_Adder FA_9584(s9584, c9584, in9584_1, in9584_2, s4116[0]);
    wire[0:0] s9585, in9585_1, in9585_2;
    wire c9585;
    assign in9585_1 = {c6950};
    assign in9585_2 = {c6951};
    Full_Adder FA_9585(s9585, c9585, in9585_1, in9585_2, c6949);
    wire[0:0] s9586, in9586_1, in9586_2;
    wire c9586;
    assign in9586_1 = {c6953};
    assign in9586_2 = {c6954};
    Full_Adder FA_9586(s9586, c9586, in9586_1, in9586_2, c6952);
    wire[0:0] s9587, in9587_1, in9587_2;
    wire c9587;
    assign in9587_1 = {c6956};
    assign in9587_2 = {c6957};
    Full_Adder FA_9587(s9587, c9587, in9587_1, in9587_2, c6955);
    wire[0:0] s9588, in9588_1, in9588_2;
    wire c9588;
    assign in9588_1 = {c6959};
    assign in9588_2 = {c6960};
    Full_Adder FA_9588(s9588, c9588, in9588_1, in9588_2, c6958);
    wire[0:0] s9589, in9589_1, in9589_2;
    wire c9589;
    assign in9589_1 = {c6962};
    assign in9589_2 = {c6963};
    Full_Adder FA_9589(s9589, c9589, in9589_1, in9589_2, c6961);
    wire[0:0] s9590, in9590_1, in9590_2;
    wire c9590;
    assign in9590_1 = {c6965};
    assign in9590_2 = {s6966[0]};
    Full_Adder FA_9590(s9590, c9590, in9590_1, in9590_2, c6964);
    wire[0:0] s9591, in9591_1, in9591_2;
    wire c9591;
    assign in9591_1 = {s6968[0]};
    assign in9591_2 = {s6969[0]};
    Full_Adder FA_9591(s9591, c9591, in9591_1, in9591_2, s6967[0]);
    wire[0:0] s9592, in9592_1, in9592_2;
    wire c9592;
    assign in9592_1 = {s6971[0]};
    assign in9592_2 = {s6972[0]};
    Full_Adder FA_9592(s9592, c9592, in9592_1, in9592_2, s6970[0]);
    wire[0:0] s9593, in9593_1, in9593_2;
    wire c9593;
    assign in9593_1 = {s6974[0]};
    assign in9593_2 = {s6975[0]};
    Full_Adder FA_9593(s9593, c9593, in9593_1, in9593_2, s6973[0]);
    wire[0:0] s9594, in9594_1, in9594_2;
    wire c9594;
    assign in9594_1 = {s6977[0]};
    assign in9594_2 = {s6978[0]};
    Full_Adder FA_9594(s9594, c9594, in9594_1, in9594_2, s6976[0]);
    wire[0:0] s9595, in9595_1, in9595_2;
    wire c9595;
    assign in9595_1 = {s6980[0]};
    assign in9595_2 = {s6981[0]};
    Full_Adder FA_9595(s9595, c9595, in9595_1, in9595_2, s6979[0]);
    wire[0:0] s9596, in9596_1, in9596_2;
    wire c9596;
    assign in9596_1 = {s6983[0]};
    assign in9596_2 = {s6984[0]};
    Full_Adder FA_9596(s9596, c9596, in9596_1, in9596_2, s6982[0]);
    wire[0:0] s9597, in9597_1, in9597_2;
    wire c9597;
    assign in9597_1 = {c6966};
    assign in9597_2 = {c6967};
    Full_Adder FA_9597(s9597, c9597, in9597_1, in9597_2, s4144[0]);
    wire[0:0] s9598, in9598_1, in9598_2;
    wire c9598;
    assign in9598_1 = {c6969};
    assign in9598_2 = {c6970};
    Full_Adder FA_9598(s9598, c9598, in9598_1, in9598_2, c6968);
    wire[0:0] s9599, in9599_1, in9599_2;
    wire c9599;
    assign in9599_1 = {c6972};
    assign in9599_2 = {c6973};
    Full_Adder FA_9599(s9599, c9599, in9599_1, in9599_2, c6971);
    wire[0:0] s9600, in9600_1, in9600_2;
    wire c9600;
    assign in9600_1 = {c6975};
    assign in9600_2 = {c6976};
    Full_Adder FA_9600(s9600, c9600, in9600_1, in9600_2, c6974);
    wire[0:0] s9601, in9601_1, in9601_2;
    wire c9601;
    assign in9601_1 = {c6978};
    assign in9601_2 = {c6979};
    Full_Adder FA_9601(s9601, c9601, in9601_1, in9601_2, c6977);
    wire[0:0] s9602, in9602_1, in9602_2;
    wire c9602;
    assign in9602_1 = {c6981};
    assign in9602_2 = {c6982};
    Full_Adder FA_9602(s9602, c9602, in9602_1, in9602_2, c6980);
    wire[0:0] s9603, in9603_1, in9603_2;
    wire c9603;
    assign in9603_1 = {c6984};
    assign in9603_2 = {s6985[0]};
    Full_Adder FA_9603(s9603, c9603, in9603_1, in9603_2, c6983);
    wire[0:0] s9604, in9604_1, in9604_2;
    wire c9604;
    assign in9604_1 = {s6987[0]};
    assign in9604_2 = {s6988[0]};
    Full_Adder FA_9604(s9604, c9604, in9604_1, in9604_2, s6986[0]);
    wire[0:0] s9605, in9605_1, in9605_2;
    wire c9605;
    assign in9605_1 = {s6990[0]};
    assign in9605_2 = {s6991[0]};
    Full_Adder FA_9605(s9605, c9605, in9605_1, in9605_2, s6989[0]);
    wire[0:0] s9606, in9606_1, in9606_2;
    wire c9606;
    assign in9606_1 = {s6993[0]};
    assign in9606_2 = {s6994[0]};
    Full_Adder FA_9606(s9606, c9606, in9606_1, in9606_2, s6992[0]);
    wire[0:0] s9607, in9607_1, in9607_2;
    wire c9607;
    assign in9607_1 = {s6996[0]};
    assign in9607_2 = {s6997[0]};
    Full_Adder FA_9607(s9607, c9607, in9607_1, in9607_2, s6995[0]);
    wire[0:0] s9608, in9608_1, in9608_2;
    wire c9608;
    assign in9608_1 = {s6999[0]};
    assign in9608_2 = {s7000[0]};
    Full_Adder FA_9608(s9608, c9608, in9608_1, in9608_2, s6998[0]);
    wire[0:0] s9609, in9609_1, in9609_2;
    wire c9609;
    assign in9609_1 = {s7002[0]};
    assign in9609_2 = {s7003[0]};
    Full_Adder FA_9609(s9609, c9609, in9609_1, in9609_2, s7001[0]);
    wire[0:0] s9610, in9610_1, in9610_2;
    wire c9610;
    assign in9610_1 = {c6985};
    assign in9610_2 = {c6986};
    Full_Adder FA_9610(s9610, c9610, in9610_1, in9610_2, s4172[0]);
    wire[0:0] s9611, in9611_1, in9611_2;
    wire c9611;
    assign in9611_1 = {c6988};
    assign in9611_2 = {c6989};
    Full_Adder FA_9611(s9611, c9611, in9611_1, in9611_2, c6987);
    wire[0:0] s9612, in9612_1, in9612_2;
    wire c9612;
    assign in9612_1 = {c6991};
    assign in9612_2 = {c6992};
    Full_Adder FA_9612(s9612, c9612, in9612_1, in9612_2, c6990);
    wire[0:0] s9613, in9613_1, in9613_2;
    wire c9613;
    assign in9613_1 = {c6994};
    assign in9613_2 = {c6995};
    Full_Adder FA_9613(s9613, c9613, in9613_1, in9613_2, c6993);
    wire[0:0] s9614, in9614_1, in9614_2;
    wire c9614;
    assign in9614_1 = {c6997};
    assign in9614_2 = {c6998};
    Full_Adder FA_9614(s9614, c9614, in9614_1, in9614_2, c6996);
    wire[0:0] s9615, in9615_1, in9615_2;
    wire c9615;
    assign in9615_1 = {c7000};
    assign in9615_2 = {c7001};
    Full_Adder FA_9615(s9615, c9615, in9615_1, in9615_2, c6999);
    wire[0:0] s9616, in9616_1, in9616_2;
    wire c9616;
    assign in9616_1 = {c7003};
    assign in9616_2 = {s7004[0]};
    Full_Adder FA_9616(s9616, c9616, in9616_1, in9616_2, c7002);
    wire[0:0] s9617, in9617_1, in9617_2;
    wire c9617;
    assign in9617_1 = {s7006[0]};
    assign in9617_2 = {s7007[0]};
    Full_Adder FA_9617(s9617, c9617, in9617_1, in9617_2, s7005[0]);
    wire[0:0] s9618, in9618_1, in9618_2;
    wire c9618;
    assign in9618_1 = {s7009[0]};
    assign in9618_2 = {s7010[0]};
    Full_Adder FA_9618(s9618, c9618, in9618_1, in9618_2, s7008[0]);
    wire[0:0] s9619, in9619_1, in9619_2;
    wire c9619;
    assign in9619_1 = {s7012[0]};
    assign in9619_2 = {s7013[0]};
    Full_Adder FA_9619(s9619, c9619, in9619_1, in9619_2, s7011[0]);
    wire[0:0] s9620, in9620_1, in9620_2;
    wire c9620;
    assign in9620_1 = {s7015[0]};
    assign in9620_2 = {s7016[0]};
    Full_Adder FA_9620(s9620, c9620, in9620_1, in9620_2, s7014[0]);
    wire[0:0] s9621, in9621_1, in9621_2;
    wire c9621;
    assign in9621_1 = {s7018[0]};
    assign in9621_2 = {s7019[0]};
    Full_Adder FA_9621(s9621, c9621, in9621_1, in9621_2, s7017[0]);
    wire[0:0] s9622, in9622_1, in9622_2;
    wire c9622;
    assign in9622_1 = {s7021[0]};
    assign in9622_2 = {s7022[0]};
    Full_Adder FA_9622(s9622, c9622, in9622_1, in9622_2, s7020[0]);
    wire[0:0] s9623, in9623_1, in9623_2;
    wire c9623;
    assign in9623_1 = {c7004};
    assign in9623_2 = {c7005};
    Full_Adder FA_9623(s9623, c9623, in9623_1, in9623_2, s4200[0]);
    wire[0:0] s9624, in9624_1, in9624_2;
    wire c9624;
    assign in9624_1 = {c7007};
    assign in9624_2 = {c7008};
    Full_Adder FA_9624(s9624, c9624, in9624_1, in9624_2, c7006);
    wire[0:0] s9625, in9625_1, in9625_2;
    wire c9625;
    assign in9625_1 = {c7010};
    assign in9625_2 = {c7011};
    Full_Adder FA_9625(s9625, c9625, in9625_1, in9625_2, c7009);
    wire[0:0] s9626, in9626_1, in9626_2;
    wire c9626;
    assign in9626_1 = {c7013};
    assign in9626_2 = {c7014};
    Full_Adder FA_9626(s9626, c9626, in9626_1, in9626_2, c7012);
    wire[0:0] s9627, in9627_1, in9627_2;
    wire c9627;
    assign in9627_1 = {c7016};
    assign in9627_2 = {c7017};
    Full_Adder FA_9627(s9627, c9627, in9627_1, in9627_2, c7015);
    wire[0:0] s9628, in9628_1, in9628_2;
    wire c9628;
    assign in9628_1 = {c7019};
    assign in9628_2 = {c7020};
    Full_Adder FA_9628(s9628, c9628, in9628_1, in9628_2, c7018);
    wire[0:0] s9629, in9629_1, in9629_2;
    wire c9629;
    assign in9629_1 = {c7022};
    assign in9629_2 = {s7023[0]};
    Full_Adder FA_9629(s9629, c9629, in9629_1, in9629_2, c7021);
    wire[0:0] s9630, in9630_1, in9630_2;
    wire c9630;
    assign in9630_1 = {s7025[0]};
    assign in9630_2 = {s7026[0]};
    Full_Adder FA_9630(s9630, c9630, in9630_1, in9630_2, s7024[0]);
    wire[0:0] s9631, in9631_1, in9631_2;
    wire c9631;
    assign in9631_1 = {s7028[0]};
    assign in9631_2 = {s7029[0]};
    Full_Adder FA_9631(s9631, c9631, in9631_1, in9631_2, s7027[0]);
    wire[0:0] s9632, in9632_1, in9632_2;
    wire c9632;
    assign in9632_1 = {s7031[0]};
    assign in9632_2 = {s7032[0]};
    Full_Adder FA_9632(s9632, c9632, in9632_1, in9632_2, s7030[0]);
    wire[0:0] s9633, in9633_1, in9633_2;
    wire c9633;
    assign in9633_1 = {s7034[0]};
    assign in9633_2 = {s7035[0]};
    Full_Adder FA_9633(s9633, c9633, in9633_1, in9633_2, s7033[0]);
    wire[0:0] s9634, in9634_1, in9634_2;
    wire c9634;
    assign in9634_1 = {s7037[0]};
    assign in9634_2 = {s7038[0]};
    Full_Adder FA_9634(s9634, c9634, in9634_1, in9634_2, s7036[0]);
    wire[0:0] s9635, in9635_1, in9635_2;
    wire c9635;
    assign in9635_1 = {s7040[0]};
    assign in9635_2 = {s7041[0]};
    Full_Adder FA_9635(s9635, c9635, in9635_1, in9635_2, s7039[0]);
    wire[0:0] s9636, in9636_1, in9636_2;
    wire c9636;
    assign in9636_1 = {c7023};
    assign in9636_2 = {c7024};
    Full_Adder FA_9636(s9636, c9636, in9636_1, in9636_2, s4228[0]);
    wire[0:0] s9637, in9637_1, in9637_2;
    wire c9637;
    assign in9637_1 = {c7026};
    assign in9637_2 = {c7027};
    Full_Adder FA_9637(s9637, c9637, in9637_1, in9637_2, c7025);
    wire[0:0] s9638, in9638_1, in9638_2;
    wire c9638;
    assign in9638_1 = {c7029};
    assign in9638_2 = {c7030};
    Full_Adder FA_9638(s9638, c9638, in9638_1, in9638_2, c7028);
    wire[0:0] s9639, in9639_1, in9639_2;
    wire c9639;
    assign in9639_1 = {c7032};
    assign in9639_2 = {c7033};
    Full_Adder FA_9639(s9639, c9639, in9639_1, in9639_2, c7031);
    wire[0:0] s9640, in9640_1, in9640_2;
    wire c9640;
    assign in9640_1 = {c7035};
    assign in9640_2 = {c7036};
    Full_Adder FA_9640(s9640, c9640, in9640_1, in9640_2, c7034);
    wire[0:0] s9641, in9641_1, in9641_2;
    wire c9641;
    assign in9641_1 = {c7038};
    assign in9641_2 = {c7039};
    Full_Adder FA_9641(s9641, c9641, in9641_1, in9641_2, c7037);
    wire[0:0] s9642, in9642_1, in9642_2;
    wire c9642;
    assign in9642_1 = {c7041};
    assign in9642_2 = {s7042[0]};
    Full_Adder FA_9642(s9642, c9642, in9642_1, in9642_2, c7040);
    wire[0:0] s9643, in9643_1, in9643_2;
    wire c9643;
    assign in9643_1 = {s7044[0]};
    assign in9643_2 = {s7045[0]};
    Full_Adder FA_9643(s9643, c9643, in9643_1, in9643_2, s7043[0]);
    wire[0:0] s9644, in9644_1, in9644_2;
    wire c9644;
    assign in9644_1 = {s7047[0]};
    assign in9644_2 = {s7048[0]};
    Full_Adder FA_9644(s9644, c9644, in9644_1, in9644_2, s7046[0]);
    wire[0:0] s9645, in9645_1, in9645_2;
    wire c9645;
    assign in9645_1 = {s7050[0]};
    assign in9645_2 = {s7051[0]};
    Full_Adder FA_9645(s9645, c9645, in9645_1, in9645_2, s7049[0]);
    wire[0:0] s9646, in9646_1, in9646_2;
    wire c9646;
    assign in9646_1 = {s7053[0]};
    assign in9646_2 = {s7054[0]};
    Full_Adder FA_9646(s9646, c9646, in9646_1, in9646_2, s7052[0]);
    wire[0:0] s9647, in9647_1, in9647_2;
    wire c9647;
    assign in9647_1 = {s7056[0]};
    assign in9647_2 = {s7057[0]};
    Full_Adder FA_9647(s9647, c9647, in9647_1, in9647_2, s7055[0]);
    wire[0:0] s9648, in9648_1, in9648_2;
    wire c9648;
    assign in9648_1 = {s7059[0]};
    assign in9648_2 = {s7060[0]};
    Full_Adder FA_9648(s9648, c9648, in9648_1, in9648_2, s7058[0]);
    wire[0:0] s9649, in9649_1, in9649_2;
    wire c9649;
    assign in9649_1 = {c7042};
    assign in9649_2 = {c7043};
    Full_Adder FA_9649(s9649, c9649, in9649_1, in9649_2, s4256[0]);
    wire[0:0] s9650, in9650_1, in9650_2;
    wire c9650;
    assign in9650_1 = {c7045};
    assign in9650_2 = {c7046};
    Full_Adder FA_9650(s9650, c9650, in9650_1, in9650_2, c7044);
    wire[0:0] s9651, in9651_1, in9651_2;
    wire c9651;
    assign in9651_1 = {c7048};
    assign in9651_2 = {c7049};
    Full_Adder FA_9651(s9651, c9651, in9651_1, in9651_2, c7047);
    wire[0:0] s9652, in9652_1, in9652_2;
    wire c9652;
    assign in9652_1 = {c7051};
    assign in9652_2 = {c7052};
    Full_Adder FA_9652(s9652, c9652, in9652_1, in9652_2, c7050);
    wire[0:0] s9653, in9653_1, in9653_2;
    wire c9653;
    assign in9653_1 = {c7054};
    assign in9653_2 = {c7055};
    Full_Adder FA_9653(s9653, c9653, in9653_1, in9653_2, c7053);
    wire[0:0] s9654, in9654_1, in9654_2;
    wire c9654;
    assign in9654_1 = {c7057};
    assign in9654_2 = {c7058};
    Full_Adder FA_9654(s9654, c9654, in9654_1, in9654_2, c7056);
    wire[0:0] s9655, in9655_1, in9655_2;
    wire c9655;
    assign in9655_1 = {c7060};
    assign in9655_2 = {s7061[0]};
    Full_Adder FA_9655(s9655, c9655, in9655_1, in9655_2, c7059);
    wire[0:0] s9656, in9656_1, in9656_2;
    wire c9656;
    assign in9656_1 = {s7063[0]};
    assign in9656_2 = {s7064[0]};
    Full_Adder FA_9656(s9656, c9656, in9656_1, in9656_2, s7062[0]);
    wire[0:0] s9657, in9657_1, in9657_2;
    wire c9657;
    assign in9657_1 = {s7066[0]};
    assign in9657_2 = {s7067[0]};
    Full_Adder FA_9657(s9657, c9657, in9657_1, in9657_2, s7065[0]);
    wire[0:0] s9658, in9658_1, in9658_2;
    wire c9658;
    assign in9658_1 = {s7069[0]};
    assign in9658_2 = {s7070[0]};
    Full_Adder FA_9658(s9658, c9658, in9658_1, in9658_2, s7068[0]);
    wire[0:0] s9659, in9659_1, in9659_2;
    wire c9659;
    assign in9659_1 = {s7072[0]};
    assign in9659_2 = {s7073[0]};
    Full_Adder FA_9659(s9659, c9659, in9659_1, in9659_2, s7071[0]);
    wire[0:0] s9660, in9660_1, in9660_2;
    wire c9660;
    assign in9660_1 = {s7075[0]};
    assign in9660_2 = {s7076[0]};
    Full_Adder FA_9660(s9660, c9660, in9660_1, in9660_2, s7074[0]);
    wire[0:0] s9661, in9661_1, in9661_2;
    wire c9661;
    assign in9661_1 = {s7078[0]};
    assign in9661_2 = {s7079[0]};
    Full_Adder FA_9661(s9661, c9661, in9661_1, in9661_2, s7077[0]);
    wire[0:0] s9662, in9662_1, in9662_2;
    wire c9662;
    assign in9662_1 = {c7061};
    assign in9662_2 = {c7062};
    Full_Adder FA_9662(s9662, c9662, in9662_1, in9662_2, s4284[0]);
    wire[0:0] s9663, in9663_1, in9663_2;
    wire c9663;
    assign in9663_1 = {c7064};
    assign in9663_2 = {c7065};
    Full_Adder FA_9663(s9663, c9663, in9663_1, in9663_2, c7063);
    wire[0:0] s9664, in9664_1, in9664_2;
    wire c9664;
    assign in9664_1 = {c7067};
    assign in9664_2 = {c7068};
    Full_Adder FA_9664(s9664, c9664, in9664_1, in9664_2, c7066);
    wire[0:0] s9665, in9665_1, in9665_2;
    wire c9665;
    assign in9665_1 = {c7070};
    assign in9665_2 = {c7071};
    Full_Adder FA_9665(s9665, c9665, in9665_1, in9665_2, c7069);
    wire[0:0] s9666, in9666_1, in9666_2;
    wire c9666;
    assign in9666_1 = {c7073};
    assign in9666_2 = {c7074};
    Full_Adder FA_9666(s9666, c9666, in9666_1, in9666_2, c7072);
    wire[0:0] s9667, in9667_1, in9667_2;
    wire c9667;
    assign in9667_1 = {c7076};
    assign in9667_2 = {c7077};
    Full_Adder FA_9667(s9667, c9667, in9667_1, in9667_2, c7075);
    wire[0:0] s9668, in9668_1, in9668_2;
    wire c9668;
    assign in9668_1 = {c7079};
    assign in9668_2 = {s7080[0]};
    Full_Adder FA_9668(s9668, c9668, in9668_1, in9668_2, c7078);
    wire[0:0] s9669, in9669_1, in9669_2;
    wire c9669;
    assign in9669_1 = {s7082[0]};
    assign in9669_2 = {s7083[0]};
    Full_Adder FA_9669(s9669, c9669, in9669_1, in9669_2, s7081[0]);
    wire[0:0] s9670, in9670_1, in9670_2;
    wire c9670;
    assign in9670_1 = {s7085[0]};
    assign in9670_2 = {s7086[0]};
    Full_Adder FA_9670(s9670, c9670, in9670_1, in9670_2, s7084[0]);
    wire[0:0] s9671, in9671_1, in9671_2;
    wire c9671;
    assign in9671_1 = {s7088[0]};
    assign in9671_2 = {s7089[0]};
    Full_Adder FA_9671(s9671, c9671, in9671_1, in9671_2, s7087[0]);
    wire[0:0] s9672, in9672_1, in9672_2;
    wire c9672;
    assign in9672_1 = {s7091[0]};
    assign in9672_2 = {s7092[0]};
    Full_Adder FA_9672(s9672, c9672, in9672_1, in9672_2, s7090[0]);
    wire[0:0] s9673, in9673_1, in9673_2;
    wire c9673;
    assign in9673_1 = {s7094[0]};
    assign in9673_2 = {s7095[0]};
    Full_Adder FA_9673(s9673, c9673, in9673_1, in9673_2, s7093[0]);
    wire[0:0] s9674, in9674_1, in9674_2;
    wire c9674;
    assign in9674_1 = {s7097[0]};
    assign in9674_2 = {s7098[0]};
    Full_Adder FA_9674(s9674, c9674, in9674_1, in9674_2, s7096[0]);
    wire[0:0] s9675, in9675_1, in9675_2;
    wire c9675;
    assign in9675_1 = {c7080};
    assign in9675_2 = {c7081};
    Full_Adder FA_9675(s9675, c9675, in9675_1, in9675_2, s4312[0]);
    wire[0:0] s9676, in9676_1, in9676_2;
    wire c9676;
    assign in9676_1 = {c7083};
    assign in9676_2 = {c7084};
    Full_Adder FA_9676(s9676, c9676, in9676_1, in9676_2, c7082);
    wire[0:0] s9677, in9677_1, in9677_2;
    wire c9677;
    assign in9677_1 = {c7086};
    assign in9677_2 = {c7087};
    Full_Adder FA_9677(s9677, c9677, in9677_1, in9677_2, c7085);
    wire[0:0] s9678, in9678_1, in9678_2;
    wire c9678;
    assign in9678_1 = {c7089};
    assign in9678_2 = {c7090};
    Full_Adder FA_9678(s9678, c9678, in9678_1, in9678_2, c7088);
    wire[0:0] s9679, in9679_1, in9679_2;
    wire c9679;
    assign in9679_1 = {c7092};
    assign in9679_2 = {c7093};
    Full_Adder FA_9679(s9679, c9679, in9679_1, in9679_2, c7091);
    wire[0:0] s9680, in9680_1, in9680_2;
    wire c9680;
    assign in9680_1 = {c7095};
    assign in9680_2 = {c7096};
    Full_Adder FA_9680(s9680, c9680, in9680_1, in9680_2, c7094);
    wire[0:0] s9681, in9681_1, in9681_2;
    wire c9681;
    assign in9681_1 = {c7098};
    assign in9681_2 = {s7099[0]};
    Full_Adder FA_9681(s9681, c9681, in9681_1, in9681_2, c7097);
    wire[0:0] s9682, in9682_1, in9682_2;
    wire c9682;
    assign in9682_1 = {s7101[0]};
    assign in9682_2 = {s7102[0]};
    Full_Adder FA_9682(s9682, c9682, in9682_1, in9682_2, s7100[0]);
    wire[0:0] s9683, in9683_1, in9683_2;
    wire c9683;
    assign in9683_1 = {s7104[0]};
    assign in9683_2 = {s7105[0]};
    Full_Adder FA_9683(s9683, c9683, in9683_1, in9683_2, s7103[0]);
    wire[0:0] s9684, in9684_1, in9684_2;
    wire c9684;
    assign in9684_1 = {s7107[0]};
    assign in9684_2 = {s7108[0]};
    Full_Adder FA_9684(s9684, c9684, in9684_1, in9684_2, s7106[0]);
    wire[0:0] s9685, in9685_1, in9685_2;
    wire c9685;
    assign in9685_1 = {s7110[0]};
    assign in9685_2 = {s7111[0]};
    Full_Adder FA_9685(s9685, c9685, in9685_1, in9685_2, s7109[0]);
    wire[0:0] s9686, in9686_1, in9686_2;
    wire c9686;
    assign in9686_1 = {s7113[0]};
    assign in9686_2 = {s7114[0]};
    Full_Adder FA_9686(s9686, c9686, in9686_1, in9686_2, s7112[0]);
    wire[0:0] s9687, in9687_1, in9687_2;
    wire c9687;
    assign in9687_1 = {s7116[0]};
    assign in9687_2 = {s7117[0]};
    Full_Adder FA_9687(s9687, c9687, in9687_1, in9687_2, s7115[0]);
    wire[0:0] s9688, in9688_1, in9688_2;
    wire c9688;
    assign in9688_1 = {c7099};
    assign in9688_2 = {c7100};
    Full_Adder FA_9688(s9688, c9688, in9688_1, in9688_2, s4340[0]);
    wire[0:0] s9689, in9689_1, in9689_2;
    wire c9689;
    assign in9689_1 = {c7102};
    assign in9689_2 = {c7103};
    Full_Adder FA_9689(s9689, c9689, in9689_1, in9689_2, c7101);
    wire[0:0] s9690, in9690_1, in9690_2;
    wire c9690;
    assign in9690_1 = {c7105};
    assign in9690_2 = {c7106};
    Full_Adder FA_9690(s9690, c9690, in9690_1, in9690_2, c7104);
    wire[0:0] s9691, in9691_1, in9691_2;
    wire c9691;
    assign in9691_1 = {c7108};
    assign in9691_2 = {c7109};
    Full_Adder FA_9691(s9691, c9691, in9691_1, in9691_2, c7107);
    wire[0:0] s9692, in9692_1, in9692_2;
    wire c9692;
    assign in9692_1 = {c7111};
    assign in9692_2 = {c7112};
    Full_Adder FA_9692(s9692, c9692, in9692_1, in9692_2, c7110);
    wire[0:0] s9693, in9693_1, in9693_2;
    wire c9693;
    assign in9693_1 = {c7114};
    assign in9693_2 = {c7115};
    Full_Adder FA_9693(s9693, c9693, in9693_1, in9693_2, c7113);
    wire[0:0] s9694, in9694_1, in9694_2;
    wire c9694;
    assign in9694_1 = {c7117};
    assign in9694_2 = {s7118[0]};
    Full_Adder FA_9694(s9694, c9694, in9694_1, in9694_2, c7116);
    wire[0:0] s9695, in9695_1, in9695_2;
    wire c9695;
    assign in9695_1 = {s7120[0]};
    assign in9695_2 = {s7121[0]};
    Full_Adder FA_9695(s9695, c9695, in9695_1, in9695_2, s7119[0]);
    wire[0:0] s9696, in9696_1, in9696_2;
    wire c9696;
    assign in9696_1 = {s7123[0]};
    assign in9696_2 = {s7124[0]};
    Full_Adder FA_9696(s9696, c9696, in9696_1, in9696_2, s7122[0]);
    wire[0:0] s9697, in9697_1, in9697_2;
    wire c9697;
    assign in9697_1 = {s7126[0]};
    assign in9697_2 = {s7127[0]};
    Full_Adder FA_9697(s9697, c9697, in9697_1, in9697_2, s7125[0]);
    wire[0:0] s9698, in9698_1, in9698_2;
    wire c9698;
    assign in9698_1 = {s7129[0]};
    assign in9698_2 = {s7130[0]};
    Full_Adder FA_9698(s9698, c9698, in9698_1, in9698_2, s7128[0]);
    wire[0:0] s9699, in9699_1, in9699_2;
    wire c9699;
    assign in9699_1 = {s7132[0]};
    assign in9699_2 = {s7133[0]};
    Full_Adder FA_9699(s9699, c9699, in9699_1, in9699_2, s7131[0]);
    wire[0:0] s9700, in9700_1, in9700_2;
    wire c9700;
    assign in9700_1 = {s7135[0]};
    assign in9700_2 = {s7136[0]};
    Full_Adder FA_9700(s9700, c9700, in9700_1, in9700_2, s7134[0]);
    wire[0:0] s9701, in9701_1, in9701_2;
    wire c9701;
    assign in9701_1 = {c7118};
    assign in9701_2 = {c7119};
    Full_Adder FA_9701(s9701, c9701, in9701_1, in9701_2, s4368[0]);
    wire[0:0] s9702, in9702_1, in9702_2;
    wire c9702;
    assign in9702_1 = {c7121};
    assign in9702_2 = {c7122};
    Full_Adder FA_9702(s9702, c9702, in9702_1, in9702_2, c7120);
    wire[0:0] s9703, in9703_1, in9703_2;
    wire c9703;
    assign in9703_1 = {c7124};
    assign in9703_2 = {c7125};
    Full_Adder FA_9703(s9703, c9703, in9703_1, in9703_2, c7123);
    wire[0:0] s9704, in9704_1, in9704_2;
    wire c9704;
    assign in9704_1 = {c7127};
    assign in9704_2 = {c7128};
    Full_Adder FA_9704(s9704, c9704, in9704_1, in9704_2, c7126);
    wire[0:0] s9705, in9705_1, in9705_2;
    wire c9705;
    assign in9705_1 = {c7130};
    assign in9705_2 = {c7131};
    Full_Adder FA_9705(s9705, c9705, in9705_1, in9705_2, c7129);
    wire[0:0] s9706, in9706_1, in9706_2;
    wire c9706;
    assign in9706_1 = {c7133};
    assign in9706_2 = {c7134};
    Full_Adder FA_9706(s9706, c9706, in9706_1, in9706_2, c7132);
    wire[0:0] s9707, in9707_1, in9707_2;
    wire c9707;
    assign in9707_1 = {c7136};
    assign in9707_2 = {s7137[0]};
    Full_Adder FA_9707(s9707, c9707, in9707_1, in9707_2, c7135);
    wire[0:0] s9708, in9708_1, in9708_2;
    wire c9708;
    assign in9708_1 = {s7139[0]};
    assign in9708_2 = {s7140[0]};
    Full_Adder FA_9708(s9708, c9708, in9708_1, in9708_2, s7138[0]);
    wire[0:0] s9709, in9709_1, in9709_2;
    wire c9709;
    assign in9709_1 = {s7142[0]};
    assign in9709_2 = {s7143[0]};
    Full_Adder FA_9709(s9709, c9709, in9709_1, in9709_2, s7141[0]);
    wire[0:0] s9710, in9710_1, in9710_2;
    wire c9710;
    assign in9710_1 = {s7145[0]};
    assign in9710_2 = {s7146[0]};
    Full_Adder FA_9710(s9710, c9710, in9710_1, in9710_2, s7144[0]);
    wire[0:0] s9711, in9711_1, in9711_2;
    wire c9711;
    assign in9711_1 = {s7148[0]};
    assign in9711_2 = {s7149[0]};
    Full_Adder FA_9711(s9711, c9711, in9711_1, in9711_2, s7147[0]);
    wire[0:0] s9712, in9712_1, in9712_2;
    wire c9712;
    assign in9712_1 = {s7151[0]};
    assign in9712_2 = {s7152[0]};
    Full_Adder FA_9712(s9712, c9712, in9712_1, in9712_2, s7150[0]);
    wire[0:0] s9713, in9713_1, in9713_2;
    wire c9713;
    assign in9713_1 = {s7154[0]};
    assign in9713_2 = {s7155[0]};
    Full_Adder FA_9713(s9713, c9713, in9713_1, in9713_2, s7153[0]);
    wire[0:0] s9714, in9714_1, in9714_2;
    wire c9714;
    assign in9714_1 = {c7137};
    assign in9714_2 = {c7138};
    Full_Adder FA_9714(s9714, c9714, in9714_1, in9714_2, s4396[0]);
    wire[0:0] s9715, in9715_1, in9715_2;
    wire c9715;
    assign in9715_1 = {c7140};
    assign in9715_2 = {c7141};
    Full_Adder FA_9715(s9715, c9715, in9715_1, in9715_2, c7139);
    wire[0:0] s9716, in9716_1, in9716_2;
    wire c9716;
    assign in9716_1 = {c7143};
    assign in9716_2 = {c7144};
    Full_Adder FA_9716(s9716, c9716, in9716_1, in9716_2, c7142);
    wire[0:0] s9717, in9717_1, in9717_2;
    wire c9717;
    assign in9717_1 = {c7146};
    assign in9717_2 = {c7147};
    Full_Adder FA_9717(s9717, c9717, in9717_1, in9717_2, c7145);
    wire[0:0] s9718, in9718_1, in9718_2;
    wire c9718;
    assign in9718_1 = {c7149};
    assign in9718_2 = {c7150};
    Full_Adder FA_9718(s9718, c9718, in9718_1, in9718_2, c7148);
    wire[0:0] s9719, in9719_1, in9719_2;
    wire c9719;
    assign in9719_1 = {c7152};
    assign in9719_2 = {c7153};
    Full_Adder FA_9719(s9719, c9719, in9719_1, in9719_2, c7151);
    wire[0:0] s9720, in9720_1, in9720_2;
    wire c9720;
    assign in9720_1 = {c7155};
    assign in9720_2 = {s7156[0]};
    Full_Adder FA_9720(s9720, c9720, in9720_1, in9720_2, c7154);
    wire[0:0] s9721, in9721_1, in9721_2;
    wire c9721;
    assign in9721_1 = {s7158[0]};
    assign in9721_2 = {s7159[0]};
    Full_Adder FA_9721(s9721, c9721, in9721_1, in9721_2, s7157[0]);
    wire[0:0] s9722, in9722_1, in9722_2;
    wire c9722;
    assign in9722_1 = {s7161[0]};
    assign in9722_2 = {s7162[0]};
    Full_Adder FA_9722(s9722, c9722, in9722_1, in9722_2, s7160[0]);
    wire[0:0] s9723, in9723_1, in9723_2;
    wire c9723;
    assign in9723_1 = {s7164[0]};
    assign in9723_2 = {s7165[0]};
    Full_Adder FA_9723(s9723, c9723, in9723_1, in9723_2, s7163[0]);
    wire[0:0] s9724, in9724_1, in9724_2;
    wire c9724;
    assign in9724_1 = {s7167[0]};
    assign in9724_2 = {s7168[0]};
    Full_Adder FA_9724(s9724, c9724, in9724_1, in9724_2, s7166[0]);
    wire[0:0] s9725, in9725_1, in9725_2;
    wire c9725;
    assign in9725_1 = {s7170[0]};
    assign in9725_2 = {s7171[0]};
    Full_Adder FA_9725(s9725, c9725, in9725_1, in9725_2, s7169[0]);
    wire[0:0] s9726, in9726_1, in9726_2;
    wire c9726;
    assign in9726_1 = {s7173[0]};
    assign in9726_2 = {s7174[0]};
    Full_Adder FA_9726(s9726, c9726, in9726_1, in9726_2, s7172[0]);
    wire[0:0] s9727, in9727_1, in9727_2;
    wire c9727;
    assign in9727_1 = {c7156};
    assign in9727_2 = {c7157};
    Full_Adder FA_9727(s9727, c9727, in9727_1, in9727_2, s4424[0]);
    wire[0:0] s9728, in9728_1, in9728_2;
    wire c9728;
    assign in9728_1 = {c7159};
    assign in9728_2 = {c7160};
    Full_Adder FA_9728(s9728, c9728, in9728_1, in9728_2, c7158);
    wire[0:0] s9729, in9729_1, in9729_2;
    wire c9729;
    assign in9729_1 = {c7162};
    assign in9729_2 = {c7163};
    Full_Adder FA_9729(s9729, c9729, in9729_1, in9729_2, c7161);
    wire[0:0] s9730, in9730_1, in9730_2;
    wire c9730;
    assign in9730_1 = {c7165};
    assign in9730_2 = {c7166};
    Full_Adder FA_9730(s9730, c9730, in9730_1, in9730_2, c7164);
    wire[0:0] s9731, in9731_1, in9731_2;
    wire c9731;
    assign in9731_1 = {c7168};
    assign in9731_2 = {c7169};
    Full_Adder FA_9731(s9731, c9731, in9731_1, in9731_2, c7167);
    wire[0:0] s9732, in9732_1, in9732_2;
    wire c9732;
    assign in9732_1 = {c7171};
    assign in9732_2 = {c7172};
    Full_Adder FA_9732(s9732, c9732, in9732_1, in9732_2, c7170);
    wire[0:0] s9733, in9733_1, in9733_2;
    wire c9733;
    assign in9733_1 = {c7174};
    assign in9733_2 = {s7175[0]};
    Full_Adder FA_9733(s9733, c9733, in9733_1, in9733_2, c7173);
    wire[0:0] s9734, in9734_1, in9734_2;
    wire c9734;
    assign in9734_1 = {s7177[0]};
    assign in9734_2 = {s7178[0]};
    Full_Adder FA_9734(s9734, c9734, in9734_1, in9734_2, s7176[0]);
    wire[0:0] s9735, in9735_1, in9735_2;
    wire c9735;
    assign in9735_1 = {s7180[0]};
    assign in9735_2 = {s7181[0]};
    Full_Adder FA_9735(s9735, c9735, in9735_1, in9735_2, s7179[0]);
    wire[0:0] s9736, in9736_1, in9736_2;
    wire c9736;
    assign in9736_1 = {s7183[0]};
    assign in9736_2 = {s7184[0]};
    Full_Adder FA_9736(s9736, c9736, in9736_1, in9736_2, s7182[0]);
    wire[0:0] s9737, in9737_1, in9737_2;
    wire c9737;
    assign in9737_1 = {s7186[0]};
    assign in9737_2 = {s7187[0]};
    Full_Adder FA_9737(s9737, c9737, in9737_1, in9737_2, s7185[0]);
    wire[0:0] s9738, in9738_1, in9738_2;
    wire c9738;
    assign in9738_1 = {s7189[0]};
    assign in9738_2 = {s7190[0]};
    Full_Adder FA_9738(s9738, c9738, in9738_1, in9738_2, s7188[0]);
    wire[0:0] s9739, in9739_1, in9739_2;
    wire c9739;
    assign in9739_1 = {s7192[0]};
    assign in9739_2 = {s7193[0]};
    Full_Adder FA_9739(s9739, c9739, in9739_1, in9739_2, s7191[0]);
    wire[0:0] s9740, in9740_1, in9740_2;
    wire c9740;
    assign in9740_1 = {c7175};
    assign in9740_2 = {c7176};
    Full_Adder FA_9740(s9740, c9740, in9740_1, in9740_2, s4452[0]);
    wire[0:0] s9741, in9741_1, in9741_2;
    wire c9741;
    assign in9741_1 = {c7178};
    assign in9741_2 = {c7179};
    Full_Adder FA_9741(s9741, c9741, in9741_1, in9741_2, c7177);
    wire[0:0] s9742, in9742_1, in9742_2;
    wire c9742;
    assign in9742_1 = {c7181};
    assign in9742_2 = {c7182};
    Full_Adder FA_9742(s9742, c9742, in9742_1, in9742_2, c7180);
    wire[0:0] s9743, in9743_1, in9743_2;
    wire c9743;
    assign in9743_1 = {c7184};
    assign in9743_2 = {c7185};
    Full_Adder FA_9743(s9743, c9743, in9743_1, in9743_2, c7183);
    wire[0:0] s9744, in9744_1, in9744_2;
    wire c9744;
    assign in9744_1 = {c7187};
    assign in9744_2 = {c7188};
    Full_Adder FA_9744(s9744, c9744, in9744_1, in9744_2, c7186);
    wire[0:0] s9745, in9745_1, in9745_2;
    wire c9745;
    assign in9745_1 = {c7190};
    assign in9745_2 = {c7191};
    Full_Adder FA_9745(s9745, c9745, in9745_1, in9745_2, c7189);
    wire[0:0] s9746, in9746_1, in9746_2;
    wire c9746;
    assign in9746_1 = {c7193};
    assign in9746_2 = {s7194[0]};
    Full_Adder FA_9746(s9746, c9746, in9746_1, in9746_2, c7192);
    wire[0:0] s9747, in9747_1, in9747_2;
    wire c9747;
    assign in9747_1 = {s7196[0]};
    assign in9747_2 = {s7197[0]};
    Full_Adder FA_9747(s9747, c9747, in9747_1, in9747_2, s7195[0]);
    wire[0:0] s9748, in9748_1, in9748_2;
    wire c9748;
    assign in9748_1 = {s7199[0]};
    assign in9748_2 = {s7200[0]};
    Full_Adder FA_9748(s9748, c9748, in9748_1, in9748_2, s7198[0]);
    wire[0:0] s9749, in9749_1, in9749_2;
    wire c9749;
    assign in9749_1 = {s7202[0]};
    assign in9749_2 = {s7203[0]};
    Full_Adder FA_9749(s9749, c9749, in9749_1, in9749_2, s7201[0]);
    wire[0:0] s9750, in9750_1, in9750_2;
    wire c9750;
    assign in9750_1 = {s7205[0]};
    assign in9750_2 = {s7206[0]};
    Full_Adder FA_9750(s9750, c9750, in9750_1, in9750_2, s7204[0]);
    wire[0:0] s9751, in9751_1, in9751_2;
    wire c9751;
    assign in9751_1 = {s7208[0]};
    assign in9751_2 = {s7209[0]};
    Full_Adder FA_9751(s9751, c9751, in9751_1, in9751_2, s7207[0]);
    wire[0:0] s9752, in9752_1, in9752_2;
    wire c9752;
    assign in9752_1 = {s7211[0]};
    assign in9752_2 = {s7212[0]};
    Full_Adder FA_9752(s9752, c9752, in9752_1, in9752_2, s7210[0]);
    wire[0:0] s9753, in9753_1, in9753_2;
    wire c9753;
    assign in9753_1 = {c7194};
    assign in9753_2 = {c7195};
    Full_Adder FA_9753(s9753, c9753, in9753_1, in9753_2, s4480[0]);
    wire[0:0] s9754, in9754_1, in9754_2;
    wire c9754;
    assign in9754_1 = {c7197};
    assign in9754_2 = {c7198};
    Full_Adder FA_9754(s9754, c9754, in9754_1, in9754_2, c7196);
    wire[0:0] s9755, in9755_1, in9755_2;
    wire c9755;
    assign in9755_1 = {c7200};
    assign in9755_2 = {c7201};
    Full_Adder FA_9755(s9755, c9755, in9755_1, in9755_2, c7199);
    wire[0:0] s9756, in9756_1, in9756_2;
    wire c9756;
    assign in9756_1 = {c7203};
    assign in9756_2 = {c7204};
    Full_Adder FA_9756(s9756, c9756, in9756_1, in9756_2, c7202);
    wire[0:0] s9757, in9757_1, in9757_2;
    wire c9757;
    assign in9757_1 = {c7206};
    assign in9757_2 = {c7207};
    Full_Adder FA_9757(s9757, c9757, in9757_1, in9757_2, c7205);
    wire[0:0] s9758, in9758_1, in9758_2;
    wire c9758;
    assign in9758_1 = {c7209};
    assign in9758_2 = {c7210};
    Full_Adder FA_9758(s9758, c9758, in9758_1, in9758_2, c7208);
    wire[0:0] s9759, in9759_1, in9759_2;
    wire c9759;
    assign in9759_1 = {c7212};
    assign in9759_2 = {s7213[0]};
    Full_Adder FA_9759(s9759, c9759, in9759_1, in9759_2, c7211);
    wire[0:0] s9760, in9760_1, in9760_2;
    wire c9760;
    assign in9760_1 = {s7215[0]};
    assign in9760_2 = {s7216[0]};
    Full_Adder FA_9760(s9760, c9760, in9760_1, in9760_2, s7214[0]);
    wire[0:0] s9761, in9761_1, in9761_2;
    wire c9761;
    assign in9761_1 = {s7218[0]};
    assign in9761_2 = {s7219[0]};
    Full_Adder FA_9761(s9761, c9761, in9761_1, in9761_2, s7217[0]);
    wire[0:0] s9762, in9762_1, in9762_2;
    wire c9762;
    assign in9762_1 = {s7221[0]};
    assign in9762_2 = {s7222[0]};
    Full_Adder FA_9762(s9762, c9762, in9762_1, in9762_2, s7220[0]);
    wire[0:0] s9763, in9763_1, in9763_2;
    wire c9763;
    assign in9763_1 = {s7224[0]};
    assign in9763_2 = {s7225[0]};
    Full_Adder FA_9763(s9763, c9763, in9763_1, in9763_2, s7223[0]);
    wire[0:0] s9764, in9764_1, in9764_2;
    wire c9764;
    assign in9764_1 = {s7227[0]};
    assign in9764_2 = {s7228[0]};
    Full_Adder FA_9764(s9764, c9764, in9764_1, in9764_2, s7226[0]);
    wire[0:0] s9765, in9765_1, in9765_2;
    wire c9765;
    assign in9765_1 = {s7230[0]};
    assign in9765_2 = {s7231[0]};
    Full_Adder FA_9765(s9765, c9765, in9765_1, in9765_2, s7229[0]);
    wire[0:0] s9766, in9766_1, in9766_2;
    wire c9766;
    assign in9766_1 = {c7213};
    assign in9766_2 = {c7214};
    Full_Adder FA_9766(s9766, c9766, in9766_1, in9766_2, s4508[0]);
    wire[0:0] s9767, in9767_1, in9767_2;
    wire c9767;
    assign in9767_1 = {c7216};
    assign in9767_2 = {c7217};
    Full_Adder FA_9767(s9767, c9767, in9767_1, in9767_2, c7215);
    wire[0:0] s9768, in9768_1, in9768_2;
    wire c9768;
    assign in9768_1 = {c7219};
    assign in9768_2 = {c7220};
    Full_Adder FA_9768(s9768, c9768, in9768_1, in9768_2, c7218);
    wire[0:0] s9769, in9769_1, in9769_2;
    wire c9769;
    assign in9769_1 = {c7222};
    assign in9769_2 = {c7223};
    Full_Adder FA_9769(s9769, c9769, in9769_1, in9769_2, c7221);
    wire[0:0] s9770, in9770_1, in9770_2;
    wire c9770;
    assign in9770_1 = {c7225};
    assign in9770_2 = {c7226};
    Full_Adder FA_9770(s9770, c9770, in9770_1, in9770_2, c7224);
    wire[0:0] s9771, in9771_1, in9771_2;
    wire c9771;
    assign in9771_1 = {c7228};
    assign in9771_2 = {c7229};
    Full_Adder FA_9771(s9771, c9771, in9771_1, in9771_2, c7227);
    wire[0:0] s9772, in9772_1, in9772_2;
    wire c9772;
    assign in9772_1 = {c7231};
    assign in9772_2 = {s7232[0]};
    Full_Adder FA_9772(s9772, c9772, in9772_1, in9772_2, c7230);
    wire[0:0] s9773, in9773_1, in9773_2;
    wire c9773;
    assign in9773_1 = {s7234[0]};
    assign in9773_2 = {s7235[0]};
    Full_Adder FA_9773(s9773, c9773, in9773_1, in9773_2, s7233[0]);
    wire[0:0] s9774, in9774_1, in9774_2;
    wire c9774;
    assign in9774_1 = {s7237[0]};
    assign in9774_2 = {s7238[0]};
    Full_Adder FA_9774(s9774, c9774, in9774_1, in9774_2, s7236[0]);
    wire[0:0] s9775, in9775_1, in9775_2;
    wire c9775;
    assign in9775_1 = {s7240[0]};
    assign in9775_2 = {s7241[0]};
    Full_Adder FA_9775(s9775, c9775, in9775_1, in9775_2, s7239[0]);
    wire[0:0] s9776, in9776_1, in9776_2;
    wire c9776;
    assign in9776_1 = {s7243[0]};
    assign in9776_2 = {s7244[0]};
    Full_Adder FA_9776(s9776, c9776, in9776_1, in9776_2, s7242[0]);
    wire[0:0] s9777, in9777_1, in9777_2;
    wire c9777;
    assign in9777_1 = {s7246[0]};
    assign in9777_2 = {s7247[0]};
    Full_Adder FA_9777(s9777, c9777, in9777_1, in9777_2, s7245[0]);
    wire[0:0] s9778, in9778_1, in9778_2;
    wire c9778;
    assign in9778_1 = {s7249[0]};
    assign in9778_2 = {s7250[0]};
    Full_Adder FA_9778(s9778, c9778, in9778_1, in9778_2, s7248[0]);
    wire[0:0] s9779, in9779_1, in9779_2;
    wire c9779;
    assign in9779_1 = {c7232};
    assign in9779_2 = {c7233};
    Full_Adder FA_9779(s9779, c9779, in9779_1, in9779_2, s4536[0]);
    wire[0:0] s9780, in9780_1, in9780_2;
    wire c9780;
    assign in9780_1 = {c7235};
    assign in9780_2 = {c7236};
    Full_Adder FA_9780(s9780, c9780, in9780_1, in9780_2, c7234);
    wire[0:0] s9781, in9781_1, in9781_2;
    wire c9781;
    assign in9781_1 = {c7238};
    assign in9781_2 = {c7239};
    Full_Adder FA_9781(s9781, c9781, in9781_1, in9781_2, c7237);
    wire[0:0] s9782, in9782_1, in9782_2;
    wire c9782;
    assign in9782_1 = {c7241};
    assign in9782_2 = {c7242};
    Full_Adder FA_9782(s9782, c9782, in9782_1, in9782_2, c7240);
    wire[0:0] s9783, in9783_1, in9783_2;
    wire c9783;
    assign in9783_1 = {c7244};
    assign in9783_2 = {c7245};
    Full_Adder FA_9783(s9783, c9783, in9783_1, in9783_2, c7243);
    wire[0:0] s9784, in9784_1, in9784_2;
    wire c9784;
    assign in9784_1 = {c7247};
    assign in9784_2 = {c7248};
    Full_Adder FA_9784(s9784, c9784, in9784_1, in9784_2, c7246);
    wire[0:0] s9785, in9785_1, in9785_2;
    wire c9785;
    assign in9785_1 = {c7250};
    assign in9785_2 = {s7251[0]};
    Full_Adder FA_9785(s9785, c9785, in9785_1, in9785_2, c7249);
    wire[0:0] s9786, in9786_1, in9786_2;
    wire c9786;
    assign in9786_1 = {s7253[0]};
    assign in9786_2 = {s7254[0]};
    Full_Adder FA_9786(s9786, c9786, in9786_1, in9786_2, s7252[0]);
    wire[0:0] s9787, in9787_1, in9787_2;
    wire c9787;
    assign in9787_1 = {s7256[0]};
    assign in9787_2 = {s7257[0]};
    Full_Adder FA_9787(s9787, c9787, in9787_1, in9787_2, s7255[0]);
    wire[0:0] s9788, in9788_1, in9788_2;
    wire c9788;
    assign in9788_1 = {s7259[0]};
    assign in9788_2 = {s7260[0]};
    Full_Adder FA_9788(s9788, c9788, in9788_1, in9788_2, s7258[0]);
    wire[0:0] s9789, in9789_1, in9789_2;
    wire c9789;
    assign in9789_1 = {s7262[0]};
    assign in9789_2 = {s7263[0]};
    Full_Adder FA_9789(s9789, c9789, in9789_1, in9789_2, s7261[0]);
    wire[0:0] s9790, in9790_1, in9790_2;
    wire c9790;
    assign in9790_1 = {s7265[0]};
    assign in9790_2 = {s7266[0]};
    Full_Adder FA_9790(s9790, c9790, in9790_1, in9790_2, s7264[0]);
    wire[0:0] s9791, in9791_1, in9791_2;
    wire c9791;
    assign in9791_1 = {s7268[0]};
    assign in9791_2 = {s7269[0]};
    Full_Adder FA_9791(s9791, c9791, in9791_1, in9791_2, s7267[0]);
    wire[0:0] s9792, in9792_1, in9792_2;
    wire c9792;
    assign in9792_1 = {c7251};
    assign in9792_2 = {c7252};
    Full_Adder FA_9792(s9792, c9792, in9792_1, in9792_2, s4564[0]);
    wire[0:0] s9793, in9793_1, in9793_2;
    wire c9793;
    assign in9793_1 = {c7254};
    assign in9793_2 = {c7255};
    Full_Adder FA_9793(s9793, c9793, in9793_1, in9793_2, c7253);
    wire[0:0] s9794, in9794_1, in9794_2;
    wire c9794;
    assign in9794_1 = {c7257};
    assign in9794_2 = {c7258};
    Full_Adder FA_9794(s9794, c9794, in9794_1, in9794_2, c7256);
    wire[0:0] s9795, in9795_1, in9795_2;
    wire c9795;
    assign in9795_1 = {c7260};
    assign in9795_2 = {c7261};
    Full_Adder FA_9795(s9795, c9795, in9795_1, in9795_2, c7259);
    wire[0:0] s9796, in9796_1, in9796_2;
    wire c9796;
    assign in9796_1 = {c7263};
    assign in9796_2 = {c7264};
    Full_Adder FA_9796(s9796, c9796, in9796_1, in9796_2, c7262);
    wire[0:0] s9797, in9797_1, in9797_2;
    wire c9797;
    assign in9797_1 = {c7266};
    assign in9797_2 = {c7267};
    Full_Adder FA_9797(s9797, c9797, in9797_1, in9797_2, c7265);
    wire[0:0] s9798, in9798_1, in9798_2;
    wire c9798;
    assign in9798_1 = {c7269};
    assign in9798_2 = {s7270[0]};
    Full_Adder FA_9798(s9798, c9798, in9798_1, in9798_2, c7268);
    wire[0:0] s9799, in9799_1, in9799_2;
    wire c9799;
    assign in9799_1 = {s7272[0]};
    assign in9799_2 = {s7273[0]};
    Full_Adder FA_9799(s9799, c9799, in9799_1, in9799_2, s7271[0]);
    wire[0:0] s9800, in9800_1, in9800_2;
    wire c9800;
    assign in9800_1 = {s7275[0]};
    assign in9800_2 = {s7276[0]};
    Full_Adder FA_9800(s9800, c9800, in9800_1, in9800_2, s7274[0]);
    wire[0:0] s9801, in9801_1, in9801_2;
    wire c9801;
    assign in9801_1 = {s7278[0]};
    assign in9801_2 = {s7279[0]};
    Full_Adder FA_9801(s9801, c9801, in9801_1, in9801_2, s7277[0]);
    wire[0:0] s9802, in9802_1, in9802_2;
    wire c9802;
    assign in9802_1 = {s7281[0]};
    assign in9802_2 = {s7282[0]};
    Full_Adder FA_9802(s9802, c9802, in9802_1, in9802_2, s7280[0]);
    wire[0:0] s9803, in9803_1, in9803_2;
    wire c9803;
    assign in9803_1 = {s7284[0]};
    assign in9803_2 = {s7285[0]};
    Full_Adder FA_9803(s9803, c9803, in9803_1, in9803_2, s7283[0]);
    wire[0:0] s9804, in9804_1, in9804_2;
    wire c9804;
    assign in9804_1 = {s7287[0]};
    assign in9804_2 = {s7288[0]};
    Full_Adder FA_9804(s9804, c9804, in9804_1, in9804_2, s7286[0]);
    wire[0:0] s9805, in9805_1, in9805_2;
    wire c9805;
    assign in9805_1 = {c7270};
    assign in9805_2 = {c7271};
    Full_Adder FA_9805(s9805, c9805, in9805_1, in9805_2, s4592[0]);
    wire[0:0] s9806, in9806_1, in9806_2;
    wire c9806;
    assign in9806_1 = {c7273};
    assign in9806_2 = {c7274};
    Full_Adder FA_9806(s9806, c9806, in9806_1, in9806_2, c7272);
    wire[0:0] s9807, in9807_1, in9807_2;
    wire c9807;
    assign in9807_1 = {c7276};
    assign in9807_2 = {c7277};
    Full_Adder FA_9807(s9807, c9807, in9807_1, in9807_2, c7275);
    wire[0:0] s9808, in9808_1, in9808_2;
    wire c9808;
    assign in9808_1 = {c7279};
    assign in9808_2 = {c7280};
    Full_Adder FA_9808(s9808, c9808, in9808_1, in9808_2, c7278);
    wire[0:0] s9809, in9809_1, in9809_2;
    wire c9809;
    assign in9809_1 = {c7282};
    assign in9809_2 = {c7283};
    Full_Adder FA_9809(s9809, c9809, in9809_1, in9809_2, c7281);
    wire[0:0] s9810, in9810_1, in9810_2;
    wire c9810;
    assign in9810_1 = {c7285};
    assign in9810_2 = {c7286};
    Full_Adder FA_9810(s9810, c9810, in9810_1, in9810_2, c7284);
    wire[0:0] s9811, in9811_1, in9811_2;
    wire c9811;
    assign in9811_1 = {c7288};
    assign in9811_2 = {s7289[0]};
    Full_Adder FA_9811(s9811, c9811, in9811_1, in9811_2, c7287);
    wire[0:0] s9812, in9812_1, in9812_2;
    wire c9812;
    assign in9812_1 = {s7291[0]};
    assign in9812_2 = {s7292[0]};
    Full_Adder FA_9812(s9812, c9812, in9812_1, in9812_2, s7290[0]);
    wire[0:0] s9813, in9813_1, in9813_2;
    wire c9813;
    assign in9813_1 = {s7294[0]};
    assign in9813_2 = {s7295[0]};
    Full_Adder FA_9813(s9813, c9813, in9813_1, in9813_2, s7293[0]);
    wire[0:0] s9814, in9814_1, in9814_2;
    wire c9814;
    assign in9814_1 = {s7297[0]};
    assign in9814_2 = {s7298[0]};
    Full_Adder FA_9814(s9814, c9814, in9814_1, in9814_2, s7296[0]);
    wire[0:0] s9815, in9815_1, in9815_2;
    wire c9815;
    assign in9815_1 = {s7300[0]};
    assign in9815_2 = {s7301[0]};
    Full_Adder FA_9815(s9815, c9815, in9815_1, in9815_2, s7299[0]);
    wire[0:0] s9816, in9816_1, in9816_2;
    wire c9816;
    assign in9816_1 = {s7303[0]};
    assign in9816_2 = {s7304[0]};
    Full_Adder FA_9816(s9816, c9816, in9816_1, in9816_2, s7302[0]);
    wire[0:0] s9817, in9817_1, in9817_2;
    wire c9817;
    assign in9817_1 = {s7306[0]};
    assign in9817_2 = {s7307[0]};
    Full_Adder FA_9817(s9817, c9817, in9817_1, in9817_2, s7305[0]);
    wire[0:0] s9818, in9818_1, in9818_2;
    wire c9818;
    assign in9818_1 = {c7289};
    assign in9818_2 = {c7290};
    Full_Adder FA_9818(s9818, c9818, in9818_1, in9818_2, s4619[0]);
    wire[0:0] s9819, in9819_1, in9819_2;
    wire c9819;
    assign in9819_1 = {c7292};
    assign in9819_2 = {c7293};
    Full_Adder FA_9819(s9819, c9819, in9819_1, in9819_2, c7291);
    wire[0:0] s9820, in9820_1, in9820_2;
    wire c9820;
    assign in9820_1 = {c7295};
    assign in9820_2 = {c7296};
    Full_Adder FA_9820(s9820, c9820, in9820_1, in9820_2, c7294);
    wire[0:0] s9821, in9821_1, in9821_2;
    wire c9821;
    assign in9821_1 = {c7298};
    assign in9821_2 = {c7299};
    Full_Adder FA_9821(s9821, c9821, in9821_1, in9821_2, c7297);
    wire[0:0] s9822, in9822_1, in9822_2;
    wire c9822;
    assign in9822_1 = {c7301};
    assign in9822_2 = {c7302};
    Full_Adder FA_9822(s9822, c9822, in9822_1, in9822_2, c7300);
    wire[0:0] s9823, in9823_1, in9823_2;
    wire c9823;
    assign in9823_1 = {c7304};
    assign in9823_2 = {c7305};
    Full_Adder FA_9823(s9823, c9823, in9823_1, in9823_2, c7303);
    wire[0:0] s9824, in9824_1, in9824_2;
    wire c9824;
    assign in9824_1 = {c7307};
    assign in9824_2 = {s7308[0]};
    Full_Adder FA_9824(s9824, c9824, in9824_1, in9824_2, c7306);
    wire[0:0] s9825, in9825_1, in9825_2;
    wire c9825;
    assign in9825_1 = {s7310[0]};
    assign in9825_2 = {s7311[0]};
    Full_Adder FA_9825(s9825, c9825, in9825_1, in9825_2, s7309[0]);
    wire[0:0] s9826, in9826_1, in9826_2;
    wire c9826;
    assign in9826_1 = {s7313[0]};
    assign in9826_2 = {s7314[0]};
    Full_Adder FA_9826(s9826, c9826, in9826_1, in9826_2, s7312[0]);
    wire[0:0] s9827, in9827_1, in9827_2;
    wire c9827;
    assign in9827_1 = {s7316[0]};
    assign in9827_2 = {s7317[0]};
    Full_Adder FA_9827(s9827, c9827, in9827_1, in9827_2, s7315[0]);
    wire[0:0] s9828, in9828_1, in9828_2;
    wire c9828;
    assign in9828_1 = {s7319[0]};
    assign in9828_2 = {s7320[0]};
    Full_Adder FA_9828(s9828, c9828, in9828_1, in9828_2, s7318[0]);
    wire[0:0] s9829, in9829_1, in9829_2;
    wire c9829;
    assign in9829_1 = {s7322[0]};
    assign in9829_2 = {s7323[0]};
    Full_Adder FA_9829(s9829, c9829, in9829_1, in9829_2, s7321[0]);
    wire[0:0] s9830, in9830_1, in9830_2;
    wire c9830;
    assign in9830_1 = {s7325[0]};
    assign in9830_2 = {s7326[0]};
    Full_Adder FA_9830(s9830, c9830, in9830_1, in9830_2, s7324[0]);
    wire[0:0] s9831, in9831_1, in9831_2;
    wire c9831;
    assign in9831_1 = {c7308};
    assign in9831_2 = {c7309};
    Full_Adder FA_9831(s9831, c9831, in9831_1, in9831_2, s4645[0]);
    wire[0:0] s9832, in9832_1, in9832_2;
    wire c9832;
    assign in9832_1 = {c7311};
    assign in9832_2 = {c7312};
    Full_Adder FA_9832(s9832, c9832, in9832_1, in9832_2, c7310);
    wire[0:0] s9833, in9833_1, in9833_2;
    wire c9833;
    assign in9833_1 = {c7314};
    assign in9833_2 = {c7315};
    Full_Adder FA_9833(s9833, c9833, in9833_1, in9833_2, c7313);
    wire[0:0] s9834, in9834_1, in9834_2;
    wire c9834;
    assign in9834_1 = {c7317};
    assign in9834_2 = {c7318};
    Full_Adder FA_9834(s9834, c9834, in9834_1, in9834_2, c7316);
    wire[0:0] s9835, in9835_1, in9835_2;
    wire c9835;
    assign in9835_1 = {c7320};
    assign in9835_2 = {c7321};
    Full_Adder FA_9835(s9835, c9835, in9835_1, in9835_2, c7319);
    wire[0:0] s9836, in9836_1, in9836_2;
    wire c9836;
    assign in9836_1 = {c7323};
    assign in9836_2 = {c7324};
    Full_Adder FA_9836(s9836, c9836, in9836_1, in9836_2, c7322);
    wire[0:0] s9837, in9837_1, in9837_2;
    wire c9837;
    assign in9837_1 = {c7326};
    assign in9837_2 = {s7327[0]};
    Full_Adder FA_9837(s9837, c9837, in9837_1, in9837_2, c7325);
    wire[0:0] s9838, in9838_1, in9838_2;
    wire c9838;
    assign in9838_1 = {s7329[0]};
    assign in9838_2 = {s7330[0]};
    Full_Adder FA_9838(s9838, c9838, in9838_1, in9838_2, s7328[0]);
    wire[0:0] s9839, in9839_1, in9839_2;
    wire c9839;
    assign in9839_1 = {s7332[0]};
    assign in9839_2 = {s7333[0]};
    Full_Adder FA_9839(s9839, c9839, in9839_1, in9839_2, s7331[0]);
    wire[0:0] s9840, in9840_1, in9840_2;
    wire c9840;
    assign in9840_1 = {s7335[0]};
    assign in9840_2 = {s7336[0]};
    Full_Adder FA_9840(s9840, c9840, in9840_1, in9840_2, s7334[0]);
    wire[0:0] s9841, in9841_1, in9841_2;
    wire c9841;
    assign in9841_1 = {s7338[0]};
    assign in9841_2 = {s7339[0]};
    Full_Adder FA_9841(s9841, c9841, in9841_1, in9841_2, s7337[0]);
    wire[0:0] s9842, in9842_1, in9842_2;
    wire c9842;
    assign in9842_1 = {s7341[0]};
    assign in9842_2 = {s7342[0]};
    Full_Adder FA_9842(s9842, c9842, in9842_1, in9842_2, s7340[0]);
    wire[0:0] s9843, in9843_1, in9843_2;
    wire c9843;
    assign in9843_1 = {s7344[0]};
    assign in9843_2 = {s7345[0]};
    Full_Adder FA_9843(s9843, c9843, in9843_1, in9843_2, s7343[0]);
    wire[0:0] s9844, in9844_1, in9844_2;
    wire c9844;
    assign in9844_1 = {c7327};
    assign in9844_2 = {c7328};
    Full_Adder FA_9844(s9844, c9844, in9844_1, in9844_2, s4670[0]);
    wire[0:0] s9845, in9845_1, in9845_2;
    wire c9845;
    assign in9845_1 = {c7330};
    assign in9845_2 = {c7331};
    Full_Adder FA_9845(s9845, c9845, in9845_1, in9845_2, c7329);
    wire[0:0] s9846, in9846_1, in9846_2;
    wire c9846;
    assign in9846_1 = {c7333};
    assign in9846_2 = {c7334};
    Full_Adder FA_9846(s9846, c9846, in9846_1, in9846_2, c7332);
    wire[0:0] s9847, in9847_1, in9847_2;
    wire c9847;
    assign in9847_1 = {c7336};
    assign in9847_2 = {c7337};
    Full_Adder FA_9847(s9847, c9847, in9847_1, in9847_2, c7335);
    wire[0:0] s9848, in9848_1, in9848_2;
    wire c9848;
    assign in9848_1 = {c7339};
    assign in9848_2 = {c7340};
    Full_Adder FA_9848(s9848, c9848, in9848_1, in9848_2, c7338);
    wire[0:0] s9849, in9849_1, in9849_2;
    wire c9849;
    assign in9849_1 = {c7342};
    assign in9849_2 = {c7343};
    Full_Adder FA_9849(s9849, c9849, in9849_1, in9849_2, c7341);
    wire[0:0] s9850, in9850_1, in9850_2;
    wire c9850;
    assign in9850_1 = {c7345};
    assign in9850_2 = {s7346[0]};
    Full_Adder FA_9850(s9850, c9850, in9850_1, in9850_2, c7344);
    wire[0:0] s9851, in9851_1, in9851_2;
    wire c9851;
    assign in9851_1 = {s7348[0]};
    assign in9851_2 = {s7349[0]};
    Full_Adder FA_9851(s9851, c9851, in9851_1, in9851_2, s7347[0]);
    wire[0:0] s9852, in9852_1, in9852_2;
    wire c9852;
    assign in9852_1 = {s7351[0]};
    assign in9852_2 = {s7352[0]};
    Full_Adder FA_9852(s9852, c9852, in9852_1, in9852_2, s7350[0]);
    wire[0:0] s9853, in9853_1, in9853_2;
    wire c9853;
    assign in9853_1 = {s7354[0]};
    assign in9853_2 = {s7355[0]};
    Full_Adder FA_9853(s9853, c9853, in9853_1, in9853_2, s7353[0]);
    wire[0:0] s9854, in9854_1, in9854_2;
    wire c9854;
    assign in9854_1 = {s7357[0]};
    assign in9854_2 = {s7358[0]};
    Full_Adder FA_9854(s9854, c9854, in9854_1, in9854_2, s7356[0]);
    wire[0:0] s9855, in9855_1, in9855_2;
    wire c9855;
    assign in9855_1 = {s7360[0]};
    assign in9855_2 = {s7361[0]};
    Full_Adder FA_9855(s9855, c9855, in9855_1, in9855_2, s7359[0]);
    wire[0:0] s9856, in9856_1, in9856_2;
    wire c9856;
    assign in9856_1 = {s7363[0]};
    assign in9856_2 = {s7364[0]};
    Full_Adder FA_9856(s9856, c9856, in9856_1, in9856_2, s7362[0]);
    wire[0:0] s9857, in9857_1, in9857_2;
    wire c9857;
    assign in9857_1 = {c7346};
    assign in9857_2 = {c7347};
    Full_Adder FA_9857(s9857, c9857, in9857_1, in9857_2, s4694[0]);
    wire[0:0] s9858, in9858_1, in9858_2;
    wire c9858;
    assign in9858_1 = {c7349};
    assign in9858_2 = {c7350};
    Full_Adder FA_9858(s9858, c9858, in9858_1, in9858_2, c7348);
    wire[0:0] s9859, in9859_1, in9859_2;
    wire c9859;
    assign in9859_1 = {c7352};
    assign in9859_2 = {c7353};
    Full_Adder FA_9859(s9859, c9859, in9859_1, in9859_2, c7351);
    wire[0:0] s9860, in9860_1, in9860_2;
    wire c9860;
    assign in9860_1 = {c7355};
    assign in9860_2 = {c7356};
    Full_Adder FA_9860(s9860, c9860, in9860_1, in9860_2, c7354);
    wire[0:0] s9861, in9861_1, in9861_2;
    wire c9861;
    assign in9861_1 = {c7358};
    assign in9861_2 = {c7359};
    Full_Adder FA_9861(s9861, c9861, in9861_1, in9861_2, c7357);
    wire[0:0] s9862, in9862_1, in9862_2;
    wire c9862;
    assign in9862_1 = {c7361};
    assign in9862_2 = {c7362};
    Full_Adder FA_9862(s9862, c9862, in9862_1, in9862_2, c7360);
    wire[0:0] s9863, in9863_1, in9863_2;
    wire c9863;
    assign in9863_1 = {c7364};
    assign in9863_2 = {s7365[0]};
    Full_Adder FA_9863(s9863, c9863, in9863_1, in9863_2, c7363);
    wire[0:0] s9864, in9864_1, in9864_2;
    wire c9864;
    assign in9864_1 = {s7367[0]};
    assign in9864_2 = {s7368[0]};
    Full_Adder FA_9864(s9864, c9864, in9864_1, in9864_2, s7366[0]);
    wire[0:0] s9865, in9865_1, in9865_2;
    wire c9865;
    assign in9865_1 = {s7370[0]};
    assign in9865_2 = {s7371[0]};
    Full_Adder FA_9865(s9865, c9865, in9865_1, in9865_2, s7369[0]);
    wire[0:0] s9866, in9866_1, in9866_2;
    wire c9866;
    assign in9866_1 = {s7373[0]};
    assign in9866_2 = {s7374[0]};
    Full_Adder FA_9866(s9866, c9866, in9866_1, in9866_2, s7372[0]);
    wire[0:0] s9867, in9867_1, in9867_2;
    wire c9867;
    assign in9867_1 = {s7376[0]};
    assign in9867_2 = {s7377[0]};
    Full_Adder FA_9867(s9867, c9867, in9867_1, in9867_2, s7375[0]);
    wire[0:0] s9868, in9868_1, in9868_2;
    wire c9868;
    assign in9868_1 = {s7379[0]};
    assign in9868_2 = {s7380[0]};
    Full_Adder FA_9868(s9868, c9868, in9868_1, in9868_2, s7378[0]);
    wire[0:0] s9869, in9869_1, in9869_2;
    wire c9869;
    assign in9869_1 = {s7382[0]};
    assign in9869_2 = {s7383[0]};
    Full_Adder FA_9869(s9869, c9869, in9869_1, in9869_2, s7381[0]);
    wire[0:0] s9870, in9870_1, in9870_2;
    wire c9870;
    assign in9870_1 = {c7365};
    assign in9870_2 = {c7366};
    Full_Adder FA_9870(s9870, c9870, in9870_1, in9870_2, s4717[0]);
    wire[0:0] s9871, in9871_1, in9871_2;
    wire c9871;
    assign in9871_1 = {c7368};
    assign in9871_2 = {c7369};
    Full_Adder FA_9871(s9871, c9871, in9871_1, in9871_2, c7367);
    wire[0:0] s9872, in9872_1, in9872_2;
    wire c9872;
    assign in9872_1 = {c7371};
    assign in9872_2 = {c7372};
    Full_Adder FA_9872(s9872, c9872, in9872_1, in9872_2, c7370);
    wire[0:0] s9873, in9873_1, in9873_2;
    wire c9873;
    assign in9873_1 = {c7374};
    assign in9873_2 = {c7375};
    Full_Adder FA_9873(s9873, c9873, in9873_1, in9873_2, c7373);
    wire[0:0] s9874, in9874_1, in9874_2;
    wire c9874;
    assign in9874_1 = {c7377};
    assign in9874_2 = {c7378};
    Full_Adder FA_9874(s9874, c9874, in9874_1, in9874_2, c7376);
    wire[0:0] s9875, in9875_1, in9875_2;
    wire c9875;
    assign in9875_1 = {c7380};
    assign in9875_2 = {c7381};
    Full_Adder FA_9875(s9875, c9875, in9875_1, in9875_2, c7379);
    wire[0:0] s9876, in9876_1, in9876_2;
    wire c9876;
    assign in9876_1 = {c7383};
    assign in9876_2 = {s7384[0]};
    Full_Adder FA_9876(s9876, c9876, in9876_1, in9876_2, c7382);
    wire[0:0] s9877, in9877_1, in9877_2;
    wire c9877;
    assign in9877_1 = {s7386[0]};
    assign in9877_2 = {s7387[0]};
    Full_Adder FA_9877(s9877, c9877, in9877_1, in9877_2, s7385[0]);
    wire[0:0] s9878, in9878_1, in9878_2;
    wire c9878;
    assign in9878_1 = {s7389[0]};
    assign in9878_2 = {s7390[0]};
    Full_Adder FA_9878(s9878, c9878, in9878_1, in9878_2, s7388[0]);
    wire[0:0] s9879, in9879_1, in9879_2;
    wire c9879;
    assign in9879_1 = {s7392[0]};
    assign in9879_2 = {s7393[0]};
    Full_Adder FA_9879(s9879, c9879, in9879_1, in9879_2, s7391[0]);
    wire[0:0] s9880, in9880_1, in9880_2;
    wire c9880;
    assign in9880_1 = {s7395[0]};
    assign in9880_2 = {s7396[0]};
    Full_Adder FA_9880(s9880, c9880, in9880_1, in9880_2, s7394[0]);
    wire[0:0] s9881, in9881_1, in9881_2;
    wire c9881;
    assign in9881_1 = {s7398[0]};
    assign in9881_2 = {s7399[0]};
    Full_Adder FA_9881(s9881, c9881, in9881_1, in9881_2, s7397[0]);
    wire[0:0] s9882, in9882_1, in9882_2;
    wire c9882;
    assign in9882_1 = {s7401[0]};
    assign in9882_2 = {s7402[0]};
    Full_Adder FA_9882(s9882, c9882, in9882_1, in9882_2, s7400[0]);
    wire[0:0] s9883, in9883_1, in9883_2;
    wire c9883;
    assign in9883_1 = {c7384};
    assign in9883_2 = {c7385};
    Full_Adder FA_9883(s9883, c9883, in9883_1, in9883_2, s4739[0]);
    wire[0:0] s9884, in9884_1, in9884_2;
    wire c9884;
    assign in9884_1 = {c7387};
    assign in9884_2 = {c7388};
    Full_Adder FA_9884(s9884, c9884, in9884_1, in9884_2, c7386);
    wire[0:0] s9885, in9885_1, in9885_2;
    wire c9885;
    assign in9885_1 = {c7390};
    assign in9885_2 = {c7391};
    Full_Adder FA_9885(s9885, c9885, in9885_1, in9885_2, c7389);
    wire[0:0] s9886, in9886_1, in9886_2;
    wire c9886;
    assign in9886_1 = {c7393};
    assign in9886_2 = {c7394};
    Full_Adder FA_9886(s9886, c9886, in9886_1, in9886_2, c7392);
    wire[0:0] s9887, in9887_1, in9887_2;
    wire c9887;
    assign in9887_1 = {c7396};
    assign in9887_2 = {c7397};
    Full_Adder FA_9887(s9887, c9887, in9887_1, in9887_2, c7395);
    wire[0:0] s9888, in9888_1, in9888_2;
    wire c9888;
    assign in9888_1 = {c7399};
    assign in9888_2 = {c7400};
    Full_Adder FA_9888(s9888, c9888, in9888_1, in9888_2, c7398);
    wire[0:0] s9889, in9889_1, in9889_2;
    wire c9889;
    assign in9889_1 = {c7402};
    assign in9889_2 = {s7403[0]};
    Full_Adder FA_9889(s9889, c9889, in9889_1, in9889_2, c7401);
    wire[0:0] s9890, in9890_1, in9890_2;
    wire c9890;
    assign in9890_1 = {s7405[0]};
    assign in9890_2 = {s7406[0]};
    Full_Adder FA_9890(s9890, c9890, in9890_1, in9890_2, s7404[0]);
    wire[0:0] s9891, in9891_1, in9891_2;
    wire c9891;
    assign in9891_1 = {s7408[0]};
    assign in9891_2 = {s7409[0]};
    Full_Adder FA_9891(s9891, c9891, in9891_1, in9891_2, s7407[0]);
    wire[0:0] s9892, in9892_1, in9892_2;
    wire c9892;
    assign in9892_1 = {s7411[0]};
    assign in9892_2 = {s7412[0]};
    Full_Adder FA_9892(s9892, c9892, in9892_1, in9892_2, s7410[0]);
    wire[0:0] s9893, in9893_1, in9893_2;
    wire c9893;
    assign in9893_1 = {s7414[0]};
    assign in9893_2 = {s7415[0]};
    Full_Adder FA_9893(s9893, c9893, in9893_1, in9893_2, s7413[0]);
    wire[0:0] s9894, in9894_1, in9894_2;
    wire c9894;
    assign in9894_1 = {s7417[0]};
    assign in9894_2 = {s7418[0]};
    Full_Adder FA_9894(s9894, c9894, in9894_1, in9894_2, s7416[0]);
    wire[0:0] s9895, in9895_1, in9895_2;
    wire c9895;
    assign in9895_1 = {s7420[0]};
    assign in9895_2 = {s7421[0]};
    Full_Adder FA_9895(s9895, c9895, in9895_1, in9895_2, s7419[0]);
    wire[0:0] s9896, in9896_1, in9896_2;
    wire c9896;
    assign in9896_1 = {c7403};
    assign in9896_2 = {c7404};
    Full_Adder FA_9896(s9896, c9896, in9896_1, in9896_2, s4760[0]);
    wire[0:0] s9897, in9897_1, in9897_2;
    wire c9897;
    assign in9897_1 = {c7406};
    assign in9897_2 = {c7407};
    Full_Adder FA_9897(s9897, c9897, in9897_1, in9897_2, c7405);
    wire[0:0] s9898, in9898_1, in9898_2;
    wire c9898;
    assign in9898_1 = {c7409};
    assign in9898_2 = {c7410};
    Full_Adder FA_9898(s9898, c9898, in9898_1, in9898_2, c7408);
    wire[0:0] s9899, in9899_1, in9899_2;
    wire c9899;
    assign in9899_1 = {c7412};
    assign in9899_2 = {c7413};
    Full_Adder FA_9899(s9899, c9899, in9899_1, in9899_2, c7411);
    wire[0:0] s9900, in9900_1, in9900_2;
    wire c9900;
    assign in9900_1 = {c7415};
    assign in9900_2 = {c7416};
    Full_Adder FA_9900(s9900, c9900, in9900_1, in9900_2, c7414);
    wire[0:0] s9901, in9901_1, in9901_2;
    wire c9901;
    assign in9901_1 = {c7418};
    assign in9901_2 = {c7419};
    Full_Adder FA_9901(s9901, c9901, in9901_1, in9901_2, c7417);
    wire[0:0] s9902, in9902_1, in9902_2;
    wire c9902;
    assign in9902_1 = {c7421};
    assign in9902_2 = {s7422[0]};
    Full_Adder FA_9902(s9902, c9902, in9902_1, in9902_2, c7420);
    wire[0:0] s9903, in9903_1, in9903_2;
    wire c9903;
    assign in9903_1 = {s7424[0]};
    assign in9903_2 = {s7425[0]};
    Full_Adder FA_9903(s9903, c9903, in9903_1, in9903_2, s7423[0]);
    wire[0:0] s9904, in9904_1, in9904_2;
    wire c9904;
    assign in9904_1 = {s7427[0]};
    assign in9904_2 = {s7428[0]};
    Full_Adder FA_9904(s9904, c9904, in9904_1, in9904_2, s7426[0]);
    wire[0:0] s9905, in9905_1, in9905_2;
    wire c9905;
    assign in9905_1 = {s7430[0]};
    assign in9905_2 = {s7431[0]};
    Full_Adder FA_9905(s9905, c9905, in9905_1, in9905_2, s7429[0]);
    wire[0:0] s9906, in9906_1, in9906_2;
    wire c9906;
    assign in9906_1 = {s7433[0]};
    assign in9906_2 = {s7434[0]};
    Full_Adder FA_9906(s9906, c9906, in9906_1, in9906_2, s7432[0]);
    wire[0:0] s9907, in9907_1, in9907_2;
    wire c9907;
    assign in9907_1 = {s7436[0]};
    assign in9907_2 = {s7437[0]};
    Full_Adder FA_9907(s9907, c9907, in9907_1, in9907_2, s7435[0]);
    wire[0:0] s9908, in9908_1, in9908_2;
    wire c9908;
    assign in9908_1 = {s7439[0]};
    assign in9908_2 = {s7440[0]};
    Full_Adder FA_9908(s9908, c9908, in9908_1, in9908_2, s7438[0]);
    wire[0:0] s9909, in9909_1, in9909_2;
    wire c9909;
    assign in9909_1 = {c7422};
    assign in9909_2 = {c7423};
    Full_Adder FA_9909(s9909, c9909, in9909_1, in9909_2, s4780[0]);
    wire[0:0] s9910, in9910_1, in9910_2;
    wire c9910;
    assign in9910_1 = {c7425};
    assign in9910_2 = {c7426};
    Full_Adder FA_9910(s9910, c9910, in9910_1, in9910_2, c7424);
    wire[0:0] s9911, in9911_1, in9911_2;
    wire c9911;
    assign in9911_1 = {c7428};
    assign in9911_2 = {c7429};
    Full_Adder FA_9911(s9911, c9911, in9911_1, in9911_2, c7427);
    wire[0:0] s9912, in9912_1, in9912_2;
    wire c9912;
    assign in9912_1 = {c7431};
    assign in9912_2 = {c7432};
    Full_Adder FA_9912(s9912, c9912, in9912_1, in9912_2, c7430);
    wire[0:0] s9913, in9913_1, in9913_2;
    wire c9913;
    assign in9913_1 = {c7434};
    assign in9913_2 = {c7435};
    Full_Adder FA_9913(s9913, c9913, in9913_1, in9913_2, c7433);
    wire[0:0] s9914, in9914_1, in9914_2;
    wire c9914;
    assign in9914_1 = {c7437};
    assign in9914_2 = {c7438};
    Full_Adder FA_9914(s9914, c9914, in9914_1, in9914_2, c7436);
    wire[0:0] s9915, in9915_1, in9915_2;
    wire c9915;
    assign in9915_1 = {c7440};
    assign in9915_2 = {s7441[0]};
    Full_Adder FA_9915(s9915, c9915, in9915_1, in9915_2, c7439);
    wire[0:0] s9916, in9916_1, in9916_2;
    wire c9916;
    assign in9916_1 = {s7443[0]};
    assign in9916_2 = {s7444[0]};
    Full_Adder FA_9916(s9916, c9916, in9916_1, in9916_2, s7442[0]);
    wire[0:0] s9917, in9917_1, in9917_2;
    wire c9917;
    assign in9917_1 = {s7446[0]};
    assign in9917_2 = {s7447[0]};
    Full_Adder FA_9917(s9917, c9917, in9917_1, in9917_2, s7445[0]);
    wire[0:0] s9918, in9918_1, in9918_2;
    wire c9918;
    assign in9918_1 = {s7449[0]};
    assign in9918_2 = {s7450[0]};
    Full_Adder FA_9918(s9918, c9918, in9918_1, in9918_2, s7448[0]);
    wire[0:0] s9919, in9919_1, in9919_2;
    wire c9919;
    assign in9919_1 = {s7452[0]};
    assign in9919_2 = {s7453[0]};
    Full_Adder FA_9919(s9919, c9919, in9919_1, in9919_2, s7451[0]);
    wire[0:0] s9920, in9920_1, in9920_2;
    wire c9920;
    assign in9920_1 = {s7455[0]};
    assign in9920_2 = {s7456[0]};
    Full_Adder FA_9920(s9920, c9920, in9920_1, in9920_2, s7454[0]);
    wire[0:0] s9921, in9921_1, in9921_2;
    wire c9921;
    assign in9921_1 = {s7458[0]};
    assign in9921_2 = {s7459[0]};
    Full_Adder FA_9921(s9921, c9921, in9921_1, in9921_2, s7457[0]);
    wire[0:0] s9922, in9922_1, in9922_2;
    wire c9922;
    assign in9922_1 = {c7441};
    assign in9922_2 = {c7442};
    Full_Adder FA_9922(s9922, c9922, in9922_1, in9922_2, s4799[0]);
    wire[0:0] s9923, in9923_1, in9923_2;
    wire c9923;
    assign in9923_1 = {c7444};
    assign in9923_2 = {c7445};
    Full_Adder FA_9923(s9923, c9923, in9923_1, in9923_2, c7443);
    wire[0:0] s9924, in9924_1, in9924_2;
    wire c9924;
    assign in9924_1 = {c7447};
    assign in9924_2 = {c7448};
    Full_Adder FA_9924(s9924, c9924, in9924_1, in9924_2, c7446);
    wire[0:0] s9925, in9925_1, in9925_2;
    wire c9925;
    assign in9925_1 = {c7450};
    assign in9925_2 = {c7451};
    Full_Adder FA_9925(s9925, c9925, in9925_1, in9925_2, c7449);
    wire[0:0] s9926, in9926_1, in9926_2;
    wire c9926;
    assign in9926_1 = {c7453};
    assign in9926_2 = {c7454};
    Full_Adder FA_9926(s9926, c9926, in9926_1, in9926_2, c7452);
    wire[0:0] s9927, in9927_1, in9927_2;
    wire c9927;
    assign in9927_1 = {c7456};
    assign in9927_2 = {c7457};
    Full_Adder FA_9927(s9927, c9927, in9927_1, in9927_2, c7455);
    wire[0:0] s9928, in9928_1, in9928_2;
    wire c9928;
    assign in9928_1 = {c7459};
    assign in9928_2 = {s7460[0]};
    Full_Adder FA_9928(s9928, c9928, in9928_1, in9928_2, c7458);
    wire[0:0] s9929, in9929_1, in9929_2;
    wire c9929;
    assign in9929_1 = {s7462[0]};
    assign in9929_2 = {s7463[0]};
    Full_Adder FA_9929(s9929, c9929, in9929_1, in9929_2, s7461[0]);
    wire[0:0] s9930, in9930_1, in9930_2;
    wire c9930;
    assign in9930_1 = {s7465[0]};
    assign in9930_2 = {s7466[0]};
    Full_Adder FA_9930(s9930, c9930, in9930_1, in9930_2, s7464[0]);
    wire[0:0] s9931, in9931_1, in9931_2;
    wire c9931;
    assign in9931_1 = {s7468[0]};
    assign in9931_2 = {s7469[0]};
    Full_Adder FA_9931(s9931, c9931, in9931_1, in9931_2, s7467[0]);
    wire[0:0] s9932, in9932_1, in9932_2;
    wire c9932;
    assign in9932_1 = {s7471[0]};
    assign in9932_2 = {s7472[0]};
    Full_Adder FA_9932(s9932, c9932, in9932_1, in9932_2, s7470[0]);
    wire[0:0] s9933, in9933_1, in9933_2;
    wire c9933;
    assign in9933_1 = {s7474[0]};
    assign in9933_2 = {s7475[0]};
    Full_Adder FA_9933(s9933, c9933, in9933_1, in9933_2, s7473[0]);
    wire[0:0] s9934, in9934_1, in9934_2;
    wire c9934;
    assign in9934_1 = {s7477[0]};
    assign in9934_2 = {s7478[0]};
    Full_Adder FA_9934(s9934, c9934, in9934_1, in9934_2, s7476[0]);
    wire[0:0] s9935, in9935_1, in9935_2;
    wire c9935;
    assign in9935_1 = {c7460};
    assign in9935_2 = {c7461};
    Full_Adder FA_9935(s9935, c9935, in9935_1, in9935_2, s4817[0]);
    wire[0:0] s9936, in9936_1, in9936_2;
    wire c9936;
    assign in9936_1 = {c7463};
    assign in9936_2 = {c7464};
    Full_Adder FA_9936(s9936, c9936, in9936_1, in9936_2, c7462);
    wire[0:0] s9937, in9937_1, in9937_2;
    wire c9937;
    assign in9937_1 = {c7466};
    assign in9937_2 = {c7467};
    Full_Adder FA_9937(s9937, c9937, in9937_1, in9937_2, c7465);
    wire[0:0] s9938, in9938_1, in9938_2;
    wire c9938;
    assign in9938_1 = {c7469};
    assign in9938_2 = {c7470};
    Full_Adder FA_9938(s9938, c9938, in9938_1, in9938_2, c7468);
    wire[0:0] s9939, in9939_1, in9939_2;
    wire c9939;
    assign in9939_1 = {c7472};
    assign in9939_2 = {c7473};
    Full_Adder FA_9939(s9939, c9939, in9939_1, in9939_2, c7471);
    wire[0:0] s9940, in9940_1, in9940_2;
    wire c9940;
    assign in9940_1 = {c7475};
    assign in9940_2 = {c7476};
    Full_Adder FA_9940(s9940, c9940, in9940_1, in9940_2, c7474);
    wire[0:0] s9941, in9941_1, in9941_2;
    wire c9941;
    assign in9941_1 = {c7478};
    assign in9941_2 = {s7479[0]};
    Full_Adder FA_9941(s9941, c9941, in9941_1, in9941_2, c7477);
    wire[0:0] s9942, in9942_1, in9942_2;
    wire c9942;
    assign in9942_1 = {s7481[0]};
    assign in9942_2 = {s7482[0]};
    Full_Adder FA_9942(s9942, c9942, in9942_1, in9942_2, s7480[0]);
    wire[0:0] s9943, in9943_1, in9943_2;
    wire c9943;
    assign in9943_1 = {s7484[0]};
    assign in9943_2 = {s7485[0]};
    Full_Adder FA_9943(s9943, c9943, in9943_1, in9943_2, s7483[0]);
    wire[0:0] s9944, in9944_1, in9944_2;
    wire c9944;
    assign in9944_1 = {s7487[0]};
    assign in9944_2 = {s7488[0]};
    Full_Adder FA_9944(s9944, c9944, in9944_1, in9944_2, s7486[0]);
    wire[0:0] s9945, in9945_1, in9945_2;
    wire c9945;
    assign in9945_1 = {s7490[0]};
    assign in9945_2 = {s7491[0]};
    Full_Adder FA_9945(s9945, c9945, in9945_1, in9945_2, s7489[0]);
    wire[0:0] s9946, in9946_1, in9946_2;
    wire c9946;
    assign in9946_1 = {s7493[0]};
    assign in9946_2 = {s7494[0]};
    Full_Adder FA_9946(s9946, c9946, in9946_1, in9946_2, s7492[0]);
    wire[0:0] s9947, in9947_1, in9947_2;
    wire c9947;
    assign in9947_1 = {s7496[0]};
    assign in9947_2 = {s7497[0]};
    Full_Adder FA_9947(s9947, c9947, in9947_1, in9947_2, s7495[0]);
    wire[0:0] s9948, in9948_1, in9948_2;
    wire c9948;
    assign in9948_1 = {c7479};
    assign in9948_2 = {c7480};
    Full_Adder FA_9948(s9948, c9948, in9948_1, in9948_2, s4834[0]);
    wire[0:0] s9949, in9949_1, in9949_2;
    wire c9949;
    assign in9949_1 = {c7482};
    assign in9949_2 = {c7483};
    Full_Adder FA_9949(s9949, c9949, in9949_1, in9949_2, c7481);
    wire[0:0] s9950, in9950_1, in9950_2;
    wire c9950;
    assign in9950_1 = {c7485};
    assign in9950_2 = {c7486};
    Full_Adder FA_9950(s9950, c9950, in9950_1, in9950_2, c7484);
    wire[0:0] s9951, in9951_1, in9951_2;
    wire c9951;
    assign in9951_1 = {c7488};
    assign in9951_2 = {c7489};
    Full_Adder FA_9951(s9951, c9951, in9951_1, in9951_2, c7487);
    wire[0:0] s9952, in9952_1, in9952_2;
    wire c9952;
    assign in9952_1 = {c7491};
    assign in9952_2 = {c7492};
    Full_Adder FA_9952(s9952, c9952, in9952_1, in9952_2, c7490);
    wire[0:0] s9953, in9953_1, in9953_2;
    wire c9953;
    assign in9953_1 = {c7494};
    assign in9953_2 = {c7495};
    Full_Adder FA_9953(s9953, c9953, in9953_1, in9953_2, c7493);
    wire[0:0] s9954, in9954_1, in9954_2;
    wire c9954;
    assign in9954_1 = {c7497};
    assign in9954_2 = {s7498[0]};
    Full_Adder FA_9954(s9954, c9954, in9954_1, in9954_2, c7496);
    wire[0:0] s9955, in9955_1, in9955_2;
    wire c9955;
    assign in9955_1 = {s7500[0]};
    assign in9955_2 = {s7501[0]};
    Full_Adder FA_9955(s9955, c9955, in9955_1, in9955_2, s7499[0]);
    wire[0:0] s9956, in9956_1, in9956_2;
    wire c9956;
    assign in9956_1 = {s7503[0]};
    assign in9956_2 = {s7504[0]};
    Full_Adder FA_9956(s9956, c9956, in9956_1, in9956_2, s7502[0]);
    wire[0:0] s9957, in9957_1, in9957_2;
    wire c9957;
    assign in9957_1 = {s7506[0]};
    assign in9957_2 = {s7507[0]};
    Full_Adder FA_9957(s9957, c9957, in9957_1, in9957_2, s7505[0]);
    wire[0:0] s9958, in9958_1, in9958_2;
    wire c9958;
    assign in9958_1 = {s7509[0]};
    assign in9958_2 = {s7510[0]};
    Full_Adder FA_9958(s9958, c9958, in9958_1, in9958_2, s7508[0]);
    wire[0:0] s9959, in9959_1, in9959_2;
    wire c9959;
    assign in9959_1 = {s7512[0]};
    assign in9959_2 = {s7513[0]};
    Full_Adder FA_9959(s9959, c9959, in9959_1, in9959_2, s7511[0]);
    wire[0:0] s9960, in9960_1, in9960_2;
    wire c9960;
    assign in9960_1 = {s7515[0]};
    assign in9960_2 = {s7516[0]};
    Full_Adder FA_9960(s9960, c9960, in9960_1, in9960_2, s7514[0]);
    wire[0:0] s9961, in9961_1, in9961_2;
    wire c9961;
    assign in9961_1 = {c7498};
    assign in9961_2 = {c7499};
    Full_Adder FA_9961(s9961, c9961, in9961_1, in9961_2, s4850[0]);
    wire[0:0] s9962, in9962_1, in9962_2;
    wire c9962;
    assign in9962_1 = {c7501};
    assign in9962_2 = {c7502};
    Full_Adder FA_9962(s9962, c9962, in9962_1, in9962_2, c7500);
    wire[0:0] s9963, in9963_1, in9963_2;
    wire c9963;
    assign in9963_1 = {c7504};
    assign in9963_2 = {c7505};
    Full_Adder FA_9963(s9963, c9963, in9963_1, in9963_2, c7503);
    wire[0:0] s9964, in9964_1, in9964_2;
    wire c9964;
    assign in9964_1 = {c7507};
    assign in9964_2 = {c7508};
    Full_Adder FA_9964(s9964, c9964, in9964_1, in9964_2, c7506);
    wire[0:0] s9965, in9965_1, in9965_2;
    wire c9965;
    assign in9965_1 = {c7510};
    assign in9965_2 = {c7511};
    Full_Adder FA_9965(s9965, c9965, in9965_1, in9965_2, c7509);
    wire[0:0] s9966, in9966_1, in9966_2;
    wire c9966;
    assign in9966_1 = {c7513};
    assign in9966_2 = {c7514};
    Full_Adder FA_9966(s9966, c9966, in9966_1, in9966_2, c7512);
    wire[0:0] s9967, in9967_1, in9967_2;
    wire c9967;
    assign in9967_1 = {c7516};
    assign in9967_2 = {s7517[0]};
    Full_Adder FA_9967(s9967, c9967, in9967_1, in9967_2, c7515);
    wire[0:0] s9968, in9968_1, in9968_2;
    wire c9968;
    assign in9968_1 = {s7519[0]};
    assign in9968_2 = {s7520[0]};
    Full_Adder FA_9968(s9968, c9968, in9968_1, in9968_2, s7518[0]);
    wire[0:0] s9969, in9969_1, in9969_2;
    wire c9969;
    assign in9969_1 = {s7522[0]};
    assign in9969_2 = {s7523[0]};
    Full_Adder FA_9969(s9969, c9969, in9969_1, in9969_2, s7521[0]);
    wire[0:0] s9970, in9970_1, in9970_2;
    wire c9970;
    assign in9970_1 = {s7525[0]};
    assign in9970_2 = {s7526[0]};
    Full_Adder FA_9970(s9970, c9970, in9970_1, in9970_2, s7524[0]);
    wire[0:0] s9971, in9971_1, in9971_2;
    wire c9971;
    assign in9971_1 = {s7528[0]};
    assign in9971_2 = {s7529[0]};
    Full_Adder FA_9971(s9971, c9971, in9971_1, in9971_2, s7527[0]);
    wire[0:0] s9972, in9972_1, in9972_2;
    wire c9972;
    assign in9972_1 = {s7531[0]};
    assign in9972_2 = {s7532[0]};
    Full_Adder FA_9972(s9972, c9972, in9972_1, in9972_2, s7530[0]);
    wire[0:0] s9973, in9973_1, in9973_2;
    wire c9973;
    assign in9973_1 = {s7534[0]};
    assign in9973_2 = {s7535[0]};
    Full_Adder FA_9973(s9973, c9973, in9973_1, in9973_2, s7533[0]);
    wire[0:0] s9974, in9974_1, in9974_2;
    wire c9974;
    assign in9974_1 = {c7517};
    assign in9974_2 = {c7518};
    Full_Adder FA_9974(s9974, c9974, in9974_1, in9974_2, s4865[0]);
    wire[0:0] s9975, in9975_1, in9975_2;
    wire c9975;
    assign in9975_1 = {c7520};
    assign in9975_2 = {c7521};
    Full_Adder FA_9975(s9975, c9975, in9975_1, in9975_2, c7519);
    wire[0:0] s9976, in9976_1, in9976_2;
    wire c9976;
    assign in9976_1 = {c7523};
    assign in9976_2 = {c7524};
    Full_Adder FA_9976(s9976, c9976, in9976_1, in9976_2, c7522);
    wire[0:0] s9977, in9977_1, in9977_2;
    wire c9977;
    assign in9977_1 = {c7526};
    assign in9977_2 = {c7527};
    Full_Adder FA_9977(s9977, c9977, in9977_1, in9977_2, c7525);
    wire[0:0] s9978, in9978_1, in9978_2;
    wire c9978;
    assign in9978_1 = {c7529};
    assign in9978_2 = {c7530};
    Full_Adder FA_9978(s9978, c9978, in9978_1, in9978_2, c7528);
    wire[0:0] s9979, in9979_1, in9979_2;
    wire c9979;
    assign in9979_1 = {c7532};
    assign in9979_2 = {c7533};
    Full_Adder FA_9979(s9979, c9979, in9979_1, in9979_2, c7531);
    wire[0:0] s9980, in9980_1, in9980_2;
    wire c9980;
    assign in9980_1 = {c7535};
    assign in9980_2 = {s7536[0]};
    Full_Adder FA_9980(s9980, c9980, in9980_1, in9980_2, c7534);
    wire[0:0] s9981, in9981_1, in9981_2;
    wire c9981;
    assign in9981_1 = {s7538[0]};
    assign in9981_2 = {s7539[0]};
    Full_Adder FA_9981(s9981, c9981, in9981_1, in9981_2, s7537[0]);
    wire[0:0] s9982, in9982_1, in9982_2;
    wire c9982;
    assign in9982_1 = {s7541[0]};
    assign in9982_2 = {s7542[0]};
    Full_Adder FA_9982(s9982, c9982, in9982_1, in9982_2, s7540[0]);
    wire[0:0] s9983, in9983_1, in9983_2;
    wire c9983;
    assign in9983_1 = {s7544[0]};
    assign in9983_2 = {s7545[0]};
    Full_Adder FA_9983(s9983, c9983, in9983_1, in9983_2, s7543[0]);
    wire[0:0] s9984, in9984_1, in9984_2;
    wire c9984;
    assign in9984_1 = {s7547[0]};
    assign in9984_2 = {s7548[0]};
    Full_Adder FA_9984(s9984, c9984, in9984_1, in9984_2, s7546[0]);
    wire[0:0] s9985, in9985_1, in9985_2;
    wire c9985;
    assign in9985_1 = {s7550[0]};
    assign in9985_2 = {s7551[0]};
    Full_Adder FA_9985(s9985, c9985, in9985_1, in9985_2, s7549[0]);
    wire[0:0] s9986, in9986_1, in9986_2;
    wire c9986;
    assign in9986_1 = {s7553[0]};
    assign in9986_2 = {s7554[0]};
    Full_Adder FA_9986(s9986, c9986, in9986_1, in9986_2, s7552[0]);
    wire[0:0] s9987, in9987_1, in9987_2;
    wire c9987;
    assign in9987_1 = {c7536};
    assign in9987_2 = {c7537};
    Full_Adder FA_9987(s9987, c9987, in9987_1, in9987_2, s4879[0]);
    wire[0:0] s9988, in9988_1, in9988_2;
    wire c9988;
    assign in9988_1 = {c7539};
    assign in9988_2 = {c7540};
    Full_Adder FA_9988(s9988, c9988, in9988_1, in9988_2, c7538);
    wire[0:0] s9989, in9989_1, in9989_2;
    wire c9989;
    assign in9989_1 = {c7542};
    assign in9989_2 = {c7543};
    Full_Adder FA_9989(s9989, c9989, in9989_1, in9989_2, c7541);
    wire[0:0] s9990, in9990_1, in9990_2;
    wire c9990;
    assign in9990_1 = {c7545};
    assign in9990_2 = {c7546};
    Full_Adder FA_9990(s9990, c9990, in9990_1, in9990_2, c7544);
    wire[0:0] s9991, in9991_1, in9991_2;
    wire c9991;
    assign in9991_1 = {c7548};
    assign in9991_2 = {c7549};
    Full_Adder FA_9991(s9991, c9991, in9991_1, in9991_2, c7547);
    wire[0:0] s9992, in9992_1, in9992_2;
    wire c9992;
    assign in9992_1 = {c7551};
    assign in9992_2 = {c7552};
    Full_Adder FA_9992(s9992, c9992, in9992_1, in9992_2, c7550);
    wire[0:0] s9993, in9993_1, in9993_2;
    wire c9993;
    assign in9993_1 = {c7554};
    assign in9993_2 = {s7555[0]};
    Full_Adder FA_9993(s9993, c9993, in9993_1, in9993_2, c7553);
    wire[0:0] s9994, in9994_1, in9994_2;
    wire c9994;
    assign in9994_1 = {s7557[0]};
    assign in9994_2 = {s7558[0]};
    Full_Adder FA_9994(s9994, c9994, in9994_1, in9994_2, s7556[0]);
    wire[0:0] s9995, in9995_1, in9995_2;
    wire c9995;
    assign in9995_1 = {s7560[0]};
    assign in9995_2 = {s7561[0]};
    Full_Adder FA_9995(s9995, c9995, in9995_1, in9995_2, s7559[0]);
    wire[0:0] s9996, in9996_1, in9996_2;
    wire c9996;
    assign in9996_1 = {s7563[0]};
    assign in9996_2 = {s7564[0]};
    Full_Adder FA_9996(s9996, c9996, in9996_1, in9996_2, s7562[0]);
    wire[0:0] s9997, in9997_1, in9997_2;
    wire c9997;
    assign in9997_1 = {s7566[0]};
    assign in9997_2 = {s7567[0]};
    Full_Adder FA_9997(s9997, c9997, in9997_1, in9997_2, s7565[0]);
    wire[0:0] s9998, in9998_1, in9998_2;
    wire c9998;
    assign in9998_1 = {s7569[0]};
    assign in9998_2 = {s7570[0]};
    Full_Adder FA_9998(s9998, c9998, in9998_1, in9998_2, s7568[0]);
    wire[0:0] s9999, in9999_1, in9999_2;
    wire c9999;
    assign in9999_1 = {s7572[0]};
    assign in9999_2 = {s7573[0]};
    Full_Adder FA_9999(s9999, c9999, in9999_1, in9999_2, s7571[0]);
    wire[0:0] s10000, in10000_1, in10000_2;
    wire c10000;
    assign in10000_1 = {c7555};
    assign in10000_2 = {c7556};
    Full_Adder FA_10000(s10000, c10000, in10000_1, in10000_2, s4892[0]);
    wire[0:0] s10001, in10001_1, in10001_2;
    wire c10001;
    assign in10001_1 = {c7558};
    assign in10001_2 = {c7559};
    Full_Adder FA_10001(s10001, c10001, in10001_1, in10001_2, c7557);
    wire[0:0] s10002, in10002_1, in10002_2;
    wire c10002;
    assign in10002_1 = {c7561};
    assign in10002_2 = {c7562};
    Full_Adder FA_10002(s10002, c10002, in10002_1, in10002_2, c7560);
    wire[0:0] s10003, in10003_1, in10003_2;
    wire c10003;
    assign in10003_1 = {c7564};
    assign in10003_2 = {c7565};
    Full_Adder FA_10003(s10003, c10003, in10003_1, in10003_2, c7563);
    wire[0:0] s10004, in10004_1, in10004_2;
    wire c10004;
    assign in10004_1 = {c7567};
    assign in10004_2 = {c7568};
    Full_Adder FA_10004(s10004, c10004, in10004_1, in10004_2, c7566);
    wire[0:0] s10005, in10005_1, in10005_2;
    wire c10005;
    assign in10005_1 = {c7570};
    assign in10005_2 = {c7571};
    Full_Adder FA_10005(s10005, c10005, in10005_1, in10005_2, c7569);
    wire[0:0] s10006, in10006_1, in10006_2;
    wire c10006;
    assign in10006_1 = {c7573};
    assign in10006_2 = {s7574[0]};
    Full_Adder FA_10006(s10006, c10006, in10006_1, in10006_2, c7572);
    wire[0:0] s10007, in10007_1, in10007_2;
    wire c10007;
    assign in10007_1 = {s7576[0]};
    assign in10007_2 = {s7577[0]};
    Full_Adder FA_10007(s10007, c10007, in10007_1, in10007_2, s7575[0]);
    wire[0:0] s10008, in10008_1, in10008_2;
    wire c10008;
    assign in10008_1 = {s7579[0]};
    assign in10008_2 = {s7580[0]};
    Full_Adder FA_10008(s10008, c10008, in10008_1, in10008_2, s7578[0]);
    wire[0:0] s10009, in10009_1, in10009_2;
    wire c10009;
    assign in10009_1 = {s7582[0]};
    assign in10009_2 = {s7583[0]};
    Full_Adder FA_10009(s10009, c10009, in10009_1, in10009_2, s7581[0]);
    wire[0:0] s10010, in10010_1, in10010_2;
    wire c10010;
    assign in10010_1 = {s7585[0]};
    assign in10010_2 = {s7586[0]};
    Full_Adder FA_10010(s10010, c10010, in10010_1, in10010_2, s7584[0]);
    wire[0:0] s10011, in10011_1, in10011_2;
    wire c10011;
    assign in10011_1 = {s7588[0]};
    assign in10011_2 = {s7589[0]};
    Full_Adder FA_10011(s10011, c10011, in10011_1, in10011_2, s7587[0]);
    wire[0:0] s10012, in10012_1, in10012_2;
    wire c10012;
    assign in10012_1 = {s7591[0]};
    assign in10012_2 = {s7592[0]};
    Full_Adder FA_10012(s10012, c10012, in10012_1, in10012_2, s7590[0]);
    wire[0:0] s10013, in10013_1, in10013_2;
    wire c10013;
    assign in10013_1 = {c7574};
    assign in10013_2 = {c7575};
    Full_Adder FA_10013(s10013, c10013, in10013_1, in10013_2, s4904[0]);
    wire[0:0] s10014, in10014_1, in10014_2;
    wire c10014;
    assign in10014_1 = {c7577};
    assign in10014_2 = {c7578};
    Full_Adder FA_10014(s10014, c10014, in10014_1, in10014_2, c7576);
    wire[0:0] s10015, in10015_1, in10015_2;
    wire c10015;
    assign in10015_1 = {c7580};
    assign in10015_2 = {c7581};
    Full_Adder FA_10015(s10015, c10015, in10015_1, in10015_2, c7579);
    wire[0:0] s10016, in10016_1, in10016_2;
    wire c10016;
    assign in10016_1 = {c7583};
    assign in10016_2 = {c7584};
    Full_Adder FA_10016(s10016, c10016, in10016_1, in10016_2, c7582);
    wire[0:0] s10017, in10017_1, in10017_2;
    wire c10017;
    assign in10017_1 = {c7586};
    assign in10017_2 = {c7587};
    Full_Adder FA_10017(s10017, c10017, in10017_1, in10017_2, c7585);
    wire[0:0] s10018, in10018_1, in10018_2;
    wire c10018;
    assign in10018_1 = {c7589};
    assign in10018_2 = {c7590};
    Full_Adder FA_10018(s10018, c10018, in10018_1, in10018_2, c7588);
    wire[0:0] s10019, in10019_1, in10019_2;
    wire c10019;
    assign in10019_1 = {c7592};
    assign in10019_2 = {s7593[0]};
    Full_Adder FA_10019(s10019, c10019, in10019_1, in10019_2, c7591);
    wire[0:0] s10020, in10020_1, in10020_2;
    wire c10020;
    assign in10020_1 = {s7595[0]};
    assign in10020_2 = {s7596[0]};
    Full_Adder FA_10020(s10020, c10020, in10020_1, in10020_2, s7594[0]);
    wire[0:0] s10021, in10021_1, in10021_2;
    wire c10021;
    assign in10021_1 = {s7598[0]};
    assign in10021_2 = {s7599[0]};
    Full_Adder FA_10021(s10021, c10021, in10021_1, in10021_2, s7597[0]);
    wire[0:0] s10022, in10022_1, in10022_2;
    wire c10022;
    assign in10022_1 = {s7601[0]};
    assign in10022_2 = {s7602[0]};
    Full_Adder FA_10022(s10022, c10022, in10022_1, in10022_2, s7600[0]);
    wire[0:0] s10023, in10023_1, in10023_2;
    wire c10023;
    assign in10023_1 = {s7604[0]};
    assign in10023_2 = {s7605[0]};
    Full_Adder FA_10023(s10023, c10023, in10023_1, in10023_2, s7603[0]);
    wire[0:0] s10024, in10024_1, in10024_2;
    wire c10024;
    assign in10024_1 = {s7607[0]};
    assign in10024_2 = {s7608[0]};
    Full_Adder FA_10024(s10024, c10024, in10024_1, in10024_2, s7606[0]);
    wire[0:0] s10025, in10025_1, in10025_2;
    wire c10025;
    assign in10025_1 = {s7610[0]};
    assign in10025_2 = {s7611[0]};
    Full_Adder FA_10025(s10025, c10025, in10025_1, in10025_2, s7609[0]);
    wire[0:0] s10026, in10026_1, in10026_2;
    wire c10026;
    assign in10026_1 = {c7593};
    assign in10026_2 = {c7594};
    Full_Adder FA_10026(s10026, c10026, in10026_1, in10026_2, s4915[0]);
    wire[0:0] s10027, in10027_1, in10027_2;
    wire c10027;
    assign in10027_1 = {c7596};
    assign in10027_2 = {c7597};
    Full_Adder FA_10027(s10027, c10027, in10027_1, in10027_2, c7595);
    wire[0:0] s10028, in10028_1, in10028_2;
    wire c10028;
    assign in10028_1 = {c7599};
    assign in10028_2 = {c7600};
    Full_Adder FA_10028(s10028, c10028, in10028_1, in10028_2, c7598);
    wire[0:0] s10029, in10029_1, in10029_2;
    wire c10029;
    assign in10029_1 = {c7602};
    assign in10029_2 = {c7603};
    Full_Adder FA_10029(s10029, c10029, in10029_1, in10029_2, c7601);
    wire[0:0] s10030, in10030_1, in10030_2;
    wire c10030;
    assign in10030_1 = {c7605};
    assign in10030_2 = {c7606};
    Full_Adder FA_10030(s10030, c10030, in10030_1, in10030_2, c7604);
    wire[0:0] s10031, in10031_1, in10031_2;
    wire c10031;
    assign in10031_1 = {c7608};
    assign in10031_2 = {c7609};
    Full_Adder FA_10031(s10031, c10031, in10031_1, in10031_2, c7607);
    wire[0:0] s10032, in10032_1, in10032_2;
    wire c10032;
    assign in10032_1 = {c7611};
    assign in10032_2 = {s7612[0]};
    Full_Adder FA_10032(s10032, c10032, in10032_1, in10032_2, c7610);
    wire[0:0] s10033, in10033_1, in10033_2;
    wire c10033;
    assign in10033_1 = {s7614[0]};
    assign in10033_2 = {s7615[0]};
    Full_Adder FA_10033(s10033, c10033, in10033_1, in10033_2, s7613[0]);
    wire[0:0] s10034, in10034_1, in10034_2;
    wire c10034;
    assign in10034_1 = {s7617[0]};
    assign in10034_2 = {s7618[0]};
    Full_Adder FA_10034(s10034, c10034, in10034_1, in10034_2, s7616[0]);
    wire[0:0] s10035, in10035_1, in10035_2;
    wire c10035;
    assign in10035_1 = {s7620[0]};
    assign in10035_2 = {s7621[0]};
    Full_Adder FA_10035(s10035, c10035, in10035_1, in10035_2, s7619[0]);
    wire[0:0] s10036, in10036_1, in10036_2;
    wire c10036;
    assign in10036_1 = {s7623[0]};
    assign in10036_2 = {s7624[0]};
    Full_Adder FA_10036(s10036, c10036, in10036_1, in10036_2, s7622[0]);
    wire[0:0] s10037, in10037_1, in10037_2;
    wire c10037;
    assign in10037_1 = {s7626[0]};
    assign in10037_2 = {s7627[0]};
    Full_Adder FA_10037(s10037, c10037, in10037_1, in10037_2, s7625[0]);
    wire[0:0] s10038, in10038_1, in10038_2;
    wire c10038;
    assign in10038_1 = {s7629[0]};
    assign in10038_2 = {s7630[0]};
    Full_Adder FA_10038(s10038, c10038, in10038_1, in10038_2, s7628[0]);
    wire[0:0] s10039, in10039_1, in10039_2;
    wire c10039;
    assign in10039_1 = {c7612};
    assign in10039_2 = {c7613};
    Full_Adder FA_10039(s10039, c10039, in10039_1, in10039_2, s4925[0]);
    wire[0:0] s10040, in10040_1, in10040_2;
    wire c10040;
    assign in10040_1 = {c7615};
    assign in10040_2 = {c7616};
    Full_Adder FA_10040(s10040, c10040, in10040_1, in10040_2, c7614);
    wire[0:0] s10041, in10041_1, in10041_2;
    wire c10041;
    assign in10041_1 = {c7618};
    assign in10041_2 = {c7619};
    Full_Adder FA_10041(s10041, c10041, in10041_1, in10041_2, c7617);
    wire[0:0] s10042, in10042_1, in10042_2;
    wire c10042;
    assign in10042_1 = {c7621};
    assign in10042_2 = {c7622};
    Full_Adder FA_10042(s10042, c10042, in10042_1, in10042_2, c7620);
    wire[0:0] s10043, in10043_1, in10043_2;
    wire c10043;
    assign in10043_1 = {c7624};
    assign in10043_2 = {c7625};
    Full_Adder FA_10043(s10043, c10043, in10043_1, in10043_2, c7623);
    wire[0:0] s10044, in10044_1, in10044_2;
    wire c10044;
    assign in10044_1 = {c7627};
    assign in10044_2 = {c7628};
    Full_Adder FA_10044(s10044, c10044, in10044_1, in10044_2, c7626);
    wire[0:0] s10045, in10045_1, in10045_2;
    wire c10045;
    assign in10045_1 = {c7630};
    assign in10045_2 = {s7631[0]};
    Full_Adder FA_10045(s10045, c10045, in10045_1, in10045_2, c7629);
    wire[0:0] s10046, in10046_1, in10046_2;
    wire c10046;
    assign in10046_1 = {s7633[0]};
    assign in10046_2 = {s7634[0]};
    Full_Adder FA_10046(s10046, c10046, in10046_1, in10046_2, s7632[0]);
    wire[0:0] s10047, in10047_1, in10047_2;
    wire c10047;
    assign in10047_1 = {s7636[0]};
    assign in10047_2 = {s7637[0]};
    Full_Adder FA_10047(s10047, c10047, in10047_1, in10047_2, s7635[0]);
    wire[0:0] s10048, in10048_1, in10048_2;
    wire c10048;
    assign in10048_1 = {s7639[0]};
    assign in10048_2 = {s7640[0]};
    Full_Adder FA_10048(s10048, c10048, in10048_1, in10048_2, s7638[0]);
    wire[0:0] s10049, in10049_1, in10049_2;
    wire c10049;
    assign in10049_1 = {s7642[0]};
    assign in10049_2 = {s7643[0]};
    Full_Adder FA_10049(s10049, c10049, in10049_1, in10049_2, s7641[0]);
    wire[0:0] s10050, in10050_1, in10050_2;
    wire c10050;
    assign in10050_1 = {s7645[0]};
    assign in10050_2 = {s7646[0]};
    Full_Adder FA_10050(s10050, c10050, in10050_1, in10050_2, s7644[0]);
    wire[0:0] s10051, in10051_1, in10051_2;
    wire c10051;
    assign in10051_1 = {s7648[0]};
    assign in10051_2 = {s7649[0]};
    Full_Adder FA_10051(s10051, c10051, in10051_1, in10051_2, s7647[0]);
    wire[0:0] s10052, in10052_1, in10052_2;
    wire c10052;
    assign in10052_1 = {c7631};
    assign in10052_2 = {c7632};
    Full_Adder FA_10052(s10052, c10052, in10052_1, in10052_2, s4934[0]);
    wire[0:0] s10053, in10053_1, in10053_2;
    wire c10053;
    assign in10053_1 = {c7634};
    assign in10053_2 = {c7635};
    Full_Adder FA_10053(s10053, c10053, in10053_1, in10053_2, c7633);
    wire[0:0] s10054, in10054_1, in10054_2;
    wire c10054;
    assign in10054_1 = {c7637};
    assign in10054_2 = {c7638};
    Full_Adder FA_10054(s10054, c10054, in10054_1, in10054_2, c7636);
    wire[0:0] s10055, in10055_1, in10055_2;
    wire c10055;
    assign in10055_1 = {c7640};
    assign in10055_2 = {c7641};
    Full_Adder FA_10055(s10055, c10055, in10055_1, in10055_2, c7639);
    wire[0:0] s10056, in10056_1, in10056_2;
    wire c10056;
    assign in10056_1 = {c7643};
    assign in10056_2 = {c7644};
    Full_Adder FA_10056(s10056, c10056, in10056_1, in10056_2, c7642);
    wire[0:0] s10057, in10057_1, in10057_2;
    wire c10057;
    assign in10057_1 = {c7646};
    assign in10057_2 = {c7647};
    Full_Adder FA_10057(s10057, c10057, in10057_1, in10057_2, c7645);
    wire[0:0] s10058, in10058_1, in10058_2;
    wire c10058;
    assign in10058_1 = {c7649};
    assign in10058_2 = {s7650[0]};
    Full_Adder FA_10058(s10058, c10058, in10058_1, in10058_2, c7648);
    wire[0:0] s10059, in10059_1, in10059_2;
    wire c10059;
    assign in10059_1 = {s7652[0]};
    assign in10059_2 = {s7653[0]};
    Full_Adder FA_10059(s10059, c10059, in10059_1, in10059_2, s7651[0]);
    wire[0:0] s10060, in10060_1, in10060_2;
    wire c10060;
    assign in10060_1 = {s7655[0]};
    assign in10060_2 = {s7656[0]};
    Full_Adder FA_10060(s10060, c10060, in10060_1, in10060_2, s7654[0]);
    wire[0:0] s10061, in10061_1, in10061_2;
    wire c10061;
    assign in10061_1 = {s7658[0]};
    assign in10061_2 = {s7659[0]};
    Full_Adder FA_10061(s10061, c10061, in10061_1, in10061_2, s7657[0]);
    wire[0:0] s10062, in10062_1, in10062_2;
    wire c10062;
    assign in10062_1 = {s7661[0]};
    assign in10062_2 = {s7662[0]};
    Full_Adder FA_10062(s10062, c10062, in10062_1, in10062_2, s7660[0]);
    wire[0:0] s10063, in10063_1, in10063_2;
    wire c10063;
    assign in10063_1 = {s7664[0]};
    assign in10063_2 = {s7665[0]};
    Full_Adder FA_10063(s10063, c10063, in10063_1, in10063_2, s7663[0]);
    wire[0:0] s10064, in10064_1, in10064_2;
    wire c10064;
    assign in10064_1 = {s7667[0]};
    assign in10064_2 = {s7668[0]};
    Full_Adder FA_10064(s10064, c10064, in10064_1, in10064_2, s7666[0]);
    wire[0:0] s10065, in10065_1, in10065_2;
    wire c10065;
    assign in10065_1 = {c7650};
    assign in10065_2 = {c7651};
    Full_Adder FA_10065(s10065, c10065, in10065_1, in10065_2, s4942[0]);
    wire[0:0] s10066, in10066_1, in10066_2;
    wire c10066;
    assign in10066_1 = {c7653};
    assign in10066_2 = {c7654};
    Full_Adder FA_10066(s10066, c10066, in10066_1, in10066_2, c7652);
    wire[0:0] s10067, in10067_1, in10067_2;
    wire c10067;
    assign in10067_1 = {c7656};
    assign in10067_2 = {c7657};
    Full_Adder FA_10067(s10067, c10067, in10067_1, in10067_2, c7655);
    wire[0:0] s10068, in10068_1, in10068_2;
    wire c10068;
    assign in10068_1 = {c7659};
    assign in10068_2 = {c7660};
    Full_Adder FA_10068(s10068, c10068, in10068_1, in10068_2, c7658);
    wire[0:0] s10069, in10069_1, in10069_2;
    wire c10069;
    assign in10069_1 = {c7662};
    assign in10069_2 = {c7663};
    Full_Adder FA_10069(s10069, c10069, in10069_1, in10069_2, c7661);
    wire[0:0] s10070, in10070_1, in10070_2;
    wire c10070;
    assign in10070_1 = {c7665};
    assign in10070_2 = {c7666};
    Full_Adder FA_10070(s10070, c10070, in10070_1, in10070_2, c7664);
    wire[0:0] s10071, in10071_1, in10071_2;
    wire c10071;
    assign in10071_1 = {c7668};
    assign in10071_2 = {s7669[0]};
    Full_Adder FA_10071(s10071, c10071, in10071_1, in10071_2, c7667);
    wire[0:0] s10072, in10072_1, in10072_2;
    wire c10072;
    assign in10072_1 = {s7671[0]};
    assign in10072_2 = {s7672[0]};
    Full_Adder FA_10072(s10072, c10072, in10072_1, in10072_2, s7670[0]);
    wire[0:0] s10073, in10073_1, in10073_2;
    wire c10073;
    assign in10073_1 = {s7674[0]};
    assign in10073_2 = {s7675[0]};
    Full_Adder FA_10073(s10073, c10073, in10073_1, in10073_2, s7673[0]);
    wire[0:0] s10074, in10074_1, in10074_2;
    wire c10074;
    assign in10074_1 = {s7677[0]};
    assign in10074_2 = {s7678[0]};
    Full_Adder FA_10074(s10074, c10074, in10074_1, in10074_2, s7676[0]);
    wire[0:0] s10075, in10075_1, in10075_2;
    wire c10075;
    assign in10075_1 = {s7680[0]};
    assign in10075_2 = {s7681[0]};
    Full_Adder FA_10075(s10075, c10075, in10075_1, in10075_2, s7679[0]);
    wire[0:0] s10076, in10076_1, in10076_2;
    wire c10076;
    assign in10076_1 = {s7683[0]};
    assign in10076_2 = {s7684[0]};
    Full_Adder FA_10076(s10076, c10076, in10076_1, in10076_2, s7682[0]);
    wire[0:0] s10077, in10077_1, in10077_2;
    wire c10077;
    assign in10077_1 = {s7686[0]};
    assign in10077_2 = {s7687[0]};
    Full_Adder FA_10077(s10077, c10077, in10077_1, in10077_2, s7685[0]);
    wire[0:0] s10078, in10078_1, in10078_2;
    wire c10078;
    assign in10078_1 = {c7669};
    assign in10078_2 = {c7670};
    Full_Adder FA_10078(s10078, c10078, in10078_1, in10078_2, s4949[0]);
    wire[0:0] s10079, in10079_1, in10079_2;
    wire c10079;
    assign in10079_1 = {c7672};
    assign in10079_2 = {c7673};
    Full_Adder FA_10079(s10079, c10079, in10079_1, in10079_2, c7671);
    wire[0:0] s10080, in10080_1, in10080_2;
    wire c10080;
    assign in10080_1 = {c7675};
    assign in10080_2 = {c7676};
    Full_Adder FA_10080(s10080, c10080, in10080_1, in10080_2, c7674);
    wire[0:0] s10081, in10081_1, in10081_2;
    wire c10081;
    assign in10081_1 = {c7678};
    assign in10081_2 = {c7679};
    Full_Adder FA_10081(s10081, c10081, in10081_1, in10081_2, c7677);
    wire[0:0] s10082, in10082_1, in10082_2;
    wire c10082;
    assign in10082_1 = {c7681};
    assign in10082_2 = {c7682};
    Full_Adder FA_10082(s10082, c10082, in10082_1, in10082_2, c7680);
    wire[0:0] s10083, in10083_1, in10083_2;
    wire c10083;
    assign in10083_1 = {c7684};
    assign in10083_2 = {c7685};
    Full_Adder FA_10083(s10083, c10083, in10083_1, in10083_2, c7683);
    wire[0:0] s10084, in10084_1, in10084_2;
    wire c10084;
    assign in10084_1 = {c7687};
    assign in10084_2 = {s7688[0]};
    Full_Adder FA_10084(s10084, c10084, in10084_1, in10084_2, c7686);
    wire[0:0] s10085, in10085_1, in10085_2;
    wire c10085;
    assign in10085_1 = {s7690[0]};
    assign in10085_2 = {s7691[0]};
    Full_Adder FA_10085(s10085, c10085, in10085_1, in10085_2, s7689[0]);
    wire[0:0] s10086, in10086_1, in10086_2;
    wire c10086;
    assign in10086_1 = {s7693[0]};
    assign in10086_2 = {s7694[0]};
    Full_Adder FA_10086(s10086, c10086, in10086_1, in10086_2, s7692[0]);
    wire[0:0] s10087, in10087_1, in10087_2;
    wire c10087;
    assign in10087_1 = {s7696[0]};
    assign in10087_2 = {s7697[0]};
    Full_Adder FA_10087(s10087, c10087, in10087_1, in10087_2, s7695[0]);
    wire[0:0] s10088, in10088_1, in10088_2;
    wire c10088;
    assign in10088_1 = {s7699[0]};
    assign in10088_2 = {s7700[0]};
    Full_Adder FA_10088(s10088, c10088, in10088_1, in10088_2, s7698[0]);
    wire[0:0] s10089, in10089_1, in10089_2;
    wire c10089;
    assign in10089_1 = {s7702[0]};
    assign in10089_2 = {s7703[0]};
    Full_Adder FA_10089(s10089, c10089, in10089_1, in10089_2, s7701[0]);
    wire[0:0] s10090, in10090_1, in10090_2;
    wire c10090;
    assign in10090_1 = {s7705[0]};
    assign in10090_2 = {s7706[0]};
    Full_Adder FA_10090(s10090, c10090, in10090_1, in10090_2, s7704[0]);
    wire[0:0] s10091, in10091_1, in10091_2;
    wire c10091;
    assign in10091_1 = {c7688};
    assign in10091_2 = {c7689};
    Full_Adder FA_10091(s10091, c10091, in10091_1, in10091_2, s4955[0]);
    wire[0:0] s10092, in10092_1, in10092_2;
    wire c10092;
    assign in10092_1 = {c7691};
    assign in10092_2 = {c7692};
    Full_Adder FA_10092(s10092, c10092, in10092_1, in10092_2, c7690);
    wire[0:0] s10093, in10093_1, in10093_2;
    wire c10093;
    assign in10093_1 = {c7694};
    assign in10093_2 = {c7695};
    Full_Adder FA_10093(s10093, c10093, in10093_1, in10093_2, c7693);
    wire[0:0] s10094, in10094_1, in10094_2;
    wire c10094;
    assign in10094_1 = {c7697};
    assign in10094_2 = {c7698};
    Full_Adder FA_10094(s10094, c10094, in10094_1, in10094_2, c7696);
    wire[0:0] s10095, in10095_1, in10095_2;
    wire c10095;
    assign in10095_1 = {c7700};
    assign in10095_2 = {c7701};
    Full_Adder FA_10095(s10095, c10095, in10095_1, in10095_2, c7699);
    wire[0:0] s10096, in10096_1, in10096_2;
    wire c10096;
    assign in10096_1 = {c7703};
    assign in10096_2 = {c7704};
    Full_Adder FA_10096(s10096, c10096, in10096_1, in10096_2, c7702);
    wire[0:0] s10097, in10097_1, in10097_2;
    wire c10097;
    assign in10097_1 = {c7706};
    assign in10097_2 = {s7707[0]};
    Full_Adder FA_10097(s10097, c10097, in10097_1, in10097_2, c7705);
    wire[0:0] s10098, in10098_1, in10098_2;
    wire c10098;
    assign in10098_1 = {s7709[0]};
    assign in10098_2 = {s7710[0]};
    Full_Adder FA_10098(s10098, c10098, in10098_1, in10098_2, s7708[0]);
    wire[0:0] s10099, in10099_1, in10099_2;
    wire c10099;
    assign in10099_1 = {s7712[0]};
    assign in10099_2 = {s7713[0]};
    Full_Adder FA_10099(s10099, c10099, in10099_1, in10099_2, s7711[0]);
    wire[0:0] s10100, in10100_1, in10100_2;
    wire c10100;
    assign in10100_1 = {s7715[0]};
    assign in10100_2 = {s7716[0]};
    Full_Adder FA_10100(s10100, c10100, in10100_1, in10100_2, s7714[0]);
    wire[0:0] s10101, in10101_1, in10101_2;
    wire c10101;
    assign in10101_1 = {s7718[0]};
    assign in10101_2 = {s7719[0]};
    Full_Adder FA_10101(s10101, c10101, in10101_1, in10101_2, s7717[0]);
    wire[0:0] s10102, in10102_1, in10102_2;
    wire c10102;
    assign in10102_1 = {s7721[0]};
    assign in10102_2 = {s7722[0]};
    Full_Adder FA_10102(s10102, c10102, in10102_1, in10102_2, s7720[0]);
    wire[0:0] s10103, in10103_1, in10103_2;
    wire c10103;
    assign in10103_1 = {s7724[0]};
    assign in10103_2 = {s7725[0]};
    Full_Adder FA_10103(s10103, c10103, in10103_1, in10103_2, s7723[0]);
    wire[0:0] s10104, in10104_1, in10104_2;
    wire c10104;
    assign in10104_1 = {c7707};
    assign in10104_2 = {c7708};
    Full_Adder FA_10104(s10104, c10104, in10104_1, in10104_2, s4960[0]);
    wire[0:0] s10105, in10105_1, in10105_2;
    wire c10105;
    assign in10105_1 = {c7710};
    assign in10105_2 = {c7711};
    Full_Adder FA_10105(s10105, c10105, in10105_1, in10105_2, c7709);
    wire[0:0] s10106, in10106_1, in10106_2;
    wire c10106;
    assign in10106_1 = {c7713};
    assign in10106_2 = {c7714};
    Full_Adder FA_10106(s10106, c10106, in10106_1, in10106_2, c7712);
    wire[0:0] s10107, in10107_1, in10107_2;
    wire c10107;
    assign in10107_1 = {c7716};
    assign in10107_2 = {c7717};
    Full_Adder FA_10107(s10107, c10107, in10107_1, in10107_2, c7715);
    wire[0:0] s10108, in10108_1, in10108_2;
    wire c10108;
    assign in10108_1 = {c7719};
    assign in10108_2 = {c7720};
    Full_Adder FA_10108(s10108, c10108, in10108_1, in10108_2, c7718);
    wire[0:0] s10109, in10109_1, in10109_2;
    wire c10109;
    assign in10109_1 = {c7722};
    assign in10109_2 = {c7723};
    Full_Adder FA_10109(s10109, c10109, in10109_1, in10109_2, c7721);
    wire[0:0] s10110, in10110_1, in10110_2;
    wire c10110;
    assign in10110_1 = {c7725};
    assign in10110_2 = {s7726[0]};
    Full_Adder FA_10110(s10110, c10110, in10110_1, in10110_2, c7724);
    wire[0:0] s10111, in10111_1, in10111_2;
    wire c10111;
    assign in10111_1 = {s7728[0]};
    assign in10111_2 = {s7729[0]};
    Full_Adder FA_10111(s10111, c10111, in10111_1, in10111_2, s7727[0]);
    wire[0:0] s10112, in10112_1, in10112_2;
    wire c10112;
    assign in10112_1 = {s7731[0]};
    assign in10112_2 = {s7732[0]};
    Full_Adder FA_10112(s10112, c10112, in10112_1, in10112_2, s7730[0]);
    wire[0:0] s10113, in10113_1, in10113_2;
    wire c10113;
    assign in10113_1 = {s7734[0]};
    assign in10113_2 = {s7735[0]};
    Full_Adder FA_10113(s10113, c10113, in10113_1, in10113_2, s7733[0]);
    wire[0:0] s10114, in10114_1, in10114_2;
    wire c10114;
    assign in10114_1 = {s7737[0]};
    assign in10114_2 = {s7738[0]};
    Full_Adder FA_10114(s10114, c10114, in10114_1, in10114_2, s7736[0]);
    wire[0:0] s10115, in10115_1, in10115_2;
    wire c10115;
    assign in10115_1 = {s7740[0]};
    assign in10115_2 = {s7741[0]};
    Full_Adder FA_10115(s10115, c10115, in10115_1, in10115_2, s7739[0]);
    wire[0:0] s10116, in10116_1, in10116_2;
    wire c10116;
    assign in10116_1 = {s7743[0]};
    assign in10116_2 = {s7744[0]};
    Full_Adder FA_10116(s10116, c10116, in10116_1, in10116_2, s7742[0]);
    wire[0:0] s10117, in10117_1, in10117_2;
    wire c10117;
    assign in10117_1 = {c7726};
    assign in10117_2 = {c7727};
    Full_Adder FA_10117(s10117, c10117, in10117_1, in10117_2, s4964[0]);
    wire[0:0] s10118, in10118_1, in10118_2;
    wire c10118;
    assign in10118_1 = {c7729};
    assign in10118_2 = {c7730};
    Full_Adder FA_10118(s10118, c10118, in10118_1, in10118_2, c7728);
    wire[0:0] s10119, in10119_1, in10119_2;
    wire c10119;
    assign in10119_1 = {c7732};
    assign in10119_2 = {c7733};
    Full_Adder FA_10119(s10119, c10119, in10119_1, in10119_2, c7731);
    wire[0:0] s10120, in10120_1, in10120_2;
    wire c10120;
    assign in10120_1 = {c7735};
    assign in10120_2 = {c7736};
    Full_Adder FA_10120(s10120, c10120, in10120_1, in10120_2, c7734);
    wire[0:0] s10121, in10121_1, in10121_2;
    wire c10121;
    assign in10121_1 = {c7738};
    assign in10121_2 = {c7739};
    Full_Adder FA_10121(s10121, c10121, in10121_1, in10121_2, c7737);
    wire[0:0] s10122, in10122_1, in10122_2;
    wire c10122;
    assign in10122_1 = {c7741};
    assign in10122_2 = {c7742};
    Full_Adder FA_10122(s10122, c10122, in10122_1, in10122_2, c7740);
    wire[0:0] s10123, in10123_1, in10123_2;
    wire c10123;
    assign in10123_1 = {c7744};
    assign in10123_2 = {s7745[0]};
    Full_Adder FA_10123(s10123, c10123, in10123_1, in10123_2, c7743);
    wire[0:0] s10124, in10124_1, in10124_2;
    wire c10124;
    assign in10124_1 = {s7747[0]};
    assign in10124_2 = {s7748[0]};
    Full_Adder FA_10124(s10124, c10124, in10124_1, in10124_2, s7746[0]);
    wire[0:0] s10125, in10125_1, in10125_2;
    wire c10125;
    assign in10125_1 = {s7750[0]};
    assign in10125_2 = {s7751[0]};
    Full_Adder FA_10125(s10125, c10125, in10125_1, in10125_2, s7749[0]);
    wire[0:0] s10126, in10126_1, in10126_2;
    wire c10126;
    assign in10126_1 = {s7753[0]};
    assign in10126_2 = {s7754[0]};
    Full_Adder FA_10126(s10126, c10126, in10126_1, in10126_2, s7752[0]);
    wire[0:0] s10127, in10127_1, in10127_2;
    wire c10127;
    assign in10127_1 = {s7756[0]};
    assign in10127_2 = {s7757[0]};
    Full_Adder FA_10127(s10127, c10127, in10127_1, in10127_2, s7755[0]);
    wire[0:0] s10128, in10128_1, in10128_2;
    wire c10128;
    assign in10128_1 = {s7759[0]};
    assign in10128_2 = {s7760[0]};
    Full_Adder FA_10128(s10128, c10128, in10128_1, in10128_2, s7758[0]);
    wire[0:0] s10129, in10129_1, in10129_2;
    wire c10129;
    assign in10129_1 = {s7762[0]};
    assign in10129_2 = {s7763[0]};
    Full_Adder FA_10129(s10129, c10129, in10129_1, in10129_2, s7761[0]);
    wire[0:0] s10130, in10130_1, in10130_2;
    wire c10130;
    assign in10130_1 = {c7745};
    assign in10130_2 = {c7746};
    Full_Adder FA_10130(s10130, c10130, in10130_1, in10130_2, s4967[0]);
    wire[0:0] s10131, in10131_1, in10131_2;
    wire c10131;
    assign in10131_1 = {c7748};
    assign in10131_2 = {c7749};
    Full_Adder FA_10131(s10131, c10131, in10131_1, in10131_2, c7747);
    wire[0:0] s10132, in10132_1, in10132_2;
    wire c10132;
    assign in10132_1 = {c7751};
    assign in10132_2 = {c7752};
    Full_Adder FA_10132(s10132, c10132, in10132_1, in10132_2, c7750);
    wire[0:0] s10133, in10133_1, in10133_2;
    wire c10133;
    assign in10133_1 = {c7754};
    assign in10133_2 = {c7755};
    Full_Adder FA_10133(s10133, c10133, in10133_1, in10133_2, c7753);
    wire[0:0] s10134, in10134_1, in10134_2;
    wire c10134;
    assign in10134_1 = {c7757};
    assign in10134_2 = {c7758};
    Full_Adder FA_10134(s10134, c10134, in10134_1, in10134_2, c7756);
    wire[0:0] s10135, in10135_1, in10135_2;
    wire c10135;
    assign in10135_1 = {c7760};
    assign in10135_2 = {c7761};
    Full_Adder FA_10135(s10135, c10135, in10135_1, in10135_2, c7759);
    wire[0:0] s10136, in10136_1, in10136_2;
    wire c10136;
    assign in10136_1 = {c7763};
    assign in10136_2 = {s7764[0]};
    Full_Adder FA_10136(s10136, c10136, in10136_1, in10136_2, c7762);
    wire[0:0] s10137, in10137_1, in10137_2;
    wire c10137;
    assign in10137_1 = {s7766[0]};
    assign in10137_2 = {s7767[0]};
    Full_Adder FA_10137(s10137, c10137, in10137_1, in10137_2, s7765[0]);
    wire[0:0] s10138, in10138_1, in10138_2;
    wire c10138;
    assign in10138_1 = {s7769[0]};
    assign in10138_2 = {s7770[0]};
    Full_Adder FA_10138(s10138, c10138, in10138_1, in10138_2, s7768[0]);
    wire[0:0] s10139, in10139_1, in10139_2;
    wire c10139;
    assign in10139_1 = {s7772[0]};
    assign in10139_2 = {s7773[0]};
    Full_Adder FA_10139(s10139, c10139, in10139_1, in10139_2, s7771[0]);
    wire[0:0] s10140, in10140_1, in10140_2;
    wire c10140;
    assign in10140_1 = {s7775[0]};
    assign in10140_2 = {s7776[0]};
    Full_Adder FA_10140(s10140, c10140, in10140_1, in10140_2, s7774[0]);
    wire[0:0] s10141, in10141_1, in10141_2;
    wire c10141;
    assign in10141_1 = {s7778[0]};
    assign in10141_2 = {s7779[0]};
    Full_Adder FA_10141(s10141, c10141, in10141_1, in10141_2, s7777[0]);
    wire[0:0] s10142, in10142_1, in10142_2;
    wire c10142;
    assign in10142_1 = {s7781[0]};
    assign in10142_2 = {s7782[0]};
    Full_Adder FA_10142(s10142, c10142, in10142_1, in10142_2, s7780[0]);
    wire[0:0] s10143, in10143_1, in10143_2;
    wire c10143;
    assign in10143_1 = {c7764};
    assign in10143_2 = {c7765};
    Full_Adder FA_10143(s10143, c10143, in10143_1, in10143_2, s4969[0]);
    wire[0:0] s10144, in10144_1, in10144_2;
    wire c10144;
    assign in10144_1 = {c7767};
    assign in10144_2 = {c7768};
    Full_Adder FA_10144(s10144, c10144, in10144_1, in10144_2, c7766);
    wire[0:0] s10145, in10145_1, in10145_2;
    wire c10145;
    assign in10145_1 = {c7770};
    assign in10145_2 = {c7771};
    Full_Adder FA_10145(s10145, c10145, in10145_1, in10145_2, c7769);
    wire[0:0] s10146, in10146_1, in10146_2;
    wire c10146;
    assign in10146_1 = {c7773};
    assign in10146_2 = {c7774};
    Full_Adder FA_10146(s10146, c10146, in10146_1, in10146_2, c7772);
    wire[0:0] s10147, in10147_1, in10147_2;
    wire c10147;
    assign in10147_1 = {c7776};
    assign in10147_2 = {c7777};
    Full_Adder FA_10147(s10147, c10147, in10147_1, in10147_2, c7775);
    wire[0:0] s10148, in10148_1, in10148_2;
    wire c10148;
    assign in10148_1 = {c7779};
    assign in10148_2 = {c7780};
    Full_Adder FA_10148(s10148, c10148, in10148_1, in10148_2, c7778);
    wire[0:0] s10149, in10149_1, in10149_2;
    wire c10149;
    assign in10149_1 = {c7782};
    assign in10149_2 = {s7783[0]};
    Full_Adder FA_10149(s10149, c10149, in10149_1, in10149_2, c7781);
    wire[0:0] s10150, in10150_1, in10150_2;
    wire c10150;
    assign in10150_1 = {s7785[0]};
    assign in10150_2 = {s7786[0]};
    Full_Adder FA_10150(s10150, c10150, in10150_1, in10150_2, s7784[0]);
    wire[0:0] s10151, in10151_1, in10151_2;
    wire c10151;
    assign in10151_1 = {s7788[0]};
    assign in10151_2 = {s7789[0]};
    Full_Adder FA_10151(s10151, c10151, in10151_1, in10151_2, s7787[0]);
    wire[0:0] s10152, in10152_1, in10152_2;
    wire c10152;
    assign in10152_1 = {s7791[0]};
    assign in10152_2 = {s7792[0]};
    Full_Adder FA_10152(s10152, c10152, in10152_1, in10152_2, s7790[0]);
    wire[0:0] s10153, in10153_1, in10153_2;
    wire c10153;
    assign in10153_1 = {s7794[0]};
    assign in10153_2 = {s7795[0]};
    Full_Adder FA_10153(s10153, c10153, in10153_1, in10153_2, s7793[0]);
    wire[0:0] s10154, in10154_1, in10154_2;
    wire c10154;
    assign in10154_1 = {s7797[0]};
    assign in10154_2 = {s7798[0]};
    Full_Adder FA_10154(s10154, c10154, in10154_1, in10154_2, s7796[0]);
    wire[0:0] s10155, in10155_1, in10155_2;
    wire c10155;
    assign in10155_1 = {s7800[0]};
    assign in10155_2 = {s7801[0]};
    Full_Adder FA_10155(s10155, c10155, in10155_1, in10155_2, s7799[0]);
    wire[0:0] s10156, in10156_1, in10156_2;
    wire c10156;
    assign in10156_1 = {c7783};
    assign in10156_2 = {c7784};
    Full_Adder FA_10156(s10156, c10156, in10156_1, in10156_2, s4970[0]);
    wire[0:0] s10157, in10157_1, in10157_2;
    wire c10157;
    assign in10157_1 = {c7786};
    assign in10157_2 = {c7787};
    Full_Adder FA_10157(s10157, c10157, in10157_1, in10157_2, c7785);
    wire[0:0] s10158, in10158_1, in10158_2;
    wire c10158;
    assign in10158_1 = {c7789};
    assign in10158_2 = {c7790};
    Full_Adder FA_10158(s10158, c10158, in10158_1, in10158_2, c7788);
    wire[0:0] s10159, in10159_1, in10159_2;
    wire c10159;
    assign in10159_1 = {c7792};
    assign in10159_2 = {c7793};
    Full_Adder FA_10159(s10159, c10159, in10159_1, in10159_2, c7791);
    wire[0:0] s10160, in10160_1, in10160_2;
    wire c10160;
    assign in10160_1 = {c7795};
    assign in10160_2 = {c7796};
    Full_Adder FA_10160(s10160, c10160, in10160_1, in10160_2, c7794);
    wire[0:0] s10161, in10161_1, in10161_2;
    wire c10161;
    assign in10161_1 = {c7798};
    assign in10161_2 = {c7799};
    Full_Adder FA_10161(s10161, c10161, in10161_1, in10161_2, c7797);
    wire[0:0] s10162, in10162_1, in10162_2;
    wire c10162;
    assign in10162_1 = {c7801};
    assign in10162_2 = {s7802[0]};
    Full_Adder FA_10162(s10162, c10162, in10162_1, in10162_2, c7800);
    wire[0:0] s10163, in10163_1, in10163_2;
    wire c10163;
    assign in10163_1 = {s7804[0]};
    assign in10163_2 = {s7805[0]};
    Full_Adder FA_10163(s10163, c10163, in10163_1, in10163_2, s7803[0]);
    wire[0:0] s10164, in10164_1, in10164_2;
    wire c10164;
    assign in10164_1 = {s7807[0]};
    assign in10164_2 = {s7808[0]};
    Full_Adder FA_10164(s10164, c10164, in10164_1, in10164_2, s7806[0]);
    wire[0:0] s10165, in10165_1, in10165_2;
    wire c10165;
    assign in10165_1 = {s7810[0]};
    assign in10165_2 = {s7811[0]};
    Full_Adder FA_10165(s10165, c10165, in10165_1, in10165_2, s7809[0]);
    wire[0:0] s10166, in10166_1, in10166_2;
    wire c10166;
    assign in10166_1 = {s7813[0]};
    assign in10166_2 = {s7814[0]};
    Full_Adder FA_10166(s10166, c10166, in10166_1, in10166_2, s7812[0]);
    wire[0:0] s10167, in10167_1, in10167_2;
    wire c10167;
    assign in10167_1 = {s7816[0]};
    assign in10167_2 = {s7817[0]};
    Full_Adder FA_10167(s10167, c10167, in10167_1, in10167_2, s7815[0]);
    wire[0:0] s10168, in10168_1, in10168_2;
    wire c10168;
    assign in10168_1 = {s7819[0]};
    assign in10168_2 = {s7820[0]};
    Full_Adder FA_10168(s10168, c10168, in10168_1, in10168_2, s7818[0]);
    wire[0:0] s10169, in10169_1, in10169_2;
    wire c10169;
    assign in10169_1 = {c7802};
    assign in10169_2 = {c7803};
    Full_Adder FA_10169(s10169, c10169, in10169_1, in10169_2, c4970);
    wire[0:0] s10170, in10170_1, in10170_2;
    wire c10170;
    assign in10170_1 = {c7805};
    assign in10170_2 = {c7806};
    Full_Adder FA_10170(s10170, c10170, in10170_1, in10170_2, c7804);
    wire[0:0] s10171, in10171_1, in10171_2;
    wire c10171;
    assign in10171_1 = {c7808};
    assign in10171_2 = {c7809};
    Full_Adder FA_10171(s10171, c10171, in10171_1, in10171_2, c7807);
    wire[0:0] s10172, in10172_1, in10172_2;
    wire c10172;
    assign in10172_1 = {c7811};
    assign in10172_2 = {c7812};
    Full_Adder FA_10172(s10172, c10172, in10172_1, in10172_2, c7810);
    wire[0:0] s10173, in10173_1, in10173_2;
    wire c10173;
    assign in10173_1 = {c7814};
    assign in10173_2 = {c7815};
    Full_Adder FA_10173(s10173, c10173, in10173_1, in10173_2, c7813);
    wire[0:0] s10174, in10174_1, in10174_2;
    wire c10174;
    assign in10174_1 = {c7817};
    assign in10174_2 = {c7818};
    Full_Adder FA_10174(s10174, c10174, in10174_1, in10174_2, c7816);
    wire[0:0] s10175, in10175_1, in10175_2;
    wire c10175;
    assign in10175_1 = {c7820};
    assign in10175_2 = {s7821[0]};
    Full_Adder FA_10175(s10175, c10175, in10175_1, in10175_2, c7819);
    wire[0:0] s10176, in10176_1, in10176_2;
    wire c10176;
    assign in10176_1 = {s7823[0]};
    assign in10176_2 = {s7824[0]};
    Full_Adder FA_10176(s10176, c10176, in10176_1, in10176_2, s7822[0]);
    wire[0:0] s10177, in10177_1, in10177_2;
    wire c10177;
    assign in10177_1 = {s7826[0]};
    assign in10177_2 = {s7827[0]};
    Full_Adder FA_10177(s10177, c10177, in10177_1, in10177_2, s7825[0]);
    wire[0:0] s10178, in10178_1, in10178_2;
    wire c10178;
    assign in10178_1 = {s7829[0]};
    assign in10178_2 = {s7830[0]};
    Full_Adder FA_10178(s10178, c10178, in10178_1, in10178_2, s7828[0]);
    wire[0:0] s10179, in10179_1, in10179_2;
    wire c10179;
    assign in10179_1 = {s7832[0]};
    assign in10179_2 = {s7833[0]};
    Full_Adder FA_10179(s10179, c10179, in10179_1, in10179_2, s7831[0]);
    wire[0:0] s10180, in10180_1, in10180_2;
    wire c10180;
    assign in10180_1 = {s7835[0]};
    assign in10180_2 = {s7836[0]};
    Full_Adder FA_10180(s10180, c10180, in10180_1, in10180_2, s7834[0]);
    wire[0:0] s10181, in10181_1, in10181_2;
    wire c10181;
    assign in10181_1 = {s7838[0]};
    assign in10181_2 = {s7839[0]};
    Full_Adder FA_10181(s10181, c10181, in10181_1, in10181_2, s7837[0]);
    wire[0:0] s10182, in10182_1, in10182_2;
    wire c10182;
    assign in10182_1 = {pp127[72]};
    assign in10182_2 = {c7821};
    Full_Adder FA_10182(s10182, c10182, in10182_1, in10182_2, pp126[73]);
    wire[0:0] s10183, in10183_1, in10183_2;
    wire c10183;
    assign in10183_1 = {c7823};
    assign in10183_2 = {c7824};
    Full_Adder FA_10183(s10183, c10183, in10183_1, in10183_2, c7822);
    wire[0:0] s10184, in10184_1, in10184_2;
    wire c10184;
    assign in10184_1 = {c7826};
    assign in10184_2 = {c7827};
    Full_Adder FA_10184(s10184, c10184, in10184_1, in10184_2, c7825);
    wire[0:0] s10185, in10185_1, in10185_2;
    wire c10185;
    assign in10185_1 = {c7829};
    assign in10185_2 = {c7830};
    Full_Adder FA_10185(s10185, c10185, in10185_1, in10185_2, c7828);
    wire[0:0] s10186, in10186_1, in10186_2;
    wire c10186;
    assign in10186_1 = {c7832};
    assign in10186_2 = {c7833};
    Full_Adder FA_10186(s10186, c10186, in10186_1, in10186_2, c7831);
    wire[0:0] s10187, in10187_1, in10187_2;
    wire c10187;
    assign in10187_1 = {c7835};
    assign in10187_2 = {c7836};
    Full_Adder FA_10187(s10187, c10187, in10187_1, in10187_2, c7834);
    wire[0:0] s10188, in10188_1, in10188_2;
    wire c10188;
    assign in10188_1 = {c7838};
    assign in10188_2 = {c7839};
    Full_Adder FA_10188(s10188, c10188, in10188_1, in10188_2, c7837);
    wire[0:0] s10189, in10189_1, in10189_2;
    wire c10189;
    assign in10189_1 = {s7841[0]};
    assign in10189_2 = {s7842[0]};
    Full_Adder FA_10189(s10189, c10189, in10189_1, in10189_2, s7840[0]);
    wire[0:0] s10190, in10190_1, in10190_2;
    wire c10190;
    assign in10190_1 = {s7844[0]};
    assign in10190_2 = {s7845[0]};
    Full_Adder FA_10190(s10190, c10190, in10190_1, in10190_2, s7843[0]);
    wire[0:0] s10191, in10191_1, in10191_2;
    wire c10191;
    assign in10191_1 = {s7847[0]};
    assign in10191_2 = {s7848[0]};
    Full_Adder FA_10191(s10191, c10191, in10191_1, in10191_2, s7846[0]);
    wire[0:0] s10192, in10192_1, in10192_2;
    wire c10192;
    assign in10192_1 = {s7850[0]};
    assign in10192_2 = {s7851[0]};
    Full_Adder FA_10192(s10192, c10192, in10192_1, in10192_2, s7849[0]);
    wire[0:0] s10193, in10193_1, in10193_2;
    wire c10193;
    assign in10193_1 = {s7853[0]};
    assign in10193_2 = {s7854[0]};
    Full_Adder FA_10193(s10193, c10193, in10193_1, in10193_2, s7852[0]);
    wire[0:0] s10194, in10194_1, in10194_2;
    wire c10194;
    assign in10194_1 = {s7856[0]};
    assign in10194_2 = {s7857[0]};
    Full_Adder FA_10194(s10194, c10194, in10194_1, in10194_2, s7855[0]);
    wire[0:0] s10195, in10195_1, in10195_2;
    wire c10195;
    assign in10195_1 = {pp125[75]};
    assign in10195_2 = {pp126[74]};
    Full_Adder FA_10195(s10195, c10195, in10195_1, in10195_2, pp124[76]);
    wire[0:0] s10196, in10196_1, in10196_2;
    wire c10196;
    assign in10196_1 = {c7840};
    assign in10196_2 = {c7841};
    Full_Adder FA_10196(s10196, c10196, in10196_1, in10196_2, pp127[73]);
    wire[0:0] s10197, in10197_1, in10197_2;
    wire c10197;
    assign in10197_1 = {c7843};
    assign in10197_2 = {c7844};
    Full_Adder FA_10197(s10197, c10197, in10197_1, in10197_2, c7842);
    wire[0:0] s10198, in10198_1, in10198_2;
    wire c10198;
    assign in10198_1 = {c7846};
    assign in10198_2 = {c7847};
    Full_Adder FA_10198(s10198, c10198, in10198_1, in10198_2, c7845);
    wire[0:0] s10199, in10199_1, in10199_2;
    wire c10199;
    assign in10199_1 = {c7849};
    assign in10199_2 = {c7850};
    Full_Adder FA_10199(s10199, c10199, in10199_1, in10199_2, c7848);
    wire[0:0] s10200, in10200_1, in10200_2;
    wire c10200;
    assign in10200_1 = {c7852};
    assign in10200_2 = {c7853};
    Full_Adder FA_10200(s10200, c10200, in10200_1, in10200_2, c7851);
    wire[0:0] s10201, in10201_1, in10201_2;
    wire c10201;
    assign in10201_1 = {c7855};
    assign in10201_2 = {c7856};
    Full_Adder FA_10201(s10201, c10201, in10201_1, in10201_2, c7854);
    wire[0:0] s10202, in10202_1, in10202_2;
    wire c10202;
    assign in10202_1 = {s7858[0]};
    assign in10202_2 = {s7859[0]};
    Full_Adder FA_10202(s10202, c10202, in10202_1, in10202_2, c7857);
    wire[0:0] s10203, in10203_1, in10203_2;
    wire c10203;
    assign in10203_1 = {s7861[0]};
    assign in10203_2 = {s7862[0]};
    Full_Adder FA_10203(s10203, c10203, in10203_1, in10203_2, s7860[0]);
    wire[0:0] s10204, in10204_1, in10204_2;
    wire c10204;
    assign in10204_1 = {s7864[0]};
    assign in10204_2 = {s7865[0]};
    Full_Adder FA_10204(s10204, c10204, in10204_1, in10204_2, s7863[0]);
    wire[0:0] s10205, in10205_1, in10205_2;
    wire c10205;
    assign in10205_1 = {s7867[0]};
    assign in10205_2 = {s7868[0]};
    Full_Adder FA_10205(s10205, c10205, in10205_1, in10205_2, s7866[0]);
    wire[0:0] s10206, in10206_1, in10206_2;
    wire c10206;
    assign in10206_1 = {s7870[0]};
    assign in10206_2 = {s7871[0]};
    Full_Adder FA_10206(s10206, c10206, in10206_1, in10206_2, s7869[0]);
    wire[0:0] s10207, in10207_1, in10207_2;
    wire c10207;
    assign in10207_1 = {s7873[0]};
    assign in10207_2 = {s7874[0]};
    Full_Adder FA_10207(s10207, c10207, in10207_1, in10207_2, s7872[0]);
    wire[0:0] s10208, in10208_1, in10208_2;
    wire c10208;
    assign in10208_1 = {pp123[78]};
    assign in10208_2 = {pp124[77]};
    Full_Adder FA_10208(s10208, c10208, in10208_1, in10208_2, pp122[79]);
    wire[0:0] s10209, in10209_1, in10209_2;
    wire c10209;
    assign in10209_1 = {pp126[75]};
    assign in10209_2 = {pp127[74]};
    Full_Adder FA_10209(s10209, c10209, in10209_1, in10209_2, pp125[76]);
    wire[0:0] s10210, in10210_1, in10210_2;
    wire c10210;
    assign in10210_1 = {c7859};
    assign in10210_2 = {c7860};
    Full_Adder FA_10210(s10210, c10210, in10210_1, in10210_2, c7858);
    wire[0:0] s10211, in10211_1, in10211_2;
    wire c10211;
    assign in10211_1 = {c7862};
    assign in10211_2 = {c7863};
    Full_Adder FA_10211(s10211, c10211, in10211_1, in10211_2, c7861);
    wire[0:0] s10212, in10212_1, in10212_2;
    wire c10212;
    assign in10212_1 = {c7865};
    assign in10212_2 = {c7866};
    Full_Adder FA_10212(s10212, c10212, in10212_1, in10212_2, c7864);
    wire[0:0] s10213, in10213_1, in10213_2;
    wire c10213;
    assign in10213_1 = {c7868};
    assign in10213_2 = {c7869};
    Full_Adder FA_10213(s10213, c10213, in10213_1, in10213_2, c7867);
    wire[0:0] s10214, in10214_1, in10214_2;
    wire c10214;
    assign in10214_1 = {c7871};
    assign in10214_2 = {c7872};
    Full_Adder FA_10214(s10214, c10214, in10214_1, in10214_2, c7870);
    wire[0:0] s10215, in10215_1, in10215_2;
    wire c10215;
    assign in10215_1 = {c7874};
    assign in10215_2 = {s7875[0]};
    Full_Adder FA_10215(s10215, c10215, in10215_1, in10215_2, c7873);
    wire[0:0] s10216, in10216_1, in10216_2;
    wire c10216;
    assign in10216_1 = {s7877[0]};
    assign in10216_2 = {s7878[0]};
    Full_Adder FA_10216(s10216, c10216, in10216_1, in10216_2, s7876[0]);
    wire[0:0] s10217, in10217_1, in10217_2;
    wire c10217;
    assign in10217_1 = {s7880[0]};
    assign in10217_2 = {s7881[0]};
    Full_Adder FA_10217(s10217, c10217, in10217_1, in10217_2, s7879[0]);
    wire[0:0] s10218, in10218_1, in10218_2;
    wire c10218;
    assign in10218_1 = {s7883[0]};
    assign in10218_2 = {s7884[0]};
    Full_Adder FA_10218(s10218, c10218, in10218_1, in10218_2, s7882[0]);
    wire[0:0] s10219, in10219_1, in10219_2;
    wire c10219;
    assign in10219_1 = {s7886[0]};
    assign in10219_2 = {s7887[0]};
    Full_Adder FA_10219(s10219, c10219, in10219_1, in10219_2, s7885[0]);
    wire[0:0] s10220, in10220_1, in10220_2;
    wire c10220;
    assign in10220_1 = {s7889[0]};
    assign in10220_2 = {s7890[0]};
    Full_Adder FA_10220(s10220, c10220, in10220_1, in10220_2, s7888[0]);
    wire[0:0] s10221, in10221_1, in10221_2;
    wire c10221;
    assign in10221_1 = {pp121[81]};
    assign in10221_2 = {pp122[80]};
    Full_Adder FA_10221(s10221, c10221, in10221_1, in10221_2, pp120[82]);
    wire[0:0] s10222, in10222_1, in10222_2;
    wire c10222;
    assign in10222_1 = {pp124[78]};
    assign in10222_2 = {pp125[77]};
    Full_Adder FA_10222(s10222, c10222, in10222_1, in10222_2, pp123[79]);
    wire[0:0] s10223, in10223_1, in10223_2;
    wire c10223;
    assign in10223_1 = {pp127[75]};
    assign in10223_2 = {c7875};
    Full_Adder FA_10223(s10223, c10223, in10223_1, in10223_2, pp126[76]);
    wire[0:0] s10224, in10224_1, in10224_2;
    wire c10224;
    assign in10224_1 = {c7877};
    assign in10224_2 = {c7878};
    Full_Adder FA_10224(s10224, c10224, in10224_1, in10224_2, c7876);
    wire[0:0] s10225, in10225_1, in10225_2;
    wire c10225;
    assign in10225_1 = {c7880};
    assign in10225_2 = {c7881};
    Full_Adder FA_10225(s10225, c10225, in10225_1, in10225_2, c7879);
    wire[0:0] s10226, in10226_1, in10226_2;
    wire c10226;
    assign in10226_1 = {c7883};
    assign in10226_2 = {c7884};
    Full_Adder FA_10226(s10226, c10226, in10226_1, in10226_2, c7882);
    wire[0:0] s10227, in10227_1, in10227_2;
    wire c10227;
    assign in10227_1 = {c7886};
    assign in10227_2 = {c7887};
    Full_Adder FA_10227(s10227, c10227, in10227_1, in10227_2, c7885);
    wire[0:0] s10228, in10228_1, in10228_2;
    wire c10228;
    assign in10228_1 = {c7889};
    assign in10228_2 = {c7890};
    Full_Adder FA_10228(s10228, c10228, in10228_1, in10228_2, c7888);
    wire[0:0] s10229, in10229_1, in10229_2;
    wire c10229;
    assign in10229_1 = {s7892[0]};
    assign in10229_2 = {s7893[0]};
    Full_Adder FA_10229(s10229, c10229, in10229_1, in10229_2, s7891[0]);
    wire[0:0] s10230, in10230_1, in10230_2;
    wire c10230;
    assign in10230_1 = {s7895[0]};
    assign in10230_2 = {s7896[0]};
    Full_Adder FA_10230(s10230, c10230, in10230_1, in10230_2, s7894[0]);
    wire[0:0] s10231, in10231_1, in10231_2;
    wire c10231;
    assign in10231_1 = {s7898[0]};
    assign in10231_2 = {s7899[0]};
    Full_Adder FA_10231(s10231, c10231, in10231_1, in10231_2, s7897[0]);
    wire[0:0] s10232, in10232_1, in10232_2;
    wire c10232;
    assign in10232_1 = {s7901[0]};
    assign in10232_2 = {s7902[0]};
    Full_Adder FA_10232(s10232, c10232, in10232_1, in10232_2, s7900[0]);
    wire[0:0] s10233, in10233_1, in10233_2;
    wire c10233;
    assign in10233_1 = {s7904[0]};
    assign in10233_2 = {s7905[0]};
    Full_Adder FA_10233(s10233, c10233, in10233_1, in10233_2, s7903[0]);
    wire[0:0] s10234, in10234_1, in10234_2;
    wire c10234;
    assign in10234_1 = {pp119[84]};
    assign in10234_2 = {pp120[83]};
    Full_Adder FA_10234(s10234, c10234, in10234_1, in10234_2, pp118[85]);
    wire[0:0] s10235, in10235_1, in10235_2;
    wire c10235;
    assign in10235_1 = {pp122[81]};
    assign in10235_2 = {pp123[80]};
    Full_Adder FA_10235(s10235, c10235, in10235_1, in10235_2, pp121[82]);
    wire[0:0] s10236, in10236_1, in10236_2;
    wire c10236;
    assign in10236_1 = {pp125[78]};
    assign in10236_2 = {pp126[77]};
    Full_Adder FA_10236(s10236, c10236, in10236_1, in10236_2, pp124[79]);
    wire[0:0] s10237, in10237_1, in10237_2;
    wire c10237;
    assign in10237_1 = {c7891};
    assign in10237_2 = {c7892};
    Full_Adder FA_10237(s10237, c10237, in10237_1, in10237_2, pp127[76]);
    wire[0:0] s10238, in10238_1, in10238_2;
    wire c10238;
    assign in10238_1 = {c7894};
    assign in10238_2 = {c7895};
    Full_Adder FA_10238(s10238, c10238, in10238_1, in10238_2, c7893);
    wire[0:0] s10239, in10239_1, in10239_2;
    wire c10239;
    assign in10239_1 = {c7897};
    assign in10239_2 = {c7898};
    Full_Adder FA_10239(s10239, c10239, in10239_1, in10239_2, c7896);
    wire[0:0] s10240, in10240_1, in10240_2;
    wire c10240;
    assign in10240_1 = {c7900};
    assign in10240_2 = {c7901};
    Full_Adder FA_10240(s10240, c10240, in10240_1, in10240_2, c7899);
    wire[0:0] s10241, in10241_1, in10241_2;
    wire c10241;
    assign in10241_1 = {c7903};
    assign in10241_2 = {c7904};
    Full_Adder FA_10241(s10241, c10241, in10241_1, in10241_2, c7902);
    wire[0:0] s10242, in10242_1, in10242_2;
    wire c10242;
    assign in10242_1 = {s7906[0]};
    assign in10242_2 = {s7907[0]};
    Full_Adder FA_10242(s10242, c10242, in10242_1, in10242_2, c7905);
    wire[0:0] s10243, in10243_1, in10243_2;
    wire c10243;
    assign in10243_1 = {s7909[0]};
    assign in10243_2 = {s7910[0]};
    Full_Adder FA_10243(s10243, c10243, in10243_1, in10243_2, s7908[0]);
    wire[0:0] s10244, in10244_1, in10244_2;
    wire c10244;
    assign in10244_1 = {s7912[0]};
    assign in10244_2 = {s7913[0]};
    Full_Adder FA_10244(s10244, c10244, in10244_1, in10244_2, s7911[0]);
    wire[0:0] s10245, in10245_1, in10245_2;
    wire c10245;
    assign in10245_1 = {s7915[0]};
    assign in10245_2 = {s7916[0]};
    Full_Adder FA_10245(s10245, c10245, in10245_1, in10245_2, s7914[0]);
    wire[0:0] s10246, in10246_1, in10246_2;
    wire c10246;
    assign in10246_1 = {s7918[0]};
    assign in10246_2 = {s7919[0]};
    Full_Adder FA_10246(s10246, c10246, in10246_1, in10246_2, s7917[0]);
    wire[0:0] s10247, in10247_1, in10247_2;
    wire c10247;
    assign in10247_1 = {pp117[87]};
    assign in10247_2 = {pp118[86]};
    Full_Adder FA_10247(s10247, c10247, in10247_1, in10247_2, pp116[88]);
    wire[0:0] s10248, in10248_1, in10248_2;
    wire c10248;
    assign in10248_1 = {pp120[84]};
    assign in10248_2 = {pp121[83]};
    Full_Adder FA_10248(s10248, c10248, in10248_1, in10248_2, pp119[85]);
    wire[0:0] s10249, in10249_1, in10249_2;
    wire c10249;
    assign in10249_1 = {pp123[81]};
    assign in10249_2 = {pp124[80]};
    Full_Adder FA_10249(s10249, c10249, in10249_1, in10249_2, pp122[82]);
    wire[0:0] s10250, in10250_1, in10250_2;
    wire c10250;
    assign in10250_1 = {pp126[78]};
    assign in10250_2 = {pp127[77]};
    Full_Adder FA_10250(s10250, c10250, in10250_1, in10250_2, pp125[79]);
    wire[0:0] s10251, in10251_1, in10251_2;
    wire c10251;
    assign in10251_1 = {c7907};
    assign in10251_2 = {c7908};
    Full_Adder FA_10251(s10251, c10251, in10251_1, in10251_2, c7906);
    wire[0:0] s10252, in10252_1, in10252_2;
    wire c10252;
    assign in10252_1 = {c7910};
    assign in10252_2 = {c7911};
    Full_Adder FA_10252(s10252, c10252, in10252_1, in10252_2, c7909);
    wire[0:0] s10253, in10253_1, in10253_2;
    wire c10253;
    assign in10253_1 = {c7913};
    assign in10253_2 = {c7914};
    Full_Adder FA_10253(s10253, c10253, in10253_1, in10253_2, c7912);
    wire[0:0] s10254, in10254_1, in10254_2;
    wire c10254;
    assign in10254_1 = {c7916};
    assign in10254_2 = {c7917};
    Full_Adder FA_10254(s10254, c10254, in10254_1, in10254_2, c7915);
    wire[0:0] s10255, in10255_1, in10255_2;
    wire c10255;
    assign in10255_1 = {c7919};
    assign in10255_2 = {s7920[0]};
    Full_Adder FA_10255(s10255, c10255, in10255_1, in10255_2, c7918);
    wire[0:0] s10256, in10256_1, in10256_2;
    wire c10256;
    assign in10256_1 = {s7922[0]};
    assign in10256_2 = {s7923[0]};
    Full_Adder FA_10256(s10256, c10256, in10256_1, in10256_2, s7921[0]);
    wire[0:0] s10257, in10257_1, in10257_2;
    wire c10257;
    assign in10257_1 = {s7925[0]};
    assign in10257_2 = {s7926[0]};
    Full_Adder FA_10257(s10257, c10257, in10257_1, in10257_2, s7924[0]);
    wire[0:0] s10258, in10258_1, in10258_2;
    wire c10258;
    assign in10258_1 = {s7928[0]};
    assign in10258_2 = {s7929[0]};
    Full_Adder FA_10258(s10258, c10258, in10258_1, in10258_2, s7927[0]);
    wire[0:0] s10259, in10259_1, in10259_2;
    wire c10259;
    assign in10259_1 = {s7931[0]};
    assign in10259_2 = {s7932[0]};
    Full_Adder FA_10259(s10259, c10259, in10259_1, in10259_2, s7930[0]);
    wire[0:0] s10260, in10260_1, in10260_2;
    wire c10260;
    assign in10260_1 = {pp115[90]};
    assign in10260_2 = {pp116[89]};
    Full_Adder FA_10260(s10260, c10260, in10260_1, in10260_2, pp114[91]);
    wire[0:0] s10261, in10261_1, in10261_2;
    wire c10261;
    assign in10261_1 = {pp118[87]};
    assign in10261_2 = {pp119[86]};
    Full_Adder FA_10261(s10261, c10261, in10261_1, in10261_2, pp117[88]);
    wire[0:0] s10262, in10262_1, in10262_2;
    wire c10262;
    assign in10262_1 = {pp121[84]};
    assign in10262_2 = {pp122[83]};
    Full_Adder FA_10262(s10262, c10262, in10262_1, in10262_2, pp120[85]);
    wire[0:0] s10263, in10263_1, in10263_2;
    wire c10263;
    assign in10263_1 = {pp124[81]};
    assign in10263_2 = {pp125[80]};
    Full_Adder FA_10263(s10263, c10263, in10263_1, in10263_2, pp123[82]);
    wire[0:0] s10264, in10264_1, in10264_2;
    wire c10264;
    assign in10264_1 = {pp127[78]};
    assign in10264_2 = {c7920};
    Full_Adder FA_10264(s10264, c10264, in10264_1, in10264_2, pp126[79]);
    wire[0:0] s10265, in10265_1, in10265_2;
    wire c10265;
    assign in10265_1 = {c7922};
    assign in10265_2 = {c7923};
    Full_Adder FA_10265(s10265, c10265, in10265_1, in10265_2, c7921);
    wire[0:0] s10266, in10266_1, in10266_2;
    wire c10266;
    assign in10266_1 = {c7925};
    assign in10266_2 = {c7926};
    Full_Adder FA_10266(s10266, c10266, in10266_1, in10266_2, c7924);
    wire[0:0] s10267, in10267_1, in10267_2;
    wire c10267;
    assign in10267_1 = {c7928};
    assign in10267_2 = {c7929};
    Full_Adder FA_10267(s10267, c10267, in10267_1, in10267_2, c7927);
    wire[0:0] s10268, in10268_1, in10268_2;
    wire c10268;
    assign in10268_1 = {c7931};
    assign in10268_2 = {c7932};
    Full_Adder FA_10268(s10268, c10268, in10268_1, in10268_2, c7930);
    wire[0:0] s10269, in10269_1, in10269_2;
    wire c10269;
    assign in10269_1 = {s7934[0]};
    assign in10269_2 = {s7935[0]};
    Full_Adder FA_10269(s10269, c10269, in10269_1, in10269_2, s7933[0]);
    wire[0:0] s10270, in10270_1, in10270_2;
    wire c10270;
    assign in10270_1 = {s7937[0]};
    assign in10270_2 = {s7938[0]};
    Full_Adder FA_10270(s10270, c10270, in10270_1, in10270_2, s7936[0]);
    wire[0:0] s10271, in10271_1, in10271_2;
    wire c10271;
    assign in10271_1 = {s7940[0]};
    assign in10271_2 = {s7941[0]};
    Full_Adder FA_10271(s10271, c10271, in10271_1, in10271_2, s7939[0]);
    wire[0:0] s10272, in10272_1, in10272_2;
    wire c10272;
    assign in10272_1 = {s7943[0]};
    assign in10272_2 = {s7944[0]};
    Full_Adder FA_10272(s10272, c10272, in10272_1, in10272_2, s7942[0]);
    wire[0:0] s10273, in10273_1, in10273_2;
    wire c10273;
    assign in10273_1 = {pp113[93]};
    assign in10273_2 = {pp114[92]};
    Full_Adder FA_10273(s10273, c10273, in10273_1, in10273_2, pp112[94]);
    wire[0:0] s10274, in10274_1, in10274_2;
    wire c10274;
    assign in10274_1 = {pp116[90]};
    assign in10274_2 = {pp117[89]};
    Full_Adder FA_10274(s10274, c10274, in10274_1, in10274_2, pp115[91]);
    wire[0:0] s10275, in10275_1, in10275_2;
    wire c10275;
    assign in10275_1 = {pp119[87]};
    assign in10275_2 = {pp120[86]};
    Full_Adder FA_10275(s10275, c10275, in10275_1, in10275_2, pp118[88]);
    wire[0:0] s10276, in10276_1, in10276_2;
    wire c10276;
    assign in10276_1 = {pp122[84]};
    assign in10276_2 = {pp123[83]};
    Full_Adder FA_10276(s10276, c10276, in10276_1, in10276_2, pp121[85]);
    wire[0:0] s10277, in10277_1, in10277_2;
    wire c10277;
    assign in10277_1 = {pp125[81]};
    assign in10277_2 = {pp126[80]};
    Full_Adder FA_10277(s10277, c10277, in10277_1, in10277_2, pp124[82]);
    wire[0:0] s10278, in10278_1, in10278_2;
    wire c10278;
    assign in10278_1 = {c7933};
    assign in10278_2 = {c7934};
    Full_Adder FA_10278(s10278, c10278, in10278_1, in10278_2, pp127[79]);
    wire[0:0] s10279, in10279_1, in10279_2;
    wire c10279;
    assign in10279_1 = {c7936};
    assign in10279_2 = {c7937};
    Full_Adder FA_10279(s10279, c10279, in10279_1, in10279_2, c7935);
    wire[0:0] s10280, in10280_1, in10280_2;
    wire c10280;
    assign in10280_1 = {c7939};
    assign in10280_2 = {c7940};
    Full_Adder FA_10280(s10280, c10280, in10280_1, in10280_2, c7938);
    wire[0:0] s10281, in10281_1, in10281_2;
    wire c10281;
    assign in10281_1 = {c7942};
    assign in10281_2 = {c7943};
    Full_Adder FA_10281(s10281, c10281, in10281_1, in10281_2, c7941);
    wire[0:0] s10282, in10282_1, in10282_2;
    wire c10282;
    assign in10282_1 = {s7945[0]};
    assign in10282_2 = {s7946[0]};
    Full_Adder FA_10282(s10282, c10282, in10282_1, in10282_2, c7944);
    wire[0:0] s10283, in10283_1, in10283_2;
    wire c10283;
    assign in10283_1 = {s7948[0]};
    assign in10283_2 = {s7949[0]};
    Full_Adder FA_10283(s10283, c10283, in10283_1, in10283_2, s7947[0]);
    wire[0:0] s10284, in10284_1, in10284_2;
    wire c10284;
    assign in10284_1 = {s7951[0]};
    assign in10284_2 = {s7952[0]};
    Full_Adder FA_10284(s10284, c10284, in10284_1, in10284_2, s7950[0]);
    wire[0:0] s10285, in10285_1, in10285_2;
    wire c10285;
    assign in10285_1 = {s7954[0]};
    assign in10285_2 = {s7955[0]};
    Full_Adder FA_10285(s10285, c10285, in10285_1, in10285_2, s7953[0]);
    wire[0:0] s10286, in10286_1, in10286_2;
    wire c10286;
    assign in10286_1 = {pp111[96]};
    assign in10286_2 = {pp112[95]};
    Full_Adder FA_10286(s10286, c10286, in10286_1, in10286_2, pp110[97]);
    wire[0:0] s10287, in10287_1, in10287_2;
    wire c10287;
    assign in10287_1 = {pp114[93]};
    assign in10287_2 = {pp115[92]};
    Full_Adder FA_10287(s10287, c10287, in10287_1, in10287_2, pp113[94]);
    wire[0:0] s10288, in10288_1, in10288_2;
    wire c10288;
    assign in10288_1 = {pp117[90]};
    assign in10288_2 = {pp118[89]};
    Full_Adder FA_10288(s10288, c10288, in10288_1, in10288_2, pp116[91]);
    wire[0:0] s10289, in10289_1, in10289_2;
    wire c10289;
    assign in10289_1 = {pp120[87]};
    assign in10289_2 = {pp121[86]};
    Full_Adder FA_10289(s10289, c10289, in10289_1, in10289_2, pp119[88]);
    wire[0:0] s10290, in10290_1, in10290_2;
    wire c10290;
    assign in10290_1 = {pp123[84]};
    assign in10290_2 = {pp124[83]};
    Full_Adder FA_10290(s10290, c10290, in10290_1, in10290_2, pp122[85]);
    wire[0:0] s10291, in10291_1, in10291_2;
    wire c10291;
    assign in10291_1 = {pp126[81]};
    assign in10291_2 = {pp127[80]};
    Full_Adder FA_10291(s10291, c10291, in10291_1, in10291_2, pp125[82]);
    wire[0:0] s10292, in10292_1, in10292_2;
    wire c10292;
    assign in10292_1 = {c7946};
    assign in10292_2 = {c7947};
    Full_Adder FA_10292(s10292, c10292, in10292_1, in10292_2, c7945);
    wire[0:0] s10293, in10293_1, in10293_2;
    wire c10293;
    assign in10293_1 = {c7949};
    assign in10293_2 = {c7950};
    Full_Adder FA_10293(s10293, c10293, in10293_1, in10293_2, c7948);
    wire[0:0] s10294, in10294_1, in10294_2;
    wire c10294;
    assign in10294_1 = {c7952};
    assign in10294_2 = {c7953};
    Full_Adder FA_10294(s10294, c10294, in10294_1, in10294_2, c7951);
    wire[0:0] s10295, in10295_1, in10295_2;
    wire c10295;
    assign in10295_1 = {c7955};
    assign in10295_2 = {s7956[0]};
    Full_Adder FA_10295(s10295, c10295, in10295_1, in10295_2, c7954);
    wire[0:0] s10296, in10296_1, in10296_2;
    wire c10296;
    assign in10296_1 = {s7958[0]};
    assign in10296_2 = {s7959[0]};
    Full_Adder FA_10296(s10296, c10296, in10296_1, in10296_2, s7957[0]);
    wire[0:0] s10297, in10297_1, in10297_2;
    wire c10297;
    assign in10297_1 = {s7961[0]};
    assign in10297_2 = {s7962[0]};
    Full_Adder FA_10297(s10297, c10297, in10297_1, in10297_2, s7960[0]);
    wire[0:0] s10298, in10298_1, in10298_2;
    wire c10298;
    assign in10298_1 = {s7964[0]};
    assign in10298_2 = {s7965[0]};
    Full_Adder FA_10298(s10298, c10298, in10298_1, in10298_2, s7963[0]);
    wire[0:0] s10299, in10299_1, in10299_2;
    wire c10299;
    assign in10299_1 = {pp109[99]};
    assign in10299_2 = {pp110[98]};
    Full_Adder FA_10299(s10299, c10299, in10299_1, in10299_2, pp108[100]);
    wire[0:0] s10300, in10300_1, in10300_2;
    wire c10300;
    assign in10300_1 = {pp112[96]};
    assign in10300_2 = {pp113[95]};
    Full_Adder FA_10300(s10300, c10300, in10300_1, in10300_2, pp111[97]);
    wire[0:0] s10301, in10301_1, in10301_2;
    wire c10301;
    assign in10301_1 = {pp115[93]};
    assign in10301_2 = {pp116[92]};
    Full_Adder FA_10301(s10301, c10301, in10301_1, in10301_2, pp114[94]);
    wire[0:0] s10302, in10302_1, in10302_2;
    wire c10302;
    assign in10302_1 = {pp118[90]};
    assign in10302_2 = {pp119[89]};
    Full_Adder FA_10302(s10302, c10302, in10302_1, in10302_2, pp117[91]);
    wire[0:0] s10303, in10303_1, in10303_2;
    wire c10303;
    assign in10303_1 = {pp121[87]};
    assign in10303_2 = {pp122[86]};
    Full_Adder FA_10303(s10303, c10303, in10303_1, in10303_2, pp120[88]);
    wire[0:0] s10304, in10304_1, in10304_2;
    wire c10304;
    assign in10304_1 = {pp124[84]};
    assign in10304_2 = {pp125[83]};
    Full_Adder FA_10304(s10304, c10304, in10304_1, in10304_2, pp123[85]);
    wire[0:0] s10305, in10305_1, in10305_2;
    wire c10305;
    assign in10305_1 = {pp127[81]};
    assign in10305_2 = {c7956};
    Full_Adder FA_10305(s10305, c10305, in10305_1, in10305_2, pp126[82]);
    wire[0:0] s10306, in10306_1, in10306_2;
    wire c10306;
    assign in10306_1 = {c7958};
    assign in10306_2 = {c7959};
    Full_Adder FA_10306(s10306, c10306, in10306_1, in10306_2, c7957);
    wire[0:0] s10307, in10307_1, in10307_2;
    wire c10307;
    assign in10307_1 = {c7961};
    assign in10307_2 = {c7962};
    Full_Adder FA_10307(s10307, c10307, in10307_1, in10307_2, c7960);
    wire[0:0] s10308, in10308_1, in10308_2;
    wire c10308;
    assign in10308_1 = {c7964};
    assign in10308_2 = {c7965};
    Full_Adder FA_10308(s10308, c10308, in10308_1, in10308_2, c7963);
    wire[0:0] s10309, in10309_1, in10309_2;
    wire c10309;
    assign in10309_1 = {s7967[0]};
    assign in10309_2 = {s7968[0]};
    Full_Adder FA_10309(s10309, c10309, in10309_1, in10309_2, s7966[0]);
    wire[0:0] s10310, in10310_1, in10310_2;
    wire c10310;
    assign in10310_1 = {s7970[0]};
    assign in10310_2 = {s7971[0]};
    Full_Adder FA_10310(s10310, c10310, in10310_1, in10310_2, s7969[0]);
    wire[0:0] s10311, in10311_1, in10311_2;
    wire c10311;
    assign in10311_1 = {s7973[0]};
    assign in10311_2 = {s7974[0]};
    Full_Adder FA_10311(s10311, c10311, in10311_1, in10311_2, s7972[0]);
    wire[0:0] s10312, in10312_1, in10312_2;
    wire c10312;
    assign in10312_1 = {pp107[102]};
    assign in10312_2 = {pp108[101]};
    Full_Adder FA_10312(s10312, c10312, in10312_1, in10312_2, pp106[103]);
    wire[0:0] s10313, in10313_1, in10313_2;
    wire c10313;
    assign in10313_1 = {pp110[99]};
    assign in10313_2 = {pp111[98]};
    Full_Adder FA_10313(s10313, c10313, in10313_1, in10313_2, pp109[100]);
    wire[0:0] s10314, in10314_1, in10314_2;
    wire c10314;
    assign in10314_1 = {pp113[96]};
    assign in10314_2 = {pp114[95]};
    Full_Adder FA_10314(s10314, c10314, in10314_1, in10314_2, pp112[97]);
    wire[0:0] s10315, in10315_1, in10315_2;
    wire c10315;
    assign in10315_1 = {pp116[93]};
    assign in10315_2 = {pp117[92]};
    Full_Adder FA_10315(s10315, c10315, in10315_1, in10315_2, pp115[94]);
    wire[0:0] s10316, in10316_1, in10316_2;
    wire c10316;
    assign in10316_1 = {pp119[90]};
    assign in10316_2 = {pp120[89]};
    Full_Adder FA_10316(s10316, c10316, in10316_1, in10316_2, pp118[91]);
    wire[0:0] s10317, in10317_1, in10317_2;
    wire c10317;
    assign in10317_1 = {pp122[87]};
    assign in10317_2 = {pp123[86]};
    Full_Adder FA_10317(s10317, c10317, in10317_1, in10317_2, pp121[88]);
    wire[0:0] s10318, in10318_1, in10318_2;
    wire c10318;
    assign in10318_1 = {pp125[84]};
    assign in10318_2 = {pp126[83]};
    Full_Adder FA_10318(s10318, c10318, in10318_1, in10318_2, pp124[85]);
    wire[0:0] s10319, in10319_1, in10319_2;
    wire c10319;
    assign in10319_1 = {c7966};
    assign in10319_2 = {c7967};
    Full_Adder FA_10319(s10319, c10319, in10319_1, in10319_2, pp127[82]);
    wire[0:0] s10320, in10320_1, in10320_2;
    wire c10320;
    assign in10320_1 = {c7969};
    assign in10320_2 = {c7970};
    Full_Adder FA_10320(s10320, c10320, in10320_1, in10320_2, c7968);
    wire[0:0] s10321, in10321_1, in10321_2;
    wire c10321;
    assign in10321_1 = {c7972};
    assign in10321_2 = {c7973};
    Full_Adder FA_10321(s10321, c10321, in10321_1, in10321_2, c7971);
    wire[0:0] s10322, in10322_1, in10322_2;
    wire c10322;
    assign in10322_1 = {s7975[0]};
    assign in10322_2 = {s7976[0]};
    Full_Adder FA_10322(s10322, c10322, in10322_1, in10322_2, c7974);
    wire[0:0] s10323, in10323_1, in10323_2;
    wire c10323;
    assign in10323_1 = {s7978[0]};
    assign in10323_2 = {s7979[0]};
    Full_Adder FA_10323(s10323, c10323, in10323_1, in10323_2, s7977[0]);
    wire[0:0] s10324, in10324_1, in10324_2;
    wire c10324;
    assign in10324_1 = {s7981[0]};
    assign in10324_2 = {s7982[0]};
    Full_Adder FA_10324(s10324, c10324, in10324_1, in10324_2, s7980[0]);
    wire[0:0] s10325, in10325_1, in10325_2;
    wire c10325;
    assign in10325_1 = {pp105[105]};
    assign in10325_2 = {pp106[104]};
    Full_Adder FA_10325(s10325, c10325, in10325_1, in10325_2, pp104[106]);
    wire[0:0] s10326, in10326_1, in10326_2;
    wire c10326;
    assign in10326_1 = {pp108[102]};
    assign in10326_2 = {pp109[101]};
    Full_Adder FA_10326(s10326, c10326, in10326_1, in10326_2, pp107[103]);
    wire[0:0] s10327, in10327_1, in10327_2;
    wire c10327;
    assign in10327_1 = {pp111[99]};
    assign in10327_2 = {pp112[98]};
    Full_Adder FA_10327(s10327, c10327, in10327_1, in10327_2, pp110[100]);
    wire[0:0] s10328, in10328_1, in10328_2;
    wire c10328;
    assign in10328_1 = {pp114[96]};
    assign in10328_2 = {pp115[95]};
    Full_Adder FA_10328(s10328, c10328, in10328_1, in10328_2, pp113[97]);
    wire[0:0] s10329, in10329_1, in10329_2;
    wire c10329;
    assign in10329_1 = {pp117[93]};
    assign in10329_2 = {pp118[92]};
    Full_Adder FA_10329(s10329, c10329, in10329_1, in10329_2, pp116[94]);
    wire[0:0] s10330, in10330_1, in10330_2;
    wire c10330;
    assign in10330_1 = {pp120[90]};
    assign in10330_2 = {pp121[89]};
    Full_Adder FA_10330(s10330, c10330, in10330_1, in10330_2, pp119[91]);
    wire[0:0] s10331, in10331_1, in10331_2;
    wire c10331;
    assign in10331_1 = {pp123[87]};
    assign in10331_2 = {pp124[86]};
    Full_Adder FA_10331(s10331, c10331, in10331_1, in10331_2, pp122[88]);
    wire[0:0] s10332, in10332_1, in10332_2;
    wire c10332;
    assign in10332_1 = {pp126[84]};
    assign in10332_2 = {pp127[83]};
    Full_Adder FA_10332(s10332, c10332, in10332_1, in10332_2, pp125[85]);
    wire[0:0] s10333, in10333_1, in10333_2;
    wire c10333;
    assign in10333_1 = {c7976};
    assign in10333_2 = {c7977};
    Full_Adder FA_10333(s10333, c10333, in10333_1, in10333_2, c7975);
    wire[0:0] s10334, in10334_1, in10334_2;
    wire c10334;
    assign in10334_1 = {c7979};
    assign in10334_2 = {c7980};
    Full_Adder FA_10334(s10334, c10334, in10334_1, in10334_2, c7978);
    wire[0:0] s10335, in10335_1, in10335_2;
    wire c10335;
    assign in10335_1 = {c7982};
    assign in10335_2 = {s7983[0]};
    Full_Adder FA_10335(s10335, c10335, in10335_1, in10335_2, c7981);
    wire[0:0] s10336, in10336_1, in10336_2;
    wire c10336;
    assign in10336_1 = {s7985[0]};
    assign in10336_2 = {s7986[0]};
    Full_Adder FA_10336(s10336, c10336, in10336_1, in10336_2, s7984[0]);
    wire[0:0] s10337, in10337_1, in10337_2;
    wire c10337;
    assign in10337_1 = {s7988[0]};
    assign in10337_2 = {s7989[0]};
    Full_Adder FA_10337(s10337, c10337, in10337_1, in10337_2, s7987[0]);
    wire[0:0] s10338, in10338_1, in10338_2;
    wire c10338;
    assign in10338_1 = {pp103[108]};
    assign in10338_2 = {pp104[107]};
    Full_Adder FA_10338(s10338, c10338, in10338_1, in10338_2, pp102[109]);
    wire[0:0] s10339, in10339_1, in10339_2;
    wire c10339;
    assign in10339_1 = {pp106[105]};
    assign in10339_2 = {pp107[104]};
    Full_Adder FA_10339(s10339, c10339, in10339_1, in10339_2, pp105[106]);
    wire[0:0] s10340, in10340_1, in10340_2;
    wire c10340;
    assign in10340_1 = {pp109[102]};
    assign in10340_2 = {pp110[101]};
    Full_Adder FA_10340(s10340, c10340, in10340_1, in10340_2, pp108[103]);
    wire[0:0] s10341, in10341_1, in10341_2;
    wire c10341;
    assign in10341_1 = {pp112[99]};
    assign in10341_2 = {pp113[98]};
    Full_Adder FA_10341(s10341, c10341, in10341_1, in10341_2, pp111[100]);
    wire[0:0] s10342, in10342_1, in10342_2;
    wire c10342;
    assign in10342_1 = {pp115[96]};
    assign in10342_2 = {pp116[95]};
    Full_Adder FA_10342(s10342, c10342, in10342_1, in10342_2, pp114[97]);
    wire[0:0] s10343, in10343_1, in10343_2;
    wire c10343;
    assign in10343_1 = {pp118[93]};
    assign in10343_2 = {pp119[92]};
    Full_Adder FA_10343(s10343, c10343, in10343_1, in10343_2, pp117[94]);
    wire[0:0] s10344, in10344_1, in10344_2;
    wire c10344;
    assign in10344_1 = {pp121[90]};
    assign in10344_2 = {pp122[89]};
    Full_Adder FA_10344(s10344, c10344, in10344_1, in10344_2, pp120[91]);
    wire[0:0] s10345, in10345_1, in10345_2;
    wire c10345;
    assign in10345_1 = {pp124[87]};
    assign in10345_2 = {pp125[86]};
    Full_Adder FA_10345(s10345, c10345, in10345_1, in10345_2, pp123[88]);
    wire[0:0] s10346, in10346_1, in10346_2;
    wire c10346;
    assign in10346_1 = {pp127[84]};
    assign in10346_2 = {c7983};
    Full_Adder FA_10346(s10346, c10346, in10346_1, in10346_2, pp126[85]);
    wire[0:0] s10347, in10347_1, in10347_2;
    wire c10347;
    assign in10347_1 = {c7985};
    assign in10347_2 = {c7986};
    Full_Adder FA_10347(s10347, c10347, in10347_1, in10347_2, c7984);
    wire[0:0] s10348, in10348_1, in10348_2;
    wire c10348;
    assign in10348_1 = {c7988};
    assign in10348_2 = {c7989};
    Full_Adder FA_10348(s10348, c10348, in10348_1, in10348_2, c7987);
    wire[0:0] s10349, in10349_1, in10349_2;
    wire c10349;
    assign in10349_1 = {s7991[0]};
    assign in10349_2 = {s7992[0]};
    Full_Adder FA_10349(s10349, c10349, in10349_1, in10349_2, s7990[0]);
    wire[0:0] s10350, in10350_1, in10350_2;
    wire c10350;
    assign in10350_1 = {s7994[0]};
    assign in10350_2 = {s7995[0]};
    Full_Adder FA_10350(s10350, c10350, in10350_1, in10350_2, s7993[0]);
    wire[0:0] s10351, in10351_1, in10351_2;
    wire c10351;
    assign in10351_1 = {pp101[111]};
    assign in10351_2 = {pp102[110]};
    Full_Adder FA_10351(s10351, c10351, in10351_1, in10351_2, pp100[112]);
    wire[0:0] s10352, in10352_1, in10352_2;
    wire c10352;
    assign in10352_1 = {pp104[108]};
    assign in10352_2 = {pp105[107]};
    Full_Adder FA_10352(s10352, c10352, in10352_1, in10352_2, pp103[109]);
    wire[0:0] s10353, in10353_1, in10353_2;
    wire c10353;
    assign in10353_1 = {pp107[105]};
    assign in10353_2 = {pp108[104]};
    Full_Adder FA_10353(s10353, c10353, in10353_1, in10353_2, pp106[106]);
    wire[0:0] s10354, in10354_1, in10354_2;
    wire c10354;
    assign in10354_1 = {pp110[102]};
    assign in10354_2 = {pp111[101]};
    Full_Adder FA_10354(s10354, c10354, in10354_1, in10354_2, pp109[103]);
    wire[0:0] s10355, in10355_1, in10355_2;
    wire c10355;
    assign in10355_1 = {pp113[99]};
    assign in10355_2 = {pp114[98]};
    Full_Adder FA_10355(s10355, c10355, in10355_1, in10355_2, pp112[100]);
    wire[0:0] s10356, in10356_1, in10356_2;
    wire c10356;
    assign in10356_1 = {pp116[96]};
    assign in10356_2 = {pp117[95]};
    Full_Adder FA_10356(s10356, c10356, in10356_1, in10356_2, pp115[97]);
    wire[0:0] s10357, in10357_1, in10357_2;
    wire c10357;
    assign in10357_1 = {pp119[93]};
    assign in10357_2 = {pp120[92]};
    Full_Adder FA_10357(s10357, c10357, in10357_1, in10357_2, pp118[94]);
    wire[0:0] s10358, in10358_1, in10358_2;
    wire c10358;
    assign in10358_1 = {pp122[90]};
    assign in10358_2 = {pp123[89]};
    Full_Adder FA_10358(s10358, c10358, in10358_1, in10358_2, pp121[91]);
    wire[0:0] s10359, in10359_1, in10359_2;
    wire c10359;
    assign in10359_1 = {pp125[87]};
    assign in10359_2 = {pp126[86]};
    Full_Adder FA_10359(s10359, c10359, in10359_1, in10359_2, pp124[88]);
    wire[0:0] s10360, in10360_1, in10360_2;
    wire c10360;
    assign in10360_1 = {c7990};
    assign in10360_2 = {c7991};
    Full_Adder FA_10360(s10360, c10360, in10360_1, in10360_2, pp127[85]);
    wire[0:0] s10361, in10361_1, in10361_2;
    wire c10361;
    assign in10361_1 = {c7993};
    assign in10361_2 = {c7994};
    Full_Adder FA_10361(s10361, c10361, in10361_1, in10361_2, c7992);
    wire[0:0] s10362, in10362_1, in10362_2;
    wire c10362;
    assign in10362_1 = {s7996[0]};
    assign in10362_2 = {s7997[0]};
    Full_Adder FA_10362(s10362, c10362, in10362_1, in10362_2, c7995);
    wire[0:0] s10363, in10363_1, in10363_2;
    wire c10363;
    assign in10363_1 = {s7999[0]};
    assign in10363_2 = {s8000[0]};
    Full_Adder FA_10363(s10363, c10363, in10363_1, in10363_2, s7998[0]);
    wire[0:0] s10364, in10364_1, in10364_2;
    wire c10364;
    assign in10364_1 = {pp99[114]};
    assign in10364_2 = {pp100[113]};
    Full_Adder FA_10364(s10364, c10364, in10364_1, in10364_2, pp98[115]);
    wire[0:0] s10365, in10365_1, in10365_2;
    wire c10365;
    assign in10365_1 = {pp102[111]};
    assign in10365_2 = {pp103[110]};
    Full_Adder FA_10365(s10365, c10365, in10365_1, in10365_2, pp101[112]);
    wire[0:0] s10366, in10366_1, in10366_2;
    wire c10366;
    assign in10366_1 = {pp105[108]};
    assign in10366_2 = {pp106[107]};
    Full_Adder FA_10366(s10366, c10366, in10366_1, in10366_2, pp104[109]);
    wire[0:0] s10367, in10367_1, in10367_2;
    wire c10367;
    assign in10367_1 = {pp108[105]};
    assign in10367_2 = {pp109[104]};
    Full_Adder FA_10367(s10367, c10367, in10367_1, in10367_2, pp107[106]);
    wire[0:0] s10368, in10368_1, in10368_2;
    wire c10368;
    assign in10368_1 = {pp111[102]};
    assign in10368_2 = {pp112[101]};
    Full_Adder FA_10368(s10368, c10368, in10368_1, in10368_2, pp110[103]);
    wire[0:0] s10369, in10369_1, in10369_2;
    wire c10369;
    assign in10369_1 = {pp114[99]};
    assign in10369_2 = {pp115[98]};
    Full_Adder FA_10369(s10369, c10369, in10369_1, in10369_2, pp113[100]);
    wire[0:0] s10370, in10370_1, in10370_2;
    wire c10370;
    assign in10370_1 = {pp117[96]};
    assign in10370_2 = {pp118[95]};
    Full_Adder FA_10370(s10370, c10370, in10370_1, in10370_2, pp116[97]);
    wire[0:0] s10371, in10371_1, in10371_2;
    wire c10371;
    assign in10371_1 = {pp120[93]};
    assign in10371_2 = {pp121[92]};
    Full_Adder FA_10371(s10371, c10371, in10371_1, in10371_2, pp119[94]);
    wire[0:0] s10372, in10372_1, in10372_2;
    wire c10372;
    assign in10372_1 = {pp123[90]};
    assign in10372_2 = {pp124[89]};
    Full_Adder FA_10372(s10372, c10372, in10372_1, in10372_2, pp122[91]);
    wire[0:0] s10373, in10373_1, in10373_2;
    wire c10373;
    assign in10373_1 = {pp126[87]};
    assign in10373_2 = {pp127[86]};
    Full_Adder FA_10373(s10373, c10373, in10373_1, in10373_2, pp125[88]);
    wire[0:0] s10374, in10374_1, in10374_2;
    wire c10374;
    assign in10374_1 = {c7997};
    assign in10374_2 = {c7998};
    Full_Adder FA_10374(s10374, c10374, in10374_1, in10374_2, c7996);
    wire[0:0] s10375, in10375_1, in10375_2;
    wire c10375;
    assign in10375_1 = {c8000};
    assign in10375_2 = {s8001[0]};
    Full_Adder FA_10375(s10375, c10375, in10375_1, in10375_2, c7999);
    wire[0:0] s10376, in10376_1, in10376_2;
    wire c10376;
    assign in10376_1 = {s8003[0]};
    assign in10376_2 = {s8004[0]};
    Full_Adder FA_10376(s10376, c10376, in10376_1, in10376_2, s8002[0]);
    wire[0:0] s10377, in10377_1, in10377_2;
    wire c10377;
    assign in10377_1 = {pp97[117]};
    assign in10377_2 = {pp98[116]};
    Full_Adder FA_10377(s10377, c10377, in10377_1, in10377_2, pp96[118]);
    wire[0:0] s10378, in10378_1, in10378_2;
    wire c10378;
    assign in10378_1 = {pp100[114]};
    assign in10378_2 = {pp101[113]};
    Full_Adder FA_10378(s10378, c10378, in10378_1, in10378_2, pp99[115]);
    wire[0:0] s10379, in10379_1, in10379_2;
    wire c10379;
    assign in10379_1 = {pp103[111]};
    assign in10379_2 = {pp104[110]};
    Full_Adder FA_10379(s10379, c10379, in10379_1, in10379_2, pp102[112]);
    wire[0:0] s10380, in10380_1, in10380_2;
    wire c10380;
    assign in10380_1 = {pp106[108]};
    assign in10380_2 = {pp107[107]};
    Full_Adder FA_10380(s10380, c10380, in10380_1, in10380_2, pp105[109]);
    wire[0:0] s10381, in10381_1, in10381_2;
    wire c10381;
    assign in10381_1 = {pp109[105]};
    assign in10381_2 = {pp110[104]};
    Full_Adder FA_10381(s10381, c10381, in10381_1, in10381_2, pp108[106]);
    wire[0:0] s10382, in10382_1, in10382_2;
    wire c10382;
    assign in10382_1 = {pp112[102]};
    assign in10382_2 = {pp113[101]};
    Full_Adder FA_10382(s10382, c10382, in10382_1, in10382_2, pp111[103]);
    wire[0:0] s10383, in10383_1, in10383_2;
    wire c10383;
    assign in10383_1 = {pp115[99]};
    assign in10383_2 = {pp116[98]};
    Full_Adder FA_10383(s10383, c10383, in10383_1, in10383_2, pp114[100]);
    wire[0:0] s10384, in10384_1, in10384_2;
    wire c10384;
    assign in10384_1 = {pp118[96]};
    assign in10384_2 = {pp119[95]};
    Full_Adder FA_10384(s10384, c10384, in10384_1, in10384_2, pp117[97]);
    wire[0:0] s10385, in10385_1, in10385_2;
    wire c10385;
    assign in10385_1 = {pp121[93]};
    assign in10385_2 = {pp122[92]};
    Full_Adder FA_10385(s10385, c10385, in10385_1, in10385_2, pp120[94]);
    wire[0:0] s10386, in10386_1, in10386_2;
    wire c10386;
    assign in10386_1 = {pp124[90]};
    assign in10386_2 = {pp125[89]};
    Full_Adder FA_10386(s10386, c10386, in10386_1, in10386_2, pp123[91]);
    wire[0:0] s10387, in10387_1, in10387_2;
    wire c10387;
    assign in10387_1 = {pp127[87]};
    assign in10387_2 = {c8001};
    Full_Adder FA_10387(s10387, c10387, in10387_1, in10387_2, pp126[88]);
    wire[0:0] s10388, in10388_1, in10388_2;
    wire c10388;
    assign in10388_1 = {c8003};
    assign in10388_2 = {c8004};
    Full_Adder FA_10388(s10388, c10388, in10388_1, in10388_2, c8002);
    wire[0:0] s10389, in10389_1, in10389_2;
    wire c10389;
    assign in10389_1 = {s8006[0]};
    assign in10389_2 = {s8007[0]};
    Full_Adder FA_10389(s10389, c10389, in10389_1, in10389_2, s8005[0]);
    wire[0:0] s10390, in10390_1, in10390_2;
    wire c10390;
    assign in10390_1 = {pp95[120]};
    assign in10390_2 = {pp96[119]};
    Full_Adder FA_10390(s10390, c10390, in10390_1, in10390_2, pp94[121]);
    wire[0:0] s10391, in10391_1, in10391_2;
    wire c10391;
    assign in10391_1 = {pp98[117]};
    assign in10391_2 = {pp99[116]};
    Full_Adder FA_10391(s10391, c10391, in10391_1, in10391_2, pp97[118]);
    wire[0:0] s10392, in10392_1, in10392_2;
    wire c10392;
    assign in10392_1 = {pp101[114]};
    assign in10392_2 = {pp102[113]};
    Full_Adder FA_10392(s10392, c10392, in10392_1, in10392_2, pp100[115]);
    wire[0:0] s10393, in10393_1, in10393_2;
    wire c10393;
    assign in10393_1 = {pp104[111]};
    assign in10393_2 = {pp105[110]};
    Full_Adder FA_10393(s10393, c10393, in10393_1, in10393_2, pp103[112]);
    wire[0:0] s10394, in10394_1, in10394_2;
    wire c10394;
    assign in10394_1 = {pp107[108]};
    assign in10394_2 = {pp108[107]};
    Full_Adder FA_10394(s10394, c10394, in10394_1, in10394_2, pp106[109]);
    wire[0:0] s10395, in10395_1, in10395_2;
    wire c10395;
    assign in10395_1 = {pp110[105]};
    assign in10395_2 = {pp111[104]};
    Full_Adder FA_10395(s10395, c10395, in10395_1, in10395_2, pp109[106]);
    wire[0:0] s10396, in10396_1, in10396_2;
    wire c10396;
    assign in10396_1 = {pp113[102]};
    assign in10396_2 = {pp114[101]};
    Full_Adder FA_10396(s10396, c10396, in10396_1, in10396_2, pp112[103]);
    wire[0:0] s10397, in10397_1, in10397_2;
    wire c10397;
    assign in10397_1 = {pp116[99]};
    assign in10397_2 = {pp117[98]};
    Full_Adder FA_10397(s10397, c10397, in10397_1, in10397_2, pp115[100]);
    wire[0:0] s10398, in10398_1, in10398_2;
    wire c10398;
    assign in10398_1 = {pp119[96]};
    assign in10398_2 = {pp120[95]};
    Full_Adder FA_10398(s10398, c10398, in10398_1, in10398_2, pp118[97]);
    wire[0:0] s10399, in10399_1, in10399_2;
    wire c10399;
    assign in10399_1 = {pp122[93]};
    assign in10399_2 = {pp123[92]};
    Full_Adder FA_10399(s10399, c10399, in10399_1, in10399_2, pp121[94]);
    wire[0:0] s10400, in10400_1, in10400_2;
    wire c10400;
    assign in10400_1 = {pp125[90]};
    assign in10400_2 = {pp126[89]};
    Full_Adder FA_10400(s10400, c10400, in10400_1, in10400_2, pp124[91]);
    wire[0:0] s10401, in10401_1, in10401_2;
    wire c10401;
    assign in10401_1 = {c8005};
    assign in10401_2 = {c8006};
    Full_Adder FA_10401(s10401, c10401, in10401_1, in10401_2, pp127[88]);
    wire[0:0] s10402, in10402_1, in10402_2;
    wire c10402;
    assign in10402_1 = {s8008[0]};
    assign in10402_2 = {s8009[0]};
    Full_Adder FA_10402(s10402, c10402, in10402_1, in10402_2, c8007);
    wire[0:0] s10403, in10403_1, in10403_2;
    wire c10403;
    assign in10403_1 = {pp93[123]};
    assign in10403_2 = {pp94[122]};
    Full_Adder FA_10403(s10403, c10403, in10403_1, in10403_2, pp92[124]);
    wire[0:0] s10404, in10404_1, in10404_2;
    wire c10404;
    assign in10404_1 = {pp96[120]};
    assign in10404_2 = {pp97[119]};
    Full_Adder FA_10404(s10404, c10404, in10404_1, in10404_2, pp95[121]);
    wire[0:0] s10405, in10405_1, in10405_2;
    wire c10405;
    assign in10405_1 = {pp99[117]};
    assign in10405_2 = {pp100[116]};
    Full_Adder FA_10405(s10405, c10405, in10405_1, in10405_2, pp98[118]);
    wire[0:0] s10406, in10406_1, in10406_2;
    wire c10406;
    assign in10406_1 = {pp102[114]};
    assign in10406_2 = {pp103[113]};
    Full_Adder FA_10406(s10406, c10406, in10406_1, in10406_2, pp101[115]);
    wire[0:0] s10407, in10407_1, in10407_2;
    wire c10407;
    assign in10407_1 = {pp105[111]};
    assign in10407_2 = {pp106[110]};
    Full_Adder FA_10407(s10407, c10407, in10407_1, in10407_2, pp104[112]);
    wire[0:0] s10408, in10408_1, in10408_2;
    wire c10408;
    assign in10408_1 = {pp108[108]};
    assign in10408_2 = {pp109[107]};
    Full_Adder FA_10408(s10408, c10408, in10408_1, in10408_2, pp107[109]);
    wire[0:0] s10409, in10409_1, in10409_2;
    wire c10409;
    assign in10409_1 = {pp111[105]};
    assign in10409_2 = {pp112[104]};
    Full_Adder FA_10409(s10409, c10409, in10409_1, in10409_2, pp110[106]);
    wire[0:0] s10410, in10410_1, in10410_2;
    wire c10410;
    assign in10410_1 = {pp114[102]};
    assign in10410_2 = {pp115[101]};
    Full_Adder FA_10410(s10410, c10410, in10410_1, in10410_2, pp113[103]);
    wire[0:0] s10411, in10411_1, in10411_2;
    wire c10411;
    assign in10411_1 = {pp117[99]};
    assign in10411_2 = {pp118[98]};
    Full_Adder FA_10411(s10411, c10411, in10411_1, in10411_2, pp116[100]);
    wire[0:0] s10412, in10412_1, in10412_2;
    wire c10412;
    assign in10412_1 = {pp120[96]};
    assign in10412_2 = {pp121[95]};
    Full_Adder FA_10412(s10412, c10412, in10412_1, in10412_2, pp119[97]);
    wire[0:0] s10413, in10413_1, in10413_2;
    wire c10413;
    assign in10413_1 = {pp123[93]};
    assign in10413_2 = {pp124[92]};
    Full_Adder FA_10413(s10413, c10413, in10413_1, in10413_2, pp122[94]);
    wire[0:0] s10414, in10414_1, in10414_2;
    wire c10414;
    assign in10414_1 = {pp126[90]};
    assign in10414_2 = {pp127[89]};
    Full_Adder FA_10414(s10414, c10414, in10414_1, in10414_2, pp125[91]);
    wire[0:0] s10415, in10415_1, in10415_2;
    wire c10415;
    assign in10415_1 = {c8009};
    assign in10415_2 = {s8010[0]};
    Full_Adder FA_10415(s10415, c10415, in10415_1, in10415_2, c8008);
    wire[0:0] s10416, in10416_1, in10416_2;
    wire c10416;
    assign in10416_1 = {pp91[126]};
    assign in10416_2 = {pp92[125]};
    Full_Adder FA_10416(s10416, c10416, in10416_1, in10416_2, pp90[127]);
    wire[0:0] s10417, in10417_1, in10417_2;
    wire c10417;
    assign in10417_1 = {pp94[123]};
    assign in10417_2 = {pp95[122]};
    Full_Adder FA_10417(s10417, c10417, in10417_1, in10417_2, pp93[124]);
    wire[0:0] s10418, in10418_1, in10418_2;
    wire c10418;
    assign in10418_1 = {pp97[120]};
    assign in10418_2 = {pp98[119]};
    Full_Adder FA_10418(s10418, c10418, in10418_1, in10418_2, pp96[121]);
    wire[0:0] s10419, in10419_1, in10419_2;
    wire c10419;
    assign in10419_1 = {pp100[117]};
    assign in10419_2 = {pp101[116]};
    Full_Adder FA_10419(s10419, c10419, in10419_1, in10419_2, pp99[118]);
    wire[0:0] s10420, in10420_1, in10420_2;
    wire c10420;
    assign in10420_1 = {pp103[114]};
    assign in10420_2 = {pp104[113]};
    Full_Adder FA_10420(s10420, c10420, in10420_1, in10420_2, pp102[115]);
    wire[0:0] s10421, in10421_1, in10421_2;
    wire c10421;
    assign in10421_1 = {pp106[111]};
    assign in10421_2 = {pp107[110]};
    Full_Adder FA_10421(s10421, c10421, in10421_1, in10421_2, pp105[112]);
    wire[0:0] s10422, in10422_1, in10422_2;
    wire c10422;
    assign in10422_1 = {pp109[108]};
    assign in10422_2 = {pp110[107]};
    Full_Adder FA_10422(s10422, c10422, in10422_1, in10422_2, pp108[109]);
    wire[0:0] s10423, in10423_1, in10423_2;
    wire c10423;
    assign in10423_1 = {pp112[105]};
    assign in10423_2 = {pp113[104]};
    Full_Adder FA_10423(s10423, c10423, in10423_1, in10423_2, pp111[106]);
    wire[0:0] s10424, in10424_1, in10424_2;
    wire c10424;
    assign in10424_1 = {pp115[102]};
    assign in10424_2 = {pp116[101]};
    Full_Adder FA_10424(s10424, c10424, in10424_1, in10424_2, pp114[103]);
    wire[0:0] s10425, in10425_1, in10425_2;
    wire c10425;
    assign in10425_1 = {pp118[99]};
    assign in10425_2 = {pp119[98]};
    Full_Adder FA_10425(s10425, c10425, in10425_1, in10425_2, pp117[100]);
    wire[0:0] s10426, in10426_1, in10426_2;
    wire c10426;
    assign in10426_1 = {pp121[96]};
    assign in10426_2 = {pp122[95]};
    Full_Adder FA_10426(s10426, c10426, in10426_1, in10426_2, pp120[97]);
    wire[0:0] s10427, in10427_1, in10427_2;
    wire c10427;
    assign in10427_1 = {pp124[93]};
    assign in10427_2 = {pp125[92]};
    Full_Adder FA_10427(s10427, c10427, in10427_1, in10427_2, pp123[94]);
    wire[0:0] s10428, in10428_1, in10428_2;
    wire c10428;
    assign in10428_1 = {pp127[90]};
    assign in10428_2 = {c8010};
    Full_Adder FA_10428(s10428, c10428, in10428_1, in10428_2, pp126[91]);
    wire[0:0] s10429, in10429_1, in10429_2;
    wire c10429;
    assign in10429_1 = {pp92[126]};
    assign in10429_2 = {pp93[125]};
    Full_Adder FA_10429(s10429, c10429, in10429_1, in10429_2, pp91[127]);
    wire[0:0] s10430, in10430_1, in10430_2;
    wire c10430;
    assign in10430_1 = {pp95[123]};
    assign in10430_2 = {pp96[122]};
    Full_Adder FA_10430(s10430, c10430, in10430_1, in10430_2, pp94[124]);
    wire[0:0] s10431, in10431_1, in10431_2;
    wire c10431;
    assign in10431_1 = {pp98[120]};
    assign in10431_2 = {pp99[119]};
    Full_Adder FA_10431(s10431, c10431, in10431_1, in10431_2, pp97[121]);
    wire[0:0] s10432, in10432_1, in10432_2;
    wire c10432;
    assign in10432_1 = {pp101[117]};
    assign in10432_2 = {pp102[116]};
    Full_Adder FA_10432(s10432, c10432, in10432_1, in10432_2, pp100[118]);
    wire[0:0] s10433, in10433_1, in10433_2;
    wire c10433;
    assign in10433_1 = {pp104[114]};
    assign in10433_2 = {pp105[113]};
    Full_Adder FA_10433(s10433, c10433, in10433_1, in10433_2, pp103[115]);
    wire[0:0] s10434, in10434_1, in10434_2;
    wire c10434;
    assign in10434_1 = {pp107[111]};
    assign in10434_2 = {pp108[110]};
    Full_Adder FA_10434(s10434, c10434, in10434_1, in10434_2, pp106[112]);
    wire[0:0] s10435, in10435_1, in10435_2;
    wire c10435;
    assign in10435_1 = {pp110[108]};
    assign in10435_2 = {pp111[107]};
    Full_Adder FA_10435(s10435, c10435, in10435_1, in10435_2, pp109[109]);
    wire[0:0] s10436, in10436_1, in10436_2;
    wire c10436;
    assign in10436_1 = {pp113[105]};
    assign in10436_2 = {pp114[104]};
    Full_Adder FA_10436(s10436, c10436, in10436_1, in10436_2, pp112[106]);
    wire[0:0] s10437, in10437_1, in10437_2;
    wire c10437;
    assign in10437_1 = {pp116[102]};
    assign in10437_2 = {pp117[101]};
    Full_Adder FA_10437(s10437, c10437, in10437_1, in10437_2, pp115[103]);
    wire[0:0] s10438, in10438_1, in10438_2;
    wire c10438;
    assign in10438_1 = {pp119[99]};
    assign in10438_2 = {pp120[98]};
    Full_Adder FA_10438(s10438, c10438, in10438_1, in10438_2, pp118[100]);
    wire[0:0] s10439, in10439_1, in10439_2;
    wire c10439;
    assign in10439_1 = {pp122[96]};
    assign in10439_2 = {pp123[95]};
    Full_Adder FA_10439(s10439, c10439, in10439_1, in10439_2, pp121[97]);
    wire[0:0] s10440, in10440_1, in10440_2;
    wire c10440;
    assign in10440_1 = {pp125[93]};
    assign in10440_2 = {pp126[92]};
    Full_Adder FA_10440(s10440, c10440, in10440_1, in10440_2, pp124[94]);
    wire[0:0] s10441, in10441_1, in10441_2;
    wire c10441;
    assign in10441_1 = {pp93[126]};
    assign in10441_2 = {pp94[125]};
    Full_Adder FA_10441(s10441, c10441, in10441_1, in10441_2, pp92[127]);
    wire[0:0] s10442, in10442_1, in10442_2;
    wire c10442;
    assign in10442_1 = {pp96[123]};
    assign in10442_2 = {pp97[122]};
    Full_Adder FA_10442(s10442, c10442, in10442_1, in10442_2, pp95[124]);
    wire[0:0] s10443, in10443_1, in10443_2;
    wire c10443;
    assign in10443_1 = {pp99[120]};
    assign in10443_2 = {pp100[119]};
    Full_Adder FA_10443(s10443, c10443, in10443_1, in10443_2, pp98[121]);
    wire[0:0] s10444, in10444_1, in10444_2;
    wire c10444;
    assign in10444_1 = {pp102[117]};
    assign in10444_2 = {pp103[116]};
    Full_Adder FA_10444(s10444, c10444, in10444_1, in10444_2, pp101[118]);
    wire[0:0] s10445, in10445_1, in10445_2;
    wire c10445;
    assign in10445_1 = {pp105[114]};
    assign in10445_2 = {pp106[113]};
    Full_Adder FA_10445(s10445, c10445, in10445_1, in10445_2, pp104[115]);
    wire[0:0] s10446, in10446_1, in10446_2;
    wire c10446;
    assign in10446_1 = {pp108[111]};
    assign in10446_2 = {pp109[110]};
    Full_Adder FA_10446(s10446, c10446, in10446_1, in10446_2, pp107[112]);
    wire[0:0] s10447, in10447_1, in10447_2;
    wire c10447;
    assign in10447_1 = {pp111[108]};
    assign in10447_2 = {pp112[107]};
    Full_Adder FA_10447(s10447, c10447, in10447_1, in10447_2, pp110[109]);
    wire[0:0] s10448, in10448_1, in10448_2;
    wire c10448;
    assign in10448_1 = {pp114[105]};
    assign in10448_2 = {pp115[104]};
    Full_Adder FA_10448(s10448, c10448, in10448_1, in10448_2, pp113[106]);
    wire[0:0] s10449, in10449_1, in10449_2;
    wire c10449;
    assign in10449_1 = {pp117[102]};
    assign in10449_2 = {pp118[101]};
    Full_Adder FA_10449(s10449, c10449, in10449_1, in10449_2, pp116[103]);
    wire[0:0] s10450, in10450_1, in10450_2;
    wire c10450;
    assign in10450_1 = {pp120[99]};
    assign in10450_2 = {pp121[98]};
    Full_Adder FA_10450(s10450, c10450, in10450_1, in10450_2, pp119[100]);
    wire[0:0] s10451, in10451_1, in10451_2;
    wire c10451;
    assign in10451_1 = {pp123[96]};
    assign in10451_2 = {pp124[95]};
    Full_Adder FA_10451(s10451, c10451, in10451_1, in10451_2, pp122[97]);
    wire[0:0] s10452, in10452_1, in10452_2;
    wire c10452;
    assign in10452_1 = {pp94[126]};
    assign in10452_2 = {pp95[125]};
    Full_Adder FA_10452(s10452, c10452, in10452_1, in10452_2, pp93[127]);
    wire[0:0] s10453, in10453_1, in10453_2;
    wire c10453;
    assign in10453_1 = {pp97[123]};
    assign in10453_2 = {pp98[122]};
    Full_Adder FA_10453(s10453, c10453, in10453_1, in10453_2, pp96[124]);
    wire[0:0] s10454, in10454_1, in10454_2;
    wire c10454;
    assign in10454_1 = {pp100[120]};
    assign in10454_2 = {pp101[119]};
    Full_Adder FA_10454(s10454, c10454, in10454_1, in10454_2, pp99[121]);
    wire[0:0] s10455, in10455_1, in10455_2;
    wire c10455;
    assign in10455_1 = {pp103[117]};
    assign in10455_2 = {pp104[116]};
    Full_Adder FA_10455(s10455, c10455, in10455_1, in10455_2, pp102[118]);
    wire[0:0] s10456, in10456_1, in10456_2;
    wire c10456;
    assign in10456_1 = {pp106[114]};
    assign in10456_2 = {pp107[113]};
    Full_Adder FA_10456(s10456, c10456, in10456_1, in10456_2, pp105[115]);
    wire[0:0] s10457, in10457_1, in10457_2;
    wire c10457;
    assign in10457_1 = {pp109[111]};
    assign in10457_2 = {pp110[110]};
    Full_Adder FA_10457(s10457, c10457, in10457_1, in10457_2, pp108[112]);
    wire[0:0] s10458, in10458_1, in10458_2;
    wire c10458;
    assign in10458_1 = {pp112[108]};
    assign in10458_2 = {pp113[107]};
    Full_Adder FA_10458(s10458, c10458, in10458_1, in10458_2, pp111[109]);
    wire[0:0] s10459, in10459_1, in10459_2;
    wire c10459;
    assign in10459_1 = {pp115[105]};
    assign in10459_2 = {pp116[104]};
    Full_Adder FA_10459(s10459, c10459, in10459_1, in10459_2, pp114[106]);
    wire[0:0] s10460, in10460_1, in10460_2;
    wire c10460;
    assign in10460_1 = {pp118[102]};
    assign in10460_2 = {pp119[101]};
    Full_Adder FA_10460(s10460, c10460, in10460_1, in10460_2, pp117[103]);
    wire[0:0] s10461, in10461_1, in10461_2;
    wire c10461;
    assign in10461_1 = {pp121[99]};
    assign in10461_2 = {pp122[98]};
    Full_Adder FA_10461(s10461, c10461, in10461_1, in10461_2, pp120[100]);
    wire[0:0] s10462, in10462_1, in10462_2;
    wire c10462;
    assign in10462_1 = {pp95[126]};
    assign in10462_2 = {pp96[125]};
    Full_Adder FA_10462(s10462, c10462, in10462_1, in10462_2, pp94[127]);
    wire[0:0] s10463, in10463_1, in10463_2;
    wire c10463;
    assign in10463_1 = {pp98[123]};
    assign in10463_2 = {pp99[122]};
    Full_Adder FA_10463(s10463, c10463, in10463_1, in10463_2, pp97[124]);
    wire[0:0] s10464, in10464_1, in10464_2;
    wire c10464;
    assign in10464_1 = {pp101[120]};
    assign in10464_2 = {pp102[119]};
    Full_Adder FA_10464(s10464, c10464, in10464_1, in10464_2, pp100[121]);
    wire[0:0] s10465, in10465_1, in10465_2;
    wire c10465;
    assign in10465_1 = {pp104[117]};
    assign in10465_2 = {pp105[116]};
    Full_Adder FA_10465(s10465, c10465, in10465_1, in10465_2, pp103[118]);
    wire[0:0] s10466, in10466_1, in10466_2;
    wire c10466;
    assign in10466_1 = {pp107[114]};
    assign in10466_2 = {pp108[113]};
    Full_Adder FA_10466(s10466, c10466, in10466_1, in10466_2, pp106[115]);
    wire[0:0] s10467, in10467_1, in10467_2;
    wire c10467;
    assign in10467_1 = {pp110[111]};
    assign in10467_2 = {pp111[110]};
    Full_Adder FA_10467(s10467, c10467, in10467_1, in10467_2, pp109[112]);
    wire[0:0] s10468, in10468_1, in10468_2;
    wire c10468;
    assign in10468_1 = {pp113[108]};
    assign in10468_2 = {pp114[107]};
    Full_Adder FA_10468(s10468, c10468, in10468_1, in10468_2, pp112[109]);
    wire[0:0] s10469, in10469_1, in10469_2;
    wire c10469;
    assign in10469_1 = {pp116[105]};
    assign in10469_2 = {pp117[104]};
    Full_Adder FA_10469(s10469, c10469, in10469_1, in10469_2, pp115[106]);
    wire[0:0] s10470, in10470_1, in10470_2;
    wire c10470;
    assign in10470_1 = {pp119[102]};
    assign in10470_2 = {pp120[101]};
    Full_Adder FA_10470(s10470, c10470, in10470_1, in10470_2, pp118[103]);
    wire[0:0] s10471, in10471_1, in10471_2;
    wire c10471;
    assign in10471_1 = {pp96[126]};
    assign in10471_2 = {pp97[125]};
    Full_Adder FA_10471(s10471, c10471, in10471_1, in10471_2, pp95[127]);
    wire[0:0] s10472, in10472_1, in10472_2;
    wire c10472;
    assign in10472_1 = {pp99[123]};
    assign in10472_2 = {pp100[122]};
    Full_Adder FA_10472(s10472, c10472, in10472_1, in10472_2, pp98[124]);
    wire[0:0] s10473, in10473_1, in10473_2;
    wire c10473;
    assign in10473_1 = {pp102[120]};
    assign in10473_2 = {pp103[119]};
    Full_Adder FA_10473(s10473, c10473, in10473_1, in10473_2, pp101[121]);
    wire[0:0] s10474, in10474_1, in10474_2;
    wire c10474;
    assign in10474_1 = {pp105[117]};
    assign in10474_2 = {pp106[116]};
    Full_Adder FA_10474(s10474, c10474, in10474_1, in10474_2, pp104[118]);
    wire[0:0] s10475, in10475_1, in10475_2;
    wire c10475;
    assign in10475_1 = {pp108[114]};
    assign in10475_2 = {pp109[113]};
    Full_Adder FA_10475(s10475, c10475, in10475_1, in10475_2, pp107[115]);
    wire[0:0] s10476, in10476_1, in10476_2;
    wire c10476;
    assign in10476_1 = {pp111[111]};
    assign in10476_2 = {pp112[110]};
    Full_Adder FA_10476(s10476, c10476, in10476_1, in10476_2, pp110[112]);
    wire[0:0] s10477, in10477_1, in10477_2;
    wire c10477;
    assign in10477_1 = {pp114[108]};
    assign in10477_2 = {pp115[107]};
    Full_Adder FA_10477(s10477, c10477, in10477_1, in10477_2, pp113[109]);
    wire[0:0] s10478, in10478_1, in10478_2;
    wire c10478;
    assign in10478_1 = {pp117[105]};
    assign in10478_2 = {pp118[104]};
    Full_Adder FA_10478(s10478, c10478, in10478_1, in10478_2, pp116[106]);
    wire[0:0] s10479, in10479_1, in10479_2;
    wire c10479;
    assign in10479_1 = {pp97[126]};
    assign in10479_2 = {pp98[125]};
    Full_Adder FA_10479(s10479, c10479, in10479_1, in10479_2, pp96[127]);
    wire[0:0] s10480, in10480_1, in10480_2;
    wire c10480;
    assign in10480_1 = {pp100[123]};
    assign in10480_2 = {pp101[122]};
    Full_Adder FA_10480(s10480, c10480, in10480_1, in10480_2, pp99[124]);
    wire[0:0] s10481, in10481_1, in10481_2;
    wire c10481;
    assign in10481_1 = {pp103[120]};
    assign in10481_2 = {pp104[119]};
    Full_Adder FA_10481(s10481, c10481, in10481_1, in10481_2, pp102[121]);
    wire[0:0] s10482, in10482_1, in10482_2;
    wire c10482;
    assign in10482_1 = {pp106[117]};
    assign in10482_2 = {pp107[116]};
    Full_Adder FA_10482(s10482, c10482, in10482_1, in10482_2, pp105[118]);
    wire[0:0] s10483, in10483_1, in10483_2;
    wire c10483;
    assign in10483_1 = {pp109[114]};
    assign in10483_2 = {pp110[113]};
    Full_Adder FA_10483(s10483, c10483, in10483_1, in10483_2, pp108[115]);
    wire[0:0] s10484, in10484_1, in10484_2;
    wire c10484;
    assign in10484_1 = {pp112[111]};
    assign in10484_2 = {pp113[110]};
    Full_Adder FA_10484(s10484, c10484, in10484_1, in10484_2, pp111[112]);
    wire[0:0] s10485, in10485_1, in10485_2;
    wire c10485;
    assign in10485_1 = {pp115[108]};
    assign in10485_2 = {pp116[107]};
    Full_Adder FA_10485(s10485, c10485, in10485_1, in10485_2, pp114[109]);
    wire[0:0] s10486, in10486_1, in10486_2;
    wire c10486;
    assign in10486_1 = {pp98[126]};
    assign in10486_2 = {pp99[125]};
    Full_Adder FA_10486(s10486, c10486, in10486_1, in10486_2, pp97[127]);
    wire[0:0] s10487, in10487_1, in10487_2;
    wire c10487;
    assign in10487_1 = {pp101[123]};
    assign in10487_2 = {pp102[122]};
    Full_Adder FA_10487(s10487, c10487, in10487_1, in10487_2, pp100[124]);
    wire[0:0] s10488, in10488_1, in10488_2;
    wire c10488;
    assign in10488_1 = {pp104[120]};
    assign in10488_2 = {pp105[119]};
    Full_Adder FA_10488(s10488, c10488, in10488_1, in10488_2, pp103[121]);
    wire[0:0] s10489, in10489_1, in10489_2;
    wire c10489;
    assign in10489_1 = {pp107[117]};
    assign in10489_2 = {pp108[116]};
    Full_Adder FA_10489(s10489, c10489, in10489_1, in10489_2, pp106[118]);
    wire[0:0] s10490, in10490_1, in10490_2;
    wire c10490;
    assign in10490_1 = {pp110[114]};
    assign in10490_2 = {pp111[113]};
    Full_Adder FA_10490(s10490, c10490, in10490_1, in10490_2, pp109[115]);
    wire[0:0] s10491, in10491_1, in10491_2;
    wire c10491;
    assign in10491_1 = {pp113[111]};
    assign in10491_2 = {pp114[110]};
    Full_Adder FA_10491(s10491, c10491, in10491_1, in10491_2, pp112[112]);
    wire[0:0] s10492, in10492_1, in10492_2;
    wire c10492;
    assign in10492_1 = {pp99[126]};
    assign in10492_2 = {pp100[125]};
    Full_Adder FA_10492(s10492, c10492, in10492_1, in10492_2, pp98[127]);
    wire[0:0] s10493, in10493_1, in10493_2;
    wire c10493;
    assign in10493_1 = {pp102[123]};
    assign in10493_2 = {pp103[122]};
    Full_Adder FA_10493(s10493, c10493, in10493_1, in10493_2, pp101[124]);
    wire[0:0] s10494, in10494_1, in10494_2;
    wire c10494;
    assign in10494_1 = {pp105[120]};
    assign in10494_2 = {pp106[119]};
    Full_Adder FA_10494(s10494, c10494, in10494_1, in10494_2, pp104[121]);
    wire[0:0] s10495, in10495_1, in10495_2;
    wire c10495;
    assign in10495_1 = {pp108[117]};
    assign in10495_2 = {pp109[116]};
    Full_Adder FA_10495(s10495, c10495, in10495_1, in10495_2, pp107[118]);
    wire[0:0] s10496, in10496_1, in10496_2;
    wire c10496;
    assign in10496_1 = {pp111[114]};
    assign in10496_2 = {pp112[113]};
    Full_Adder FA_10496(s10496, c10496, in10496_1, in10496_2, pp110[115]);
    wire[0:0] s10497, in10497_1, in10497_2;
    wire c10497;
    assign in10497_1 = {pp100[126]};
    assign in10497_2 = {pp101[125]};
    Full_Adder FA_10497(s10497, c10497, in10497_1, in10497_2, pp99[127]);
    wire[0:0] s10498, in10498_1, in10498_2;
    wire c10498;
    assign in10498_1 = {pp103[123]};
    assign in10498_2 = {pp104[122]};
    Full_Adder FA_10498(s10498, c10498, in10498_1, in10498_2, pp102[124]);
    wire[0:0] s10499, in10499_1, in10499_2;
    wire c10499;
    assign in10499_1 = {pp106[120]};
    assign in10499_2 = {pp107[119]};
    Full_Adder FA_10499(s10499, c10499, in10499_1, in10499_2, pp105[121]);
    wire[0:0] s10500, in10500_1, in10500_2;
    wire c10500;
    assign in10500_1 = {pp109[117]};
    assign in10500_2 = {pp110[116]};
    Full_Adder FA_10500(s10500, c10500, in10500_1, in10500_2, pp108[118]);
    wire[0:0] s10501, in10501_1, in10501_2;
    wire c10501;
    assign in10501_1 = {pp101[126]};
    assign in10501_2 = {pp102[125]};
    Full_Adder FA_10501(s10501, c10501, in10501_1, in10501_2, pp100[127]);
    wire[0:0] s10502, in10502_1, in10502_2;
    wire c10502;
    assign in10502_1 = {pp104[123]};
    assign in10502_2 = {pp105[122]};
    Full_Adder FA_10502(s10502, c10502, in10502_1, in10502_2, pp103[124]);
    wire[0:0] s10503, in10503_1, in10503_2;
    wire c10503;
    assign in10503_1 = {pp107[120]};
    assign in10503_2 = {pp108[119]};
    Full_Adder FA_10503(s10503, c10503, in10503_1, in10503_2, pp106[121]);
    wire[0:0] s10504, in10504_1, in10504_2;
    wire c10504;
    assign in10504_1 = {pp102[126]};
    assign in10504_2 = {pp103[125]};
    Full_Adder FA_10504(s10504, c10504, in10504_1, in10504_2, pp101[127]);
    wire[0:0] s10505, in10505_1, in10505_2;
    wire c10505;
    assign in10505_1 = {pp105[123]};
    assign in10505_2 = {pp106[122]};
    Full_Adder FA_10505(s10505, c10505, in10505_1, in10505_2, pp104[124]);
    wire[0:0] s10506, in10506_1, in10506_2;
    wire c10506;
    assign in10506_1 = {pp103[126]};
    assign in10506_2 = {pp104[125]};
    Full_Adder FA_10506(s10506, c10506, in10506_1, in10506_2, pp102[127]);

    /*Stage 5*/
    wire[0:0] s10507, in10507_1, in10507_2;
    wire c10507;
    assign in10507_1 = {pp0[18]};
    assign in10507_2 = {pp1[17]};
    Half_Adder HA_10507(s10507, c10507, in10507_1, in10507_2);
    wire[0:0] s10508, in10508_1, in10508_2;
    wire c10508;
    assign in10508_1 = {pp1[18]};
    assign in10508_2 = {pp2[17]};
    Full_Adder FA_10508(s10508, c10508, in10508_1, in10508_2, pp0[19]);
    wire[0:0] s10509, in10509_1, in10509_2;
    wire c10509;
    assign in10509_1 = {pp3[16]};
    assign in10509_2 = {pp4[15]};
    Half_Adder HA_10509(s10509, c10509, in10509_1, in10509_2);
    wire[0:0] s10510, in10510_1, in10510_2;
    wire c10510;
    assign in10510_1 = {pp1[19]};
    assign in10510_2 = {pp2[18]};
    Full_Adder FA_10510(s10510, c10510, in10510_1, in10510_2, pp0[20]);
    wire[0:0] s10511, in10511_1, in10511_2;
    wire c10511;
    assign in10511_1 = {pp4[16]};
    assign in10511_2 = {pp5[15]};
    Full_Adder FA_10511(s10511, c10511, in10511_1, in10511_2, pp3[17]);
    wire[0:0] s10512, in10512_1, in10512_2;
    wire c10512;
    assign in10512_1 = {pp6[14]};
    assign in10512_2 = {pp7[13]};
    Half_Adder HA_10512(s10512, c10512, in10512_1, in10512_2);
    wire[0:0] s10513, in10513_1, in10513_2;
    wire c10513;
    assign in10513_1 = {pp1[20]};
    assign in10513_2 = {pp2[19]};
    Full_Adder FA_10513(s10513, c10513, in10513_1, in10513_2, pp0[21]);
    wire[0:0] s10514, in10514_1, in10514_2;
    wire c10514;
    assign in10514_1 = {pp4[17]};
    assign in10514_2 = {pp5[16]};
    Full_Adder FA_10514(s10514, c10514, in10514_1, in10514_2, pp3[18]);
    wire[0:0] s10515, in10515_1, in10515_2;
    wire c10515;
    assign in10515_1 = {pp7[14]};
    assign in10515_2 = {pp8[13]};
    Full_Adder FA_10515(s10515, c10515, in10515_1, in10515_2, pp6[15]);
    wire[0:0] s10516, in10516_1, in10516_2;
    wire c10516;
    assign in10516_1 = {pp9[12]};
    assign in10516_2 = {pp10[11]};
    Half_Adder HA_10516(s10516, c10516, in10516_1, in10516_2);
    wire[0:0] s10517, in10517_1, in10517_2;
    wire c10517;
    assign in10517_1 = {pp1[21]};
    assign in10517_2 = {pp2[20]};
    Full_Adder FA_10517(s10517, c10517, in10517_1, in10517_2, pp0[22]);
    wire[0:0] s10518, in10518_1, in10518_2;
    wire c10518;
    assign in10518_1 = {pp4[18]};
    assign in10518_2 = {pp5[17]};
    Full_Adder FA_10518(s10518, c10518, in10518_1, in10518_2, pp3[19]);
    wire[0:0] s10519, in10519_1, in10519_2;
    wire c10519;
    assign in10519_1 = {pp7[15]};
    assign in10519_2 = {pp8[14]};
    Full_Adder FA_10519(s10519, c10519, in10519_1, in10519_2, pp6[16]);
    wire[0:0] s10520, in10520_1, in10520_2;
    wire c10520;
    assign in10520_1 = {pp10[12]};
    assign in10520_2 = {pp11[11]};
    Full_Adder FA_10520(s10520, c10520, in10520_1, in10520_2, pp9[13]);
    wire[0:0] s10521, in10521_1, in10521_2;
    wire c10521;
    assign in10521_1 = {pp12[10]};
    assign in10521_2 = {pp13[9]};
    Half_Adder HA_10521(s10521, c10521, in10521_1, in10521_2);
    wire[0:0] s10522, in10522_1, in10522_2;
    wire c10522;
    assign in10522_1 = {pp1[22]};
    assign in10522_2 = {pp2[21]};
    Full_Adder FA_10522(s10522, c10522, in10522_1, in10522_2, pp0[23]);
    wire[0:0] s10523, in10523_1, in10523_2;
    wire c10523;
    assign in10523_1 = {pp4[19]};
    assign in10523_2 = {pp5[18]};
    Full_Adder FA_10523(s10523, c10523, in10523_1, in10523_2, pp3[20]);
    wire[0:0] s10524, in10524_1, in10524_2;
    wire c10524;
    assign in10524_1 = {pp7[16]};
    assign in10524_2 = {pp8[15]};
    Full_Adder FA_10524(s10524, c10524, in10524_1, in10524_2, pp6[17]);
    wire[0:0] s10525, in10525_1, in10525_2;
    wire c10525;
    assign in10525_1 = {pp10[13]};
    assign in10525_2 = {pp11[12]};
    Full_Adder FA_10525(s10525, c10525, in10525_1, in10525_2, pp9[14]);
    wire[0:0] s10526, in10526_1, in10526_2;
    wire c10526;
    assign in10526_1 = {pp13[10]};
    assign in10526_2 = {pp14[9]};
    Full_Adder FA_10526(s10526, c10526, in10526_1, in10526_2, pp12[11]);
    wire[0:0] s10527, in10527_1, in10527_2;
    wire c10527;
    assign in10527_1 = {pp15[8]};
    assign in10527_2 = {pp16[7]};
    Half_Adder HA_10527(s10527, c10527, in10527_1, in10527_2);
    wire[0:0] s10528, in10528_1, in10528_2;
    wire c10528;
    assign in10528_1 = {pp1[23]};
    assign in10528_2 = {pp2[22]};
    Full_Adder FA_10528(s10528, c10528, in10528_1, in10528_2, pp0[24]);
    wire[0:0] s10529, in10529_1, in10529_2;
    wire c10529;
    assign in10529_1 = {pp4[20]};
    assign in10529_2 = {pp5[19]};
    Full_Adder FA_10529(s10529, c10529, in10529_1, in10529_2, pp3[21]);
    wire[0:0] s10530, in10530_1, in10530_2;
    wire c10530;
    assign in10530_1 = {pp7[17]};
    assign in10530_2 = {pp8[16]};
    Full_Adder FA_10530(s10530, c10530, in10530_1, in10530_2, pp6[18]);
    wire[0:0] s10531, in10531_1, in10531_2;
    wire c10531;
    assign in10531_1 = {pp10[14]};
    assign in10531_2 = {pp11[13]};
    Full_Adder FA_10531(s10531, c10531, in10531_1, in10531_2, pp9[15]);
    wire[0:0] s10532, in10532_1, in10532_2;
    wire c10532;
    assign in10532_1 = {pp13[11]};
    assign in10532_2 = {pp14[10]};
    Full_Adder FA_10532(s10532, c10532, in10532_1, in10532_2, pp12[12]);
    wire[0:0] s10533, in10533_1, in10533_2;
    wire c10533;
    assign in10533_1 = {pp16[8]};
    assign in10533_2 = {pp17[7]};
    Full_Adder FA_10533(s10533, c10533, in10533_1, in10533_2, pp15[9]);
    wire[0:0] s10534, in10534_1, in10534_2;
    wire c10534;
    assign in10534_1 = {pp18[6]};
    assign in10534_2 = {pp19[5]};
    Half_Adder HA_10534(s10534, c10534, in10534_1, in10534_2);
    wire[0:0] s10535, in10535_1, in10535_2;
    wire c10535;
    assign in10535_1 = {pp1[24]};
    assign in10535_2 = {pp2[23]};
    Full_Adder FA_10535(s10535, c10535, in10535_1, in10535_2, pp0[25]);
    wire[0:0] s10536, in10536_1, in10536_2;
    wire c10536;
    assign in10536_1 = {pp4[21]};
    assign in10536_2 = {pp5[20]};
    Full_Adder FA_10536(s10536, c10536, in10536_1, in10536_2, pp3[22]);
    wire[0:0] s10537, in10537_1, in10537_2;
    wire c10537;
    assign in10537_1 = {pp7[18]};
    assign in10537_2 = {pp8[17]};
    Full_Adder FA_10537(s10537, c10537, in10537_1, in10537_2, pp6[19]);
    wire[0:0] s10538, in10538_1, in10538_2;
    wire c10538;
    assign in10538_1 = {pp10[15]};
    assign in10538_2 = {pp11[14]};
    Full_Adder FA_10538(s10538, c10538, in10538_1, in10538_2, pp9[16]);
    wire[0:0] s10539, in10539_1, in10539_2;
    wire c10539;
    assign in10539_1 = {pp13[12]};
    assign in10539_2 = {pp14[11]};
    Full_Adder FA_10539(s10539, c10539, in10539_1, in10539_2, pp12[13]);
    wire[0:0] s10540, in10540_1, in10540_2;
    wire c10540;
    assign in10540_1 = {pp16[9]};
    assign in10540_2 = {pp17[8]};
    Full_Adder FA_10540(s10540, c10540, in10540_1, in10540_2, pp15[10]);
    wire[0:0] s10541, in10541_1, in10541_2;
    wire c10541;
    assign in10541_1 = {pp19[6]};
    assign in10541_2 = {pp20[5]};
    Full_Adder FA_10541(s10541, c10541, in10541_1, in10541_2, pp18[7]);
    wire[0:0] s10542, in10542_1, in10542_2;
    wire c10542;
    assign in10542_1 = {pp21[4]};
    assign in10542_2 = {pp22[3]};
    Half_Adder HA_10542(s10542, c10542, in10542_1, in10542_2);
    wire[0:0] s10543, in10543_1, in10543_2;
    wire c10543;
    assign in10543_1 = {pp3[23]};
    assign in10543_2 = {pp4[22]};
    Full_Adder FA_10543(s10543, c10543, in10543_1, in10543_2, pp2[24]);
    wire[0:0] s10544, in10544_1, in10544_2;
    wire c10544;
    assign in10544_1 = {pp6[20]};
    assign in10544_2 = {pp7[19]};
    Full_Adder FA_10544(s10544, c10544, in10544_1, in10544_2, pp5[21]);
    wire[0:0] s10545, in10545_1, in10545_2;
    wire c10545;
    assign in10545_1 = {pp9[17]};
    assign in10545_2 = {pp10[16]};
    Full_Adder FA_10545(s10545, c10545, in10545_1, in10545_2, pp8[18]);
    wire[0:0] s10546, in10546_1, in10546_2;
    wire c10546;
    assign in10546_1 = {pp12[14]};
    assign in10546_2 = {pp13[13]};
    Full_Adder FA_10546(s10546, c10546, in10546_1, in10546_2, pp11[15]);
    wire[0:0] s10547, in10547_1, in10547_2;
    wire c10547;
    assign in10547_1 = {pp15[11]};
    assign in10547_2 = {pp16[10]};
    Full_Adder FA_10547(s10547, c10547, in10547_1, in10547_2, pp14[12]);
    wire[0:0] s10548, in10548_1, in10548_2;
    wire c10548;
    assign in10548_1 = {pp18[8]};
    assign in10548_2 = {pp19[7]};
    Full_Adder FA_10548(s10548, c10548, in10548_1, in10548_2, pp17[9]);
    wire[0:0] s10549, in10549_1, in10549_2;
    wire c10549;
    assign in10549_1 = {pp21[5]};
    assign in10549_2 = {pp22[4]};
    Full_Adder FA_10549(s10549, c10549, in10549_1, in10549_2, pp20[6]);
    wire[0:0] s10550, in10550_1, in10550_2;
    wire c10550;
    assign in10550_1 = {pp24[2]};
    assign in10550_2 = {pp25[1]};
    Full_Adder FA_10550(s10550, c10550, in10550_1, in10550_2, pp23[3]);
    wire[0:0] s10551, in10551_1, in10551_2;
    wire c10551;
    assign in10551_1 = {pp6[21]};
    assign in10551_2 = {pp7[20]};
    Full_Adder FA_10551(s10551, c10551, in10551_1, in10551_2, pp5[22]);
    wire[0:0] s10552, in10552_1, in10552_2;
    wire c10552;
    assign in10552_1 = {pp9[18]};
    assign in10552_2 = {pp10[17]};
    Full_Adder FA_10552(s10552, c10552, in10552_1, in10552_2, pp8[19]);
    wire[0:0] s10553, in10553_1, in10553_2;
    wire c10553;
    assign in10553_1 = {pp12[15]};
    assign in10553_2 = {pp13[14]};
    Full_Adder FA_10553(s10553, c10553, in10553_1, in10553_2, pp11[16]);
    wire[0:0] s10554, in10554_1, in10554_2;
    wire c10554;
    assign in10554_1 = {pp15[12]};
    assign in10554_2 = {pp16[11]};
    Full_Adder FA_10554(s10554, c10554, in10554_1, in10554_2, pp14[13]);
    wire[0:0] s10555, in10555_1, in10555_2;
    wire c10555;
    assign in10555_1 = {pp18[9]};
    assign in10555_2 = {pp19[8]};
    Full_Adder FA_10555(s10555, c10555, in10555_1, in10555_2, pp17[10]);
    wire[0:0] s10556, in10556_1, in10556_2;
    wire c10556;
    assign in10556_1 = {pp21[6]};
    assign in10556_2 = {pp22[5]};
    Full_Adder FA_10556(s10556, c10556, in10556_1, in10556_2, pp20[7]);
    wire[0:0] s10557, in10557_1, in10557_2;
    wire c10557;
    assign in10557_1 = {pp24[3]};
    assign in10557_2 = {pp25[2]};
    Full_Adder FA_10557(s10557, c10557, in10557_1, in10557_2, pp23[4]);
    wire[0:0] s10558, in10558_1, in10558_2;
    wire c10558;
    assign in10558_1 = {pp27[0]};
    assign in10558_2 = {c8011};
    Full_Adder FA_10558(s10558, c10558, in10558_1, in10558_2, pp26[1]);
    wire[0:0] s10559, in10559_1, in10559_2;
    wire c10559;
    assign in10559_1 = {pp9[19]};
    assign in10559_2 = {pp10[18]};
    Full_Adder FA_10559(s10559, c10559, in10559_1, in10559_2, pp8[20]);
    wire[0:0] s10560, in10560_1, in10560_2;
    wire c10560;
    assign in10560_1 = {pp12[16]};
    assign in10560_2 = {pp13[15]};
    Full_Adder FA_10560(s10560, c10560, in10560_1, in10560_2, pp11[17]);
    wire[0:0] s10561, in10561_1, in10561_2;
    wire c10561;
    assign in10561_1 = {pp15[13]};
    assign in10561_2 = {pp16[12]};
    Full_Adder FA_10561(s10561, c10561, in10561_1, in10561_2, pp14[14]);
    wire[0:0] s10562, in10562_1, in10562_2;
    wire c10562;
    assign in10562_1 = {pp18[10]};
    assign in10562_2 = {pp19[9]};
    Full_Adder FA_10562(s10562, c10562, in10562_1, in10562_2, pp17[11]);
    wire[0:0] s10563, in10563_1, in10563_2;
    wire c10563;
    assign in10563_1 = {pp21[7]};
    assign in10563_2 = {pp22[6]};
    Full_Adder FA_10563(s10563, c10563, in10563_1, in10563_2, pp20[8]);
    wire[0:0] s10564, in10564_1, in10564_2;
    wire c10564;
    assign in10564_1 = {pp24[4]};
    assign in10564_2 = {pp25[3]};
    Full_Adder FA_10564(s10564, c10564, in10564_1, in10564_2, pp23[5]);
    wire[0:0] s10565, in10565_1, in10565_2;
    wire c10565;
    assign in10565_1 = {pp27[1]};
    assign in10565_2 = {pp28[0]};
    Full_Adder FA_10565(s10565, c10565, in10565_1, in10565_2, pp26[2]);
    wire[0:0] s10566, in10566_1, in10566_2;
    wire c10566;
    assign in10566_1 = {c8013};
    assign in10566_2 = {s8014[0]};
    Full_Adder FA_10566(s10566, c10566, in10566_1, in10566_2, c8012);
    wire[0:0] s10567, in10567_1, in10567_2;
    wire c10567;
    assign in10567_1 = {pp12[17]};
    assign in10567_2 = {pp13[16]};
    Full_Adder FA_10567(s10567, c10567, in10567_1, in10567_2, pp11[18]);
    wire[0:0] s10568, in10568_1, in10568_2;
    wire c10568;
    assign in10568_1 = {pp15[14]};
    assign in10568_2 = {pp16[13]};
    Full_Adder FA_10568(s10568, c10568, in10568_1, in10568_2, pp14[15]);
    wire[0:0] s10569, in10569_1, in10569_2;
    wire c10569;
    assign in10569_1 = {pp18[11]};
    assign in10569_2 = {pp19[10]};
    Full_Adder FA_10569(s10569, c10569, in10569_1, in10569_2, pp17[12]);
    wire[0:0] s10570, in10570_1, in10570_2;
    wire c10570;
    assign in10570_1 = {pp21[8]};
    assign in10570_2 = {pp22[7]};
    Full_Adder FA_10570(s10570, c10570, in10570_1, in10570_2, pp20[9]);
    wire[0:0] s10571, in10571_1, in10571_2;
    wire c10571;
    assign in10571_1 = {pp24[5]};
    assign in10571_2 = {pp25[4]};
    Full_Adder FA_10571(s10571, c10571, in10571_1, in10571_2, pp23[6]);
    wire[0:0] s10572, in10572_1, in10572_2;
    wire c10572;
    assign in10572_1 = {pp27[2]};
    assign in10572_2 = {pp28[1]};
    Full_Adder FA_10572(s10572, c10572, in10572_1, in10572_2, pp26[3]);
    wire[0:0] s10573, in10573_1, in10573_2;
    wire c10573;
    assign in10573_1 = {c8014};
    assign in10573_2 = {c8015};
    Full_Adder FA_10573(s10573, c10573, in10573_1, in10573_2, pp29[0]);
    wire[0:0] s10574, in10574_1, in10574_2;
    wire c10574;
    assign in10574_1 = {s8017[0]};
    assign in10574_2 = {s8018[0]};
    Full_Adder FA_10574(s10574, c10574, in10574_1, in10574_2, c8016);
    wire[0:0] s10575, in10575_1, in10575_2;
    wire c10575;
    assign in10575_1 = {pp15[15]};
    assign in10575_2 = {pp16[14]};
    Full_Adder FA_10575(s10575, c10575, in10575_1, in10575_2, pp14[16]);
    wire[0:0] s10576, in10576_1, in10576_2;
    wire c10576;
    assign in10576_1 = {pp18[12]};
    assign in10576_2 = {pp19[11]};
    Full_Adder FA_10576(s10576, c10576, in10576_1, in10576_2, pp17[13]);
    wire[0:0] s10577, in10577_1, in10577_2;
    wire c10577;
    assign in10577_1 = {pp21[9]};
    assign in10577_2 = {pp22[8]};
    Full_Adder FA_10577(s10577, c10577, in10577_1, in10577_2, pp20[10]);
    wire[0:0] s10578, in10578_1, in10578_2;
    wire c10578;
    assign in10578_1 = {pp24[6]};
    assign in10578_2 = {pp25[5]};
    Full_Adder FA_10578(s10578, c10578, in10578_1, in10578_2, pp23[7]);
    wire[0:0] s10579, in10579_1, in10579_2;
    wire c10579;
    assign in10579_1 = {pp27[3]};
    assign in10579_2 = {pp28[2]};
    Full_Adder FA_10579(s10579, c10579, in10579_1, in10579_2, pp26[4]);
    wire[0:0] s10580, in10580_1, in10580_2;
    wire c10580;
    assign in10580_1 = {pp30[0]};
    assign in10580_2 = {c8017};
    Full_Adder FA_10580(s10580, c10580, in10580_1, in10580_2, pp29[1]);
    wire[0:0] s10581, in10581_1, in10581_2;
    wire c10581;
    assign in10581_1 = {c8019};
    assign in10581_2 = {c8020};
    Full_Adder FA_10581(s10581, c10581, in10581_1, in10581_2, c8018);
    wire[0:0] s10582, in10582_1, in10582_2;
    wire c10582;
    assign in10582_1 = {s8022[0]};
    assign in10582_2 = {s8023[0]};
    Full_Adder FA_10582(s10582, c10582, in10582_1, in10582_2, s8021[0]);
    wire[0:0] s10583, in10583_1, in10583_2;
    wire c10583;
    assign in10583_1 = {pp18[13]};
    assign in10583_2 = {pp19[12]};
    Full_Adder FA_10583(s10583, c10583, in10583_1, in10583_2, pp17[14]);
    wire[0:0] s10584, in10584_1, in10584_2;
    wire c10584;
    assign in10584_1 = {pp21[10]};
    assign in10584_2 = {pp22[9]};
    Full_Adder FA_10584(s10584, c10584, in10584_1, in10584_2, pp20[11]);
    wire[0:0] s10585, in10585_1, in10585_2;
    wire c10585;
    assign in10585_1 = {pp24[7]};
    assign in10585_2 = {pp25[6]};
    Full_Adder FA_10585(s10585, c10585, in10585_1, in10585_2, pp23[8]);
    wire[0:0] s10586, in10586_1, in10586_2;
    wire c10586;
    assign in10586_1 = {pp27[4]};
    assign in10586_2 = {pp28[3]};
    Full_Adder FA_10586(s10586, c10586, in10586_1, in10586_2, pp26[5]);
    wire[0:0] s10587, in10587_1, in10587_2;
    wire c10587;
    assign in10587_1 = {pp30[1]};
    assign in10587_2 = {pp31[0]};
    Full_Adder FA_10587(s10587, c10587, in10587_1, in10587_2, pp29[2]);
    wire[0:0] s10588, in10588_1, in10588_2;
    wire c10588;
    assign in10588_1 = {c8022};
    assign in10588_2 = {c8023};
    Full_Adder FA_10588(s10588, c10588, in10588_1, in10588_2, c8021);
    wire[0:0] s10589, in10589_1, in10589_2;
    wire c10589;
    assign in10589_1 = {c8025};
    assign in10589_2 = {s8026[0]};
    Full_Adder FA_10589(s10589, c10589, in10589_1, in10589_2, c8024);
    wire[0:0] s10590, in10590_1, in10590_2;
    wire c10590;
    assign in10590_1 = {s8028[0]};
    assign in10590_2 = {s8029[0]};
    Full_Adder FA_10590(s10590, c10590, in10590_1, in10590_2, s8027[0]);
    wire[0:0] s10591, in10591_1, in10591_2;
    wire c10591;
    assign in10591_1 = {pp21[11]};
    assign in10591_2 = {pp22[10]};
    Full_Adder FA_10591(s10591, c10591, in10591_1, in10591_2, pp20[12]);
    wire[0:0] s10592, in10592_1, in10592_2;
    wire c10592;
    assign in10592_1 = {pp24[8]};
    assign in10592_2 = {pp25[7]};
    Full_Adder FA_10592(s10592, c10592, in10592_1, in10592_2, pp23[9]);
    wire[0:0] s10593, in10593_1, in10593_2;
    wire c10593;
    assign in10593_1 = {pp27[5]};
    assign in10593_2 = {pp28[4]};
    Full_Adder FA_10593(s10593, c10593, in10593_1, in10593_2, pp26[6]);
    wire[0:0] s10594, in10594_1, in10594_2;
    wire c10594;
    assign in10594_1 = {pp30[2]};
    assign in10594_2 = {pp31[1]};
    Full_Adder FA_10594(s10594, c10594, in10594_1, in10594_2, pp29[3]);
    wire[0:0] s10595, in10595_1, in10595_2;
    wire c10595;
    assign in10595_1 = {c8026};
    assign in10595_2 = {c8027};
    Full_Adder FA_10595(s10595, c10595, in10595_1, in10595_2, pp32[0]);
    wire[0:0] s10596, in10596_1, in10596_2;
    wire c10596;
    assign in10596_1 = {c8029};
    assign in10596_2 = {c8030};
    Full_Adder FA_10596(s10596, c10596, in10596_1, in10596_2, c8028);
    wire[0:0] s10597, in10597_1, in10597_2;
    wire c10597;
    assign in10597_1 = {s8032[0]};
    assign in10597_2 = {s8033[0]};
    Full_Adder FA_10597(s10597, c10597, in10597_1, in10597_2, c8031);
    wire[0:0] s10598, in10598_1, in10598_2;
    wire c10598;
    assign in10598_1 = {s8035[0]};
    assign in10598_2 = {s8036[0]};
    Full_Adder FA_10598(s10598, c10598, in10598_1, in10598_2, s8034[0]);
    wire[0:0] s10599, in10599_1, in10599_2;
    wire c10599;
    assign in10599_1 = {pp24[9]};
    assign in10599_2 = {pp25[8]};
    Full_Adder FA_10599(s10599, c10599, in10599_1, in10599_2, pp23[10]);
    wire[0:0] s10600, in10600_1, in10600_2;
    wire c10600;
    assign in10600_1 = {pp27[6]};
    assign in10600_2 = {pp28[5]};
    Full_Adder FA_10600(s10600, c10600, in10600_1, in10600_2, pp26[7]);
    wire[0:0] s10601, in10601_1, in10601_2;
    wire c10601;
    assign in10601_1 = {pp30[3]};
    assign in10601_2 = {pp31[2]};
    Full_Adder FA_10601(s10601, c10601, in10601_1, in10601_2, pp29[4]);
    wire[0:0] s10602, in10602_1, in10602_2;
    wire c10602;
    assign in10602_1 = {pp33[0]};
    assign in10602_2 = {c8032};
    Full_Adder FA_10602(s10602, c10602, in10602_1, in10602_2, pp32[1]);
    wire[0:0] s10603, in10603_1, in10603_2;
    wire c10603;
    assign in10603_1 = {c8034};
    assign in10603_2 = {c8035};
    Full_Adder FA_10603(s10603, c10603, in10603_1, in10603_2, c8033);
    wire[0:0] s10604, in10604_1, in10604_2;
    wire c10604;
    assign in10604_1 = {c8037};
    assign in10604_2 = {c8038};
    Full_Adder FA_10604(s10604, c10604, in10604_1, in10604_2, c8036);
    wire[0:0] s10605, in10605_1, in10605_2;
    wire c10605;
    assign in10605_1 = {s8040[0]};
    assign in10605_2 = {s8041[0]};
    Full_Adder FA_10605(s10605, c10605, in10605_1, in10605_2, s8039[0]);
    wire[0:0] s10606, in10606_1, in10606_2;
    wire c10606;
    assign in10606_1 = {s8043[0]};
    assign in10606_2 = {s8044[0]};
    Full_Adder FA_10606(s10606, c10606, in10606_1, in10606_2, s8042[0]);
    wire[0:0] s10607, in10607_1, in10607_2;
    wire c10607;
    assign in10607_1 = {pp27[7]};
    assign in10607_2 = {pp28[6]};
    Full_Adder FA_10607(s10607, c10607, in10607_1, in10607_2, pp26[8]);
    wire[0:0] s10608, in10608_1, in10608_2;
    wire c10608;
    assign in10608_1 = {pp30[4]};
    assign in10608_2 = {pp31[3]};
    Full_Adder FA_10608(s10608, c10608, in10608_1, in10608_2, pp29[5]);
    wire[0:0] s10609, in10609_1, in10609_2;
    wire c10609;
    assign in10609_1 = {pp33[1]};
    assign in10609_2 = {pp34[0]};
    Full_Adder FA_10609(s10609, c10609, in10609_1, in10609_2, pp32[2]);
    wire[0:0] s10610, in10610_1, in10610_2;
    wire c10610;
    assign in10610_1 = {c8040};
    assign in10610_2 = {c8041};
    Full_Adder FA_10610(s10610, c10610, in10610_1, in10610_2, c8039);
    wire[0:0] s10611, in10611_1, in10611_2;
    wire c10611;
    assign in10611_1 = {c8043};
    assign in10611_2 = {c8044};
    Full_Adder FA_10611(s10611, c10611, in10611_1, in10611_2, c8042);
    wire[0:0] s10612, in10612_1, in10612_2;
    wire c10612;
    assign in10612_1 = {c8046};
    assign in10612_2 = {s8047[0]};
    Full_Adder FA_10612(s10612, c10612, in10612_1, in10612_2, c8045);
    wire[0:0] s10613, in10613_1, in10613_2;
    wire c10613;
    assign in10613_1 = {s8049[0]};
    assign in10613_2 = {s8050[0]};
    Full_Adder FA_10613(s10613, c10613, in10613_1, in10613_2, s8048[0]);
    wire[0:0] s10614, in10614_1, in10614_2;
    wire c10614;
    assign in10614_1 = {s8052[0]};
    assign in10614_2 = {s8053[0]};
    Full_Adder FA_10614(s10614, c10614, in10614_1, in10614_2, s8051[0]);
    wire[0:0] s10615, in10615_1, in10615_2;
    wire c10615;
    assign in10615_1 = {pp30[5]};
    assign in10615_2 = {pp31[4]};
    Full_Adder FA_10615(s10615, c10615, in10615_1, in10615_2, pp29[6]);
    wire[0:0] s10616, in10616_1, in10616_2;
    wire c10616;
    assign in10616_1 = {pp33[2]};
    assign in10616_2 = {pp34[1]};
    Full_Adder FA_10616(s10616, c10616, in10616_1, in10616_2, pp32[3]);
    wire[0:0] s10617, in10617_1, in10617_2;
    wire c10617;
    assign in10617_1 = {c8047};
    assign in10617_2 = {c8048};
    Full_Adder FA_10617(s10617, c10617, in10617_1, in10617_2, pp35[0]);
    wire[0:0] s10618, in10618_1, in10618_2;
    wire c10618;
    assign in10618_1 = {c8050};
    assign in10618_2 = {c8051};
    Full_Adder FA_10618(s10618, c10618, in10618_1, in10618_2, c8049);
    wire[0:0] s10619, in10619_1, in10619_2;
    wire c10619;
    assign in10619_1 = {c8053};
    assign in10619_2 = {c8054};
    Full_Adder FA_10619(s10619, c10619, in10619_1, in10619_2, c8052);
    wire[0:0] s10620, in10620_1, in10620_2;
    wire c10620;
    assign in10620_1 = {s8056[0]};
    assign in10620_2 = {s8057[0]};
    Full_Adder FA_10620(s10620, c10620, in10620_1, in10620_2, c8055);
    wire[0:0] s10621, in10621_1, in10621_2;
    wire c10621;
    assign in10621_1 = {s8059[0]};
    assign in10621_2 = {s8060[0]};
    Full_Adder FA_10621(s10621, c10621, in10621_1, in10621_2, s8058[0]);
    wire[0:0] s10622, in10622_1, in10622_2;
    wire c10622;
    assign in10622_1 = {s8062[0]};
    assign in10622_2 = {s8063[0]};
    Full_Adder FA_10622(s10622, c10622, in10622_1, in10622_2, s8061[0]);
    wire[0:0] s10623, in10623_1, in10623_2;
    wire c10623;
    assign in10623_1 = {pp33[3]};
    assign in10623_2 = {pp34[2]};
    Full_Adder FA_10623(s10623, c10623, in10623_1, in10623_2, pp32[4]);
    wire[0:0] s10624, in10624_1, in10624_2;
    wire c10624;
    assign in10624_1 = {pp36[0]};
    assign in10624_2 = {c8056};
    Full_Adder FA_10624(s10624, c10624, in10624_1, in10624_2, pp35[1]);
    wire[0:0] s10625, in10625_1, in10625_2;
    wire c10625;
    assign in10625_1 = {c8058};
    assign in10625_2 = {c8059};
    Full_Adder FA_10625(s10625, c10625, in10625_1, in10625_2, c8057);
    wire[0:0] s10626, in10626_1, in10626_2;
    wire c10626;
    assign in10626_1 = {c8061};
    assign in10626_2 = {c8062};
    Full_Adder FA_10626(s10626, c10626, in10626_1, in10626_2, c8060);
    wire[0:0] s10627, in10627_1, in10627_2;
    wire c10627;
    assign in10627_1 = {c8064};
    assign in10627_2 = {c8065};
    Full_Adder FA_10627(s10627, c10627, in10627_1, in10627_2, c8063);
    wire[0:0] s10628, in10628_1, in10628_2;
    wire c10628;
    assign in10628_1 = {s8067[0]};
    assign in10628_2 = {s8068[0]};
    Full_Adder FA_10628(s10628, c10628, in10628_1, in10628_2, s8066[0]);
    wire[0:0] s10629, in10629_1, in10629_2;
    wire c10629;
    assign in10629_1 = {s8070[0]};
    assign in10629_2 = {s8071[0]};
    Full_Adder FA_10629(s10629, c10629, in10629_1, in10629_2, s8069[0]);
    wire[0:0] s10630, in10630_1, in10630_2;
    wire c10630;
    assign in10630_1 = {s8073[0]};
    assign in10630_2 = {s8074[0]};
    Full_Adder FA_10630(s10630, c10630, in10630_1, in10630_2, s8072[0]);
    wire[0:0] s10631, in10631_1, in10631_2;
    wire c10631;
    assign in10631_1 = {pp36[1]};
    assign in10631_2 = {pp37[0]};
    Full_Adder FA_10631(s10631, c10631, in10631_1, in10631_2, pp35[2]);
    wire[0:0] s10632, in10632_1, in10632_2;
    wire c10632;
    assign in10632_1 = {c8067};
    assign in10632_2 = {c8068};
    Full_Adder FA_10632(s10632, c10632, in10632_1, in10632_2, c8066);
    wire[0:0] s10633, in10633_1, in10633_2;
    wire c10633;
    assign in10633_1 = {c8070};
    assign in10633_2 = {c8071};
    Full_Adder FA_10633(s10633, c10633, in10633_1, in10633_2, c8069);
    wire[0:0] s10634, in10634_1, in10634_2;
    wire c10634;
    assign in10634_1 = {c8073};
    assign in10634_2 = {c8074};
    Full_Adder FA_10634(s10634, c10634, in10634_1, in10634_2, c8072);
    wire[0:0] s10635, in10635_1, in10635_2;
    wire c10635;
    assign in10635_1 = {c8076};
    assign in10635_2 = {s8077[0]};
    Full_Adder FA_10635(s10635, c10635, in10635_1, in10635_2, c8075);
    wire[0:0] s10636, in10636_1, in10636_2;
    wire c10636;
    assign in10636_1 = {s8079[0]};
    assign in10636_2 = {s8080[0]};
    Full_Adder FA_10636(s10636, c10636, in10636_1, in10636_2, s8078[0]);
    wire[0:0] s10637, in10637_1, in10637_2;
    wire c10637;
    assign in10637_1 = {s8082[0]};
    assign in10637_2 = {s8083[0]};
    Full_Adder FA_10637(s10637, c10637, in10637_1, in10637_2, s8081[0]);
    wire[0:0] s10638, in10638_1, in10638_2;
    wire c10638;
    assign in10638_1 = {s8085[0]};
    assign in10638_2 = {s8086[0]};
    Full_Adder FA_10638(s10638, c10638, in10638_1, in10638_2, s8084[0]);
    wire[0:0] s10639, in10639_1, in10639_2;
    wire c10639;
    assign in10639_1 = {c8077};
    assign in10639_2 = {c8078};
    Full_Adder FA_10639(s10639, c10639, in10639_1, in10639_2, pp38[0]);
    wire[0:0] s10640, in10640_1, in10640_2;
    wire c10640;
    assign in10640_1 = {c8080};
    assign in10640_2 = {c8081};
    Full_Adder FA_10640(s10640, c10640, in10640_1, in10640_2, c8079);
    wire[0:0] s10641, in10641_1, in10641_2;
    wire c10641;
    assign in10641_1 = {c8083};
    assign in10641_2 = {c8084};
    Full_Adder FA_10641(s10641, c10641, in10641_1, in10641_2, c8082);
    wire[0:0] s10642, in10642_1, in10642_2;
    wire c10642;
    assign in10642_1 = {c8086};
    assign in10642_2 = {c8087};
    Full_Adder FA_10642(s10642, c10642, in10642_1, in10642_2, c8085);
    wire[0:0] s10643, in10643_1, in10643_2;
    wire c10643;
    assign in10643_1 = {s8089[0]};
    assign in10643_2 = {s8090[0]};
    Full_Adder FA_10643(s10643, c10643, in10643_1, in10643_2, c8088);
    wire[0:0] s10644, in10644_1, in10644_2;
    wire c10644;
    assign in10644_1 = {s8092[0]};
    assign in10644_2 = {s8093[0]};
    Full_Adder FA_10644(s10644, c10644, in10644_1, in10644_2, s8091[0]);
    wire[0:0] s10645, in10645_1, in10645_2;
    wire c10645;
    assign in10645_1 = {s8095[0]};
    assign in10645_2 = {s8096[0]};
    Full_Adder FA_10645(s10645, c10645, in10645_1, in10645_2, s8094[0]);
    wire[0:0] s10646, in10646_1, in10646_2;
    wire c10646;
    assign in10646_1 = {s8098[0]};
    assign in10646_2 = {s8099[0]};
    Full_Adder FA_10646(s10646, c10646, in10646_1, in10646_2, s8097[0]);
    wire[0:0] s10647, in10647_1, in10647_2;
    wire c10647;
    assign in10647_1 = {c8090};
    assign in10647_2 = {c8091};
    Full_Adder FA_10647(s10647, c10647, in10647_1, in10647_2, c8089);
    wire[0:0] s10648, in10648_1, in10648_2;
    wire c10648;
    assign in10648_1 = {c8093};
    assign in10648_2 = {c8094};
    Full_Adder FA_10648(s10648, c10648, in10648_1, in10648_2, c8092);
    wire[0:0] s10649, in10649_1, in10649_2;
    wire c10649;
    assign in10649_1 = {c8096};
    assign in10649_2 = {c8097};
    Full_Adder FA_10649(s10649, c10649, in10649_1, in10649_2, c8095);
    wire[0:0] s10650, in10650_1, in10650_2;
    wire c10650;
    assign in10650_1 = {c8099};
    assign in10650_2 = {c8100};
    Full_Adder FA_10650(s10650, c10650, in10650_1, in10650_2, c8098);
    wire[0:0] s10651, in10651_1, in10651_2;
    wire c10651;
    assign in10651_1 = {s8102[0]};
    assign in10651_2 = {s8103[0]};
    Full_Adder FA_10651(s10651, c10651, in10651_1, in10651_2, c8101);
    wire[0:0] s10652, in10652_1, in10652_2;
    wire c10652;
    assign in10652_1 = {s8105[0]};
    assign in10652_2 = {s8106[0]};
    Full_Adder FA_10652(s10652, c10652, in10652_1, in10652_2, s8104[0]);
    wire[0:0] s10653, in10653_1, in10653_2;
    wire c10653;
    assign in10653_1 = {s8108[0]};
    assign in10653_2 = {s8109[0]};
    Full_Adder FA_10653(s10653, c10653, in10653_1, in10653_2, s8107[0]);
    wire[0:0] s10654, in10654_1, in10654_2;
    wire c10654;
    assign in10654_1 = {s8111[0]};
    assign in10654_2 = {s8112[0]};
    Full_Adder FA_10654(s10654, c10654, in10654_1, in10654_2, s8110[0]);
    wire[0:0] s10655, in10655_1, in10655_2;
    wire c10655;
    assign in10655_1 = {c8103};
    assign in10655_2 = {c8104};
    Full_Adder FA_10655(s10655, c10655, in10655_1, in10655_2, c8102);
    wire[0:0] s10656, in10656_1, in10656_2;
    wire c10656;
    assign in10656_1 = {c8106};
    assign in10656_2 = {c8107};
    Full_Adder FA_10656(s10656, c10656, in10656_1, in10656_2, c8105);
    wire[0:0] s10657, in10657_1, in10657_2;
    wire c10657;
    assign in10657_1 = {c8109};
    assign in10657_2 = {c8110};
    Full_Adder FA_10657(s10657, c10657, in10657_1, in10657_2, c8108);
    wire[0:0] s10658, in10658_1, in10658_2;
    wire c10658;
    assign in10658_1 = {c8112};
    assign in10658_2 = {c8113};
    Full_Adder FA_10658(s10658, c10658, in10658_1, in10658_2, c8111);
    wire[0:0] s10659, in10659_1, in10659_2;
    wire c10659;
    assign in10659_1 = {s8115[0]};
    assign in10659_2 = {s8116[0]};
    Full_Adder FA_10659(s10659, c10659, in10659_1, in10659_2, c8114);
    wire[0:0] s10660, in10660_1, in10660_2;
    wire c10660;
    assign in10660_1 = {s8118[0]};
    assign in10660_2 = {s8119[0]};
    Full_Adder FA_10660(s10660, c10660, in10660_1, in10660_2, s8117[0]);
    wire[0:0] s10661, in10661_1, in10661_2;
    wire c10661;
    assign in10661_1 = {s8121[0]};
    assign in10661_2 = {s8122[0]};
    Full_Adder FA_10661(s10661, c10661, in10661_1, in10661_2, s8120[0]);
    wire[0:0] s10662, in10662_1, in10662_2;
    wire c10662;
    assign in10662_1 = {s8124[0]};
    assign in10662_2 = {s8125[0]};
    Full_Adder FA_10662(s10662, c10662, in10662_1, in10662_2, s8123[0]);
    wire[0:0] s10663, in10663_1, in10663_2;
    wire c10663;
    assign in10663_1 = {c8116};
    assign in10663_2 = {c8117};
    Full_Adder FA_10663(s10663, c10663, in10663_1, in10663_2, c8115);
    wire[0:0] s10664, in10664_1, in10664_2;
    wire c10664;
    assign in10664_1 = {c8119};
    assign in10664_2 = {c8120};
    Full_Adder FA_10664(s10664, c10664, in10664_1, in10664_2, c8118);
    wire[0:0] s10665, in10665_1, in10665_2;
    wire c10665;
    assign in10665_1 = {c8122};
    assign in10665_2 = {c8123};
    Full_Adder FA_10665(s10665, c10665, in10665_1, in10665_2, c8121);
    wire[0:0] s10666, in10666_1, in10666_2;
    wire c10666;
    assign in10666_1 = {c8125};
    assign in10666_2 = {c8126};
    Full_Adder FA_10666(s10666, c10666, in10666_1, in10666_2, c8124);
    wire[0:0] s10667, in10667_1, in10667_2;
    wire c10667;
    assign in10667_1 = {s8128[0]};
    assign in10667_2 = {s8129[0]};
    Full_Adder FA_10667(s10667, c10667, in10667_1, in10667_2, c8127);
    wire[0:0] s10668, in10668_1, in10668_2;
    wire c10668;
    assign in10668_1 = {s8131[0]};
    assign in10668_2 = {s8132[0]};
    Full_Adder FA_10668(s10668, c10668, in10668_1, in10668_2, s8130[0]);
    wire[0:0] s10669, in10669_1, in10669_2;
    wire c10669;
    assign in10669_1 = {s8134[0]};
    assign in10669_2 = {s8135[0]};
    Full_Adder FA_10669(s10669, c10669, in10669_1, in10669_2, s8133[0]);
    wire[0:0] s10670, in10670_1, in10670_2;
    wire c10670;
    assign in10670_1 = {s8137[0]};
    assign in10670_2 = {s8138[0]};
    Full_Adder FA_10670(s10670, c10670, in10670_1, in10670_2, s8136[0]);
    wire[0:0] s10671, in10671_1, in10671_2;
    wire c10671;
    assign in10671_1 = {c8129};
    assign in10671_2 = {c8130};
    Full_Adder FA_10671(s10671, c10671, in10671_1, in10671_2, c8128);
    wire[0:0] s10672, in10672_1, in10672_2;
    wire c10672;
    assign in10672_1 = {c8132};
    assign in10672_2 = {c8133};
    Full_Adder FA_10672(s10672, c10672, in10672_1, in10672_2, c8131);
    wire[0:0] s10673, in10673_1, in10673_2;
    wire c10673;
    assign in10673_1 = {c8135};
    assign in10673_2 = {c8136};
    Full_Adder FA_10673(s10673, c10673, in10673_1, in10673_2, c8134);
    wire[0:0] s10674, in10674_1, in10674_2;
    wire c10674;
    assign in10674_1 = {c8138};
    assign in10674_2 = {c8139};
    Full_Adder FA_10674(s10674, c10674, in10674_1, in10674_2, c8137);
    wire[0:0] s10675, in10675_1, in10675_2;
    wire c10675;
    assign in10675_1 = {s8141[0]};
    assign in10675_2 = {s8142[0]};
    Full_Adder FA_10675(s10675, c10675, in10675_1, in10675_2, c8140);
    wire[0:0] s10676, in10676_1, in10676_2;
    wire c10676;
    assign in10676_1 = {s8144[0]};
    assign in10676_2 = {s8145[0]};
    Full_Adder FA_10676(s10676, c10676, in10676_1, in10676_2, s8143[0]);
    wire[0:0] s10677, in10677_1, in10677_2;
    wire c10677;
    assign in10677_1 = {s8147[0]};
    assign in10677_2 = {s8148[0]};
    Full_Adder FA_10677(s10677, c10677, in10677_1, in10677_2, s8146[0]);
    wire[0:0] s10678, in10678_1, in10678_2;
    wire c10678;
    assign in10678_1 = {s8150[0]};
    assign in10678_2 = {s8151[0]};
    Full_Adder FA_10678(s10678, c10678, in10678_1, in10678_2, s8149[0]);
    wire[0:0] s10679, in10679_1, in10679_2;
    wire c10679;
    assign in10679_1 = {c8142};
    assign in10679_2 = {c8143};
    Full_Adder FA_10679(s10679, c10679, in10679_1, in10679_2, c8141);
    wire[0:0] s10680, in10680_1, in10680_2;
    wire c10680;
    assign in10680_1 = {c8145};
    assign in10680_2 = {c8146};
    Full_Adder FA_10680(s10680, c10680, in10680_1, in10680_2, c8144);
    wire[0:0] s10681, in10681_1, in10681_2;
    wire c10681;
    assign in10681_1 = {c8148};
    assign in10681_2 = {c8149};
    Full_Adder FA_10681(s10681, c10681, in10681_1, in10681_2, c8147);
    wire[0:0] s10682, in10682_1, in10682_2;
    wire c10682;
    assign in10682_1 = {c8151};
    assign in10682_2 = {c8152};
    Full_Adder FA_10682(s10682, c10682, in10682_1, in10682_2, c8150);
    wire[0:0] s10683, in10683_1, in10683_2;
    wire c10683;
    assign in10683_1 = {s8154[0]};
    assign in10683_2 = {s8155[0]};
    Full_Adder FA_10683(s10683, c10683, in10683_1, in10683_2, c8153);
    wire[0:0] s10684, in10684_1, in10684_2;
    wire c10684;
    assign in10684_1 = {s8157[0]};
    assign in10684_2 = {s8158[0]};
    Full_Adder FA_10684(s10684, c10684, in10684_1, in10684_2, s8156[0]);
    wire[0:0] s10685, in10685_1, in10685_2;
    wire c10685;
    assign in10685_1 = {s8160[0]};
    assign in10685_2 = {s8161[0]};
    Full_Adder FA_10685(s10685, c10685, in10685_1, in10685_2, s8159[0]);
    wire[0:0] s10686, in10686_1, in10686_2;
    wire c10686;
    assign in10686_1 = {s8163[0]};
    assign in10686_2 = {s8164[0]};
    Full_Adder FA_10686(s10686, c10686, in10686_1, in10686_2, s8162[0]);
    wire[0:0] s10687, in10687_1, in10687_2;
    wire c10687;
    assign in10687_1 = {c8155};
    assign in10687_2 = {c8156};
    Full_Adder FA_10687(s10687, c10687, in10687_1, in10687_2, c8154);
    wire[0:0] s10688, in10688_1, in10688_2;
    wire c10688;
    assign in10688_1 = {c8158};
    assign in10688_2 = {c8159};
    Full_Adder FA_10688(s10688, c10688, in10688_1, in10688_2, c8157);
    wire[0:0] s10689, in10689_1, in10689_2;
    wire c10689;
    assign in10689_1 = {c8161};
    assign in10689_2 = {c8162};
    Full_Adder FA_10689(s10689, c10689, in10689_1, in10689_2, c8160);
    wire[0:0] s10690, in10690_1, in10690_2;
    wire c10690;
    assign in10690_1 = {c8164};
    assign in10690_2 = {c8165};
    Full_Adder FA_10690(s10690, c10690, in10690_1, in10690_2, c8163);
    wire[0:0] s10691, in10691_1, in10691_2;
    wire c10691;
    assign in10691_1 = {s8167[0]};
    assign in10691_2 = {s8168[0]};
    Full_Adder FA_10691(s10691, c10691, in10691_1, in10691_2, c8166);
    wire[0:0] s10692, in10692_1, in10692_2;
    wire c10692;
    assign in10692_1 = {s8170[0]};
    assign in10692_2 = {s8171[0]};
    Full_Adder FA_10692(s10692, c10692, in10692_1, in10692_2, s8169[0]);
    wire[0:0] s10693, in10693_1, in10693_2;
    wire c10693;
    assign in10693_1 = {s8173[0]};
    assign in10693_2 = {s8174[0]};
    Full_Adder FA_10693(s10693, c10693, in10693_1, in10693_2, s8172[0]);
    wire[0:0] s10694, in10694_1, in10694_2;
    wire c10694;
    assign in10694_1 = {s8176[0]};
    assign in10694_2 = {s8177[0]};
    Full_Adder FA_10694(s10694, c10694, in10694_1, in10694_2, s8175[0]);
    wire[0:0] s10695, in10695_1, in10695_2;
    wire c10695;
    assign in10695_1 = {c8168};
    assign in10695_2 = {c8169};
    Full_Adder FA_10695(s10695, c10695, in10695_1, in10695_2, c8167);
    wire[0:0] s10696, in10696_1, in10696_2;
    wire c10696;
    assign in10696_1 = {c8171};
    assign in10696_2 = {c8172};
    Full_Adder FA_10696(s10696, c10696, in10696_1, in10696_2, c8170);
    wire[0:0] s10697, in10697_1, in10697_2;
    wire c10697;
    assign in10697_1 = {c8174};
    assign in10697_2 = {c8175};
    Full_Adder FA_10697(s10697, c10697, in10697_1, in10697_2, c8173);
    wire[0:0] s10698, in10698_1, in10698_2;
    wire c10698;
    assign in10698_1 = {c8177};
    assign in10698_2 = {c8178};
    Full_Adder FA_10698(s10698, c10698, in10698_1, in10698_2, c8176);
    wire[0:0] s10699, in10699_1, in10699_2;
    wire c10699;
    assign in10699_1 = {s8180[0]};
    assign in10699_2 = {s8181[0]};
    Full_Adder FA_10699(s10699, c10699, in10699_1, in10699_2, c8179);
    wire[0:0] s10700, in10700_1, in10700_2;
    wire c10700;
    assign in10700_1 = {s8183[0]};
    assign in10700_2 = {s8184[0]};
    Full_Adder FA_10700(s10700, c10700, in10700_1, in10700_2, s8182[0]);
    wire[0:0] s10701, in10701_1, in10701_2;
    wire c10701;
    assign in10701_1 = {s8186[0]};
    assign in10701_2 = {s8187[0]};
    Full_Adder FA_10701(s10701, c10701, in10701_1, in10701_2, s8185[0]);
    wire[0:0] s10702, in10702_1, in10702_2;
    wire c10702;
    assign in10702_1 = {s8189[0]};
    assign in10702_2 = {s8190[0]};
    Full_Adder FA_10702(s10702, c10702, in10702_1, in10702_2, s8188[0]);
    wire[0:0] s10703, in10703_1, in10703_2;
    wire c10703;
    assign in10703_1 = {c8181};
    assign in10703_2 = {c8182};
    Full_Adder FA_10703(s10703, c10703, in10703_1, in10703_2, c8180);
    wire[0:0] s10704, in10704_1, in10704_2;
    wire c10704;
    assign in10704_1 = {c8184};
    assign in10704_2 = {c8185};
    Full_Adder FA_10704(s10704, c10704, in10704_1, in10704_2, c8183);
    wire[0:0] s10705, in10705_1, in10705_2;
    wire c10705;
    assign in10705_1 = {c8187};
    assign in10705_2 = {c8188};
    Full_Adder FA_10705(s10705, c10705, in10705_1, in10705_2, c8186);
    wire[0:0] s10706, in10706_1, in10706_2;
    wire c10706;
    assign in10706_1 = {c8190};
    assign in10706_2 = {c8191};
    Full_Adder FA_10706(s10706, c10706, in10706_1, in10706_2, c8189);
    wire[0:0] s10707, in10707_1, in10707_2;
    wire c10707;
    assign in10707_1 = {s8193[0]};
    assign in10707_2 = {s8194[0]};
    Full_Adder FA_10707(s10707, c10707, in10707_1, in10707_2, c8192);
    wire[0:0] s10708, in10708_1, in10708_2;
    wire c10708;
    assign in10708_1 = {s8196[0]};
    assign in10708_2 = {s8197[0]};
    Full_Adder FA_10708(s10708, c10708, in10708_1, in10708_2, s8195[0]);
    wire[0:0] s10709, in10709_1, in10709_2;
    wire c10709;
    assign in10709_1 = {s8199[0]};
    assign in10709_2 = {s8200[0]};
    Full_Adder FA_10709(s10709, c10709, in10709_1, in10709_2, s8198[0]);
    wire[0:0] s10710, in10710_1, in10710_2;
    wire c10710;
    assign in10710_1 = {s8202[0]};
    assign in10710_2 = {s8203[0]};
    Full_Adder FA_10710(s10710, c10710, in10710_1, in10710_2, s8201[0]);
    wire[0:0] s10711, in10711_1, in10711_2;
    wire c10711;
    assign in10711_1 = {c8194};
    assign in10711_2 = {c8195};
    Full_Adder FA_10711(s10711, c10711, in10711_1, in10711_2, c8193);
    wire[0:0] s10712, in10712_1, in10712_2;
    wire c10712;
    assign in10712_1 = {c8197};
    assign in10712_2 = {c8198};
    Full_Adder FA_10712(s10712, c10712, in10712_1, in10712_2, c8196);
    wire[0:0] s10713, in10713_1, in10713_2;
    wire c10713;
    assign in10713_1 = {c8200};
    assign in10713_2 = {c8201};
    Full_Adder FA_10713(s10713, c10713, in10713_1, in10713_2, c8199);
    wire[0:0] s10714, in10714_1, in10714_2;
    wire c10714;
    assign in10714_1 = {c8203};
    assign in10714_2 = {c8204};
    Full_Adder FA_10714(s10714, c10714, in10714_1, in10714_2, c8202);
    wire[0:0] s10715, in10715_1, in10715_2;
    wire c10715;
    assign in10715_1 = {s8206[0]};
    assign in10715_2 = {s8207[0]};
    Full_Adder FA_10715(s10715, c10715, in10715_1, in10715_2, c8205);
    wire[0:0] s10716, in10716_1, in10716_2;
    wire c10716;
    assign in10716_1 = {s8209[0]};
    assign in10716_2 = {s8210[0]};
    Full_Adder FA_10716(s10716, c10716, in10716_1, in10716_2, s8208[0]);
    wire[0:0] s10717, in10717_1, in10717_2;
    wire c10717;
    assign in10717_1 = {s8212[0]};
    assign in10717_2 = {s8213[0]};
    Full_Adder FA_10717(s10717, c10717, in10717_1, in10717_2, s8211[0]);
    wire[0:0] s10718, in10718_1, in10718_2;
    wire c10718;
    assign in10718_1 = {s8215[0]};
    assign in10718_2 = {s8216[0]};
    Full_Adder FA_10718(s10718, c10718, in10718_1, in10718_2, s8214[0]);
    wire[0:0] s10719, in10719_1, in10719_2;
    wire c10719;
    assign in10719_1 = {c8207};
    assign in10719_2 = {c8208};
    Full_Adder FA_10719(s10719, c10719, in10719_1, in10719_2, c8206);
    wire[0:0] s10720, in10720_1, in10720_2;
    wire c10720;
    assign in10720_1 = {c8210};
    assign in10720_2 = {c8211};
    Full_Adder FA_10720(s10720, c10720, in10720_1, in10720_2, c8209);
    wire[0:0] s10721, in10721_1, in10721_2;
    wire c10721;
    assign in10721_1 = {c8213};
    assign in10721_2 = {c8214};
    Full_Adder FA_10721(s10721, c10721, in10721_1, in10721_2, c8212);
    wire[0:0] s10722, in10722_1, in10722_2;
    wire c10722;
    assign in10722_1 = {c8216};
    assign in10722_2 = {c8217};
    Full_Adder FA_10722(s10722, c10722, in10722_1, in10722_2, c8215);
    wire[0:0] s10723, in10723_1, in10723_2;
    wire c10723;
    assign in10723_1 = {s8219[0]};
    assign in10723_2 = {s8220[0]};
    Full_Adder FA_10723(s10723, c10723, in10723_1, in10723_2, c8218);
    wire[0:0] s10724, in10724_1, in10724_2;
    wire c10724;
    assign in10724_1 = {s8222[0]};
    assign in10724_2 = {s8223[0]};
    Full_Adder FA_10724(s10724, c10724, in10724_1, in10724_2, s8221[0]);
    wire[0:0] s10725, in10725_1, in10725_2;
    wire c10725;
    assign in10725_1 = {s8225[0]};
    assign in10725_2 = {s8226[0]};
    Full_Adder FA_10725(s10725, c10725, in10725_1, in10725_2, s8224[0]);
    wire[0:0] s10726, in10726_1, in10726_2;
    wire c10726;
    assign in10726_1 = {s8228[0]};
    assign in10726_2 = {s8229[0]};
    Full_Adder FA_10726(s10726, c10726, in10726_1, in10726_2, s8227[0]);
    wire[0:0] s10727, in10727_1, in10727_2;
    wire c10727;
    assign in10727_1 = {c8220};
    assign in10727_2 = {c8221};
    Full_Adder FA_10727(s10727, c10727, in10727_1, in10727_2, c8219);
    wire[0:0] s10728, in10728_1, in10728_2;
    wire c10728;
    assign in10728_1 = {c8223};
    assign in10728_2 = {c8224};
    Full_Adder FA_10728(s10728, c10728, in10728_1, in10728_2, c8222);
    wire[0:0] s10729, in10729_1, in10729_2;
    wire c10729;
    assign in10729_1 = {c8226};
    assign in10729_2 = {c8227};
    Full_Adder FA_10729(s10729, c10729, in10729_1, in10729_2, c8225);
    wire[0:0] s10730, in10730_1, in10730_2;
    wire c10730;
    assign in10730_1 = {c8229};
    assign in10730_2 = {c8230};
    Full_Adder FA_10730(s10730, c10730, in10730_1, in10730_2, c8228);
    wire[0:0] s10731, in10731_1, in10731_2;
    wire c10731;
    assign in10731_1 = {s8232[0]};
    assign in10731_2 = {s8233[0]};
    Full_Adder FA_10731(s10731, c10731, in10731_1, in10731_2, c8231);
    wire[0:0] s10732, in10732_1, in10732_2;
    wire c10732;
    assign in10732_1 = {s8235[0]};
    assign in10732_2 = {s8236[0]};
    Full_Adder FA_10732(s10732, c10732, in10732_1, in10732_2, s8234[0]);
    wire[0:0] s10733, in10733_1, in10733_2;
    wire c10733;
    assign in10733_1 = {s8238[0]};
    assign in10733_2 = {s8239[0]};
    Full_Adder FA_10733(s10733, c10733, in10733_1, in10733_2, s8237[0]);
    wire[0:0] s10734, in10734_1, in10734_2;
    wire c10734;
    assign in10734_1 = {s8241[0]};
    assign in10734_2 = {s8242[0]};
    Full_Adder FA_10734(s10734, c10734, in10734_1, in10734_2, s8240[0]);
    wire[0:0] s10735, in10735_1, in10735_2;
    wire c10735;
    assign in10735_1 = {c8233};
    assign in10735_2 = {c8234};
    Full_Adder FA_10735(s10735, c10735, in10735_1, in10735_2, c8232);
    wire[0:0] s10736, in10736_1, in10736_2;
    wire c10736;
    assign in10736_1 = {c8236};
    assign in10736_2 = {c8237};
    Full_Adder FA_10736(s10736, c10736, in10736_1, in10736_2, c8235);
    wire[0:0] s10737, in10737_1, in10737_2;
    wire c10737;
    assign in10737_1 = {c8239};
    assign in10737_2 = {c8240};
    Full_Adder FA_10737(s10737, c10737, in10737_1, in10737_2, c8238);
    wire[0:0] s10738, in10738_1, in10738_2;
    wire c10738;
    assign in10738_1 = {c8242};
    assign in10738_2 = {c8243};
    Full_Adder FA_10738(s10738, c10738, in10738_1, in10738_2, c8241);
    wire[0:0] s10739, in10739_1, in10739_2;
    wire c10739;
    assign in10739_1 = {s8245[0]};
    assign in10739_2 = {s8246[0]};
    Full_Adder FA_10739(s10739, c10739, in10739_1, in10739_2, c8244);
    wire[0:0] s10740, in10740_1, in10740_2;
    wire c10740;
    assign in10740_1 = {s8248[0]};
    assign in10740_2 = {s8249[0]};
    Full_Adder FA_10740(s10740, c10740, in10740_1, in10740_2, s8247[0]);
    wire[0:0] s10741, in10741_1, in10741_2;
    wire c10741;
    assign in10741_1 = {s8251[0]};
    assign in10741_2 = {s8252[0]};
    Full_Adder FA_10741(s10741, c10741, in10741_1, in10741_2, s8250[0]);
    wire[0:0] s10742, in10742_1, in10742_2;
    wire c10742;
    assign in10742_1 = {s8254[0]};
    assign in10742_2 = {s8255[0]};
    Full_Adder FA_10742(s10742, c10742, in10742_1, in10742_2, s8253[0]);
    wire[0:0] s10743, in10743_1, in10743_2;
    wire c10743;
    assign in10743_1 = {c8246};
    assign in10743_2 = {c8247};
    Full_Adder FA_10743(s10743, c10743, in10743_1, in10743_2, c8245);
    wire[0:0] s10744, in10744_1, in10744_2;
    wire c10744;
    assign in10744_1 = {c8249};
    assign in10744_2 = {c8250};
    Full_Adder FA_10744(s10744, c10744, in10744_1, in10744_2, c8248);
    wire[0:0] s10745, in10745_1, in10745_2;
    wire c10745;
    assign in10745_1 = {c8252};
    assign in10745_2 = {c8253};
    Full_Adder FA_10745(s10745, c10745, in10745_1, in10745_2, c8251);
    wire[0:0] s10746, in10746_1, in10746_2;
    wire c10746;
    assign in10746_1 = {c8255};
    assign in10746_2 = {c8256};
    Full_Adder FA_10746(s10746, c10746, in10746_1, in10746_2, c8254);
    wire[0:0] s10747, in10747_1, in10747_2;
    wire c10747;
    assign in10747_1 = {s8258[0]};
    assign in10747_2 = {s8259[0]};
    Full_Adder FA_10747(s10747, c10747, in10747_1, in10747_2, c8257);
    wire[0:0] s10748, in10748_1, in10748_2;
    wire c10748;
    assign in10748_1 = {s8261[0]};
    assign in10748_2 = {s8262[0]};
    Full_Adder FA_10748(s10748, c10748, in10748_1, in10748_2, s8260[0]);
    wire[0:0] s10749, in10749_1, in10749_2;
    wire c10749;
    assign in10749_1 = {s8264[0]};
    assign in10749_2 = {s8265[0]};
    Full_Adder FA_10749(s10749, c10749, in10749_1, in10749_2, s8263[0]);
    wire[0:0] s10750, in10750_1, in10750_2;
    wire c10750;
    assign in10750_1 = {s8267[0]};
    assign in10750_2 = {s8268[0]};
    Full_Adder FA_10750(s10750, c10750, in10750_1, in10750_2, s8266[0]);
    wire[0:0] s10751, in10751_1, in10751_2;
    wire c10751;
    assign in10751_1 = {c8259};
    assign in10751_2 = {c8260};
    Full_Adder FA_10751(s10751, c10751, in10751_1, in10751_2, c8258);
    wire[0:0] s10752, in10752_1, in10752_2;
    wire c10752;
    assign in10752_1 = {c8262};
    assign in10752_2 = {c8263};
    Full_Adder FA_10752(s10752, c10752, in10752_1, in10752_2, c8261);
    wire[0:0] s10753, in10753_1, in10753_2;
    wire c10753;
    assign in10753_1 = {c8265};
    assign in10753_2 = {c8266};
    Full_Adder FA_10753(s10753, c10753, in10753_1, in10753_2, c8264);
    wire[0:0] s10754, in10754_1, in10754_2;
    wire c10754;
    assign in10754_1 = {c8268};
    assign in10754_2 = {c8269};
    Full_Adder FA_10754(s10754, c10754, in10754_1, in10754_2, c8267);
    wire[0:0] s10755, in10755_1, in10755_2;
    wire c10755;
    assign in10755_1 = {s8271[0]};
    assign in10755_2 = {s8272[0]};
    Full_Adder FA_10755(s10755, c10755, in10755_1, in10755_2, c8270);
    wire[0:0] s10756, in10756_1, in10756_2;
    wire c10756;
    assign in10756_1 = {s8274[0]};
    assign in10756_2 = {s8275[0]};
    Full_Adder FA_10756(s10756, c10756, in10756_1, in10756_2, s8273[0]);
    wire[0:0] s10757, in10757_1, in10757_2;
    wire c10757;
    assign in10757_1 = {s8277[0]};
    assign in10757_2 = {s8278[0]};
    Full_Adder FA_10757(s10757, c10757, in10757_1, in10757_2, s8276[0]);
    wire[0:0] s10758, in10758_1, in10758_2;
    wire c10758;
    assign in10758_1 = {s8280[0]};
    assign in10758_2 = {s8281[0]};
    Full_Adder FA_10758(s10758, c10758, in10758_1, in10758_2, s8279[0]);
    wire[0:0] s10759, in10759_1, in10759_2;
    wire c10759;
    assign in10759_1 = {c8272};
    assign in10759_2 = {c8273};
    Full_Adder FA_10759(s10759, c10759, in10759_1, in10759_2, c8271);
    wire[0:0] s10760, in10760_1, in10760_2;
    wire c10760;
    assign in10760_1 = {c8275};
    assign in10760_2 = {c8276};
    Full_Adder FA_10760(s10760, c10760, in10760_1, in10760_2, c8274);
    wire[0:0] s10761, in10761_1, in10761_2;
    wire c10761;
    assign in10761_1 = {c8278};
    assign in10761_2 = {c8279};
    Full_Adder FA_10761(s10761, c10761, in10761_1, in10761_2, c8277);
    wire[0:0] s10762, in10762_1, in10762_2;
    wire c10762;
    assign in10762_1 = {c8281};
    assign in10762_2 = {c8282};
    Full_Adder FA_10762(s10762, c10762, in10762_1, in10762_2, c8280);
    wire[0:0] s10763, in10763_1, in10763_2;
    wire c10763;
    assign in10763_1 = {s8284[0]};
    assign in10763_2 = {s8285[0]};
    Full_Adder FA_10763(s10763, c10763, in10763_1, in10763_2, c8283);
    wire[0:0] s10764, in10764_1, in10764_2;
    wire c10764;
    assign in10764_1 = {s8287[0]};
    assign in10764_2 = {s8288[0]};
    Full_Adder FA_10764(s10764, c10764, in10764_1, in10764_2, s8286[0]);
    wire[0:0] s10765, in10765_1, in10765_2;
    wire c10765;
    assign in10765_1 = {s8290[0]};
    assign in10765_2 = {s8291[0]};
    Full_Adder FA_10765(s10765, c10765, in10765_1, in10765_2, s8289[0]);
    wire[0:0] s10766, in10766_1, in10766_2;
    wire c10766;
    assign in10766_1 = {s8293[0]};
    assign in10766_2 = {s8294[0]};
    Full_Adder FA_10766(s10766, c10766, in10766_1, in10766_2, s8292[0]);
    wire[0:0] s10767, in10767_1, in10767_2;
    wire c10767;
    assign in10767_1 = {c8285};
    assign in10767_2 = {c8286};
    Full_Adder FA_10767(s10767, c10767, in10767_1, in10767_2, c8284);
    wire[0:0] s10768, in10768_1, in10768_2;
    wire c10768;
    assign in10768_1 = {c8288};
    assign in10768_2 = {c8289};
    Full_Adder FA_10768(s10768, c10768, in10768_1, in10768_2, c8287);
    wire[0:0] s10769, in10769_1, in10769_2;
    wire c10769;
    assign in10769_1 = {c8291};
    assign in10769_2 = {c8292};
    Full_Adder FA_10769(s10769, c10769, in10769_1, in10769_2, c8290);
    wire[0:0] s10770, in10770_1, in10770_2;
    wire c10770;
    assign in10770_1 = {c8294};
    assign in10770_2 = {c8295};
    Full_Adder FA_10770(s10770, c10770, in10770_1, in10770_2, c8293);
    wire[0:0] s10771, in10771_1, in10771_2;
    wire c10771;
    assign in10771_1 = {s8297[0]};
    assign in10771_2 = {s8298[0]};
    Full_Adder FA_10771(s10771, c10771, in10771_1, in10771_2, c8296);
    wire[0:0] s10772, in10772_1, in10772_2;
    wire c10772;
    assign in10772_1 = {s8300[0]};
    assign in10772_2 = {s8301[0]};
    Full_Adder FA_10772(s10772, c10772, in10772_1, in10772_2, s8299[0]);
    wire[0:0] s10773, in10773_1, in10773_2;
    wire c10773;
    assign in10773_1 = {s8303[0]};
    assign in10773_2 = {s8304[0]};
    Full_Adder FA_10773(s10773, c10773, in10773_1, in10773_2, s8302[0]);
    wire[0:0] s10774, in10774_1, in10774_2;
    wire c10774;
    assign in10774_1 = {s8306[0]};
    assign in10774_2 = {s8307[0]};
    Full_Adder FA_10774(s10774, c10774, in10774_1, in10774_2, s8305[0]);
    wire[0:0] s10775, in10775_1, in10775_2;
    wire c10775;
    assign in10775_1 = {c8298};
    assign in10775_2 = {c8299};
    Full_Adder FA_10775(s10775, c10775, in10775_1, in10775_2, c8297);
    wire[0:0] s10776, in10776_1, in10776_2;
    wire c10776;
    assign in10776_1 = {c8301};
    assign in10776_2 = {c8302};
    Full_Adder FA_10776(s10776, c10776, in10776_1, in10776_2, c8300);
    wire[0:0] s10777, in10777_1, in10777_2;
    wire c10777;
    assign in10777_1 = {c8304};
    assign in10777_2 = {c8305};
    Full_Adder FA_10777(s10777, c10777, in10777_1, in10777_2, c8303);
    wire[0:0] s10778, in10778_1, in10778_2;
    wire c10778;
    assign in10778_1 = {c8307};
    assign in10778_2 = {c8308};
    Full_Adder FA_10778(s10778, c10778, in10778_1, in10778_2, c8306);
    wire[0:0] s10779, in10779_1, in10779_2;
    wire c10779;
    assign in10779_1 = {s8310[0]};
    assign in10779_2 = {s8311[0]};
    Full_Adder FA_10779(s10779, c10779, in10779_1, in10779_2, c8309);
    wire[0:0] s10780, in10780_1, in10780_2;
    wire c10780;
    assign in10780_1 = {s8313[0]};
    assign in10780_2 = {s8314[0]};
    Full_Adder FA_10780(s10780, c10780, in10780_1, in10780_2, s8312[0]);
    wire[0:0] s10781, in10781_1, in10781_2;
    wire c10781;
    assign in10781_1 = {s8316[0]};
    assign in10781_2 = {s8317[0]};
    Full_Adder FA_10781(s10781, c10781, in10781_1, in10781_2, s8315[0]);
    wire[0:0] s10782, in10782_1, in10782_2;
    wire c10782;
    assign in10782_1 = {s8319[0]};
    assign in10782_2 = {s8320[0]};
    Full_Adder FA_10782(s10782, c10782, in10782_1, in10782_2, s8318[0]);
    wire[0:0] s10783, in10783_1, in10783_2;
    wire c10783;
    assign in10783_1 = {c8311};
    assign in10783_2 = {c8312};
    Full_Adder FA_10783(s10783, c10783, in10783_1, in10783_2, c8310);
    wire[0:0] s10784, in10784_1, in10784_2;
    wire c10784;
    assign in10784_1 = {c8314};
    assign in10784_2 = {c8315};
    Full_Adder FA_10784(s10784, c10784, in10784_1, in10784_2, c8313);
    wire[0:0] s10785, in10785_1, in10785_2;
    wire c10785;
    assign in10785_1 = {c8317};
    assign in10785_2 = {c8318};
    Full_Adder FA_10785(s10785, c10785, in10785_1, in10785_2, c8316);
    wire[0:0] s10786, in10786_1, in10786_2;
    wire c10786;
    assign in10786_1 = {c8320};
    assign in10786_2 = {c8321};
    Full_Adder FA_10786(s10786, c10786, in10786_1, in10786_2, c8319);
    wire[0:0] s10787, in10787_1, in10787_2;
    wire c10787;
    assign in10787_1 = {s8323[0]};
    assign in10787_2 = {s8324[0]};
    Full_Adder FA_10787(s10787, c10787, in10787_1, in10787_2, c8322);
    wire[0:0] s10788, in10788_1, in10788_2;
    wire c10788;
    assign in10788_1 = {s8326[0]};
    assign in10788_2 = {s8327[0]};
    Full_Adder FA_10788(s10788, c10788, in10788_1, in10788_2, s8325[0]);
    wire[0:0] s10789, in10789_1, in10789_2;
    wire c10789;
    assign in10789_1 = {s8329[0]};
    assign in10789_2 = {s8330[0]};
    Full_Adder FA_10789(s10789, c10789, in10789_1, in10789_2, s8328[0]);
    wire[0:0] s10790, in10790_1, in10790_2;
    wire c10790;
    assign in10790_1 = {s8332[0]};
    assign in10790_2 = {s8333[0]};
    Full_Adder FA_10790(s10790, c10790, in10790_1, in10790_2, s8331[0]);
    wire[0:0] s10791, in10791_1, in10791_2;
    wire c10791;
    assign in10791_1 = {c8324};
    assign in10791_2 = {c8325};
    Full_Adder FA_10791(s10791, c10791, in10791_1, in10791_2, c8323);
    wire[0:0] s10792, in10792_1, in10792_2;
    wire c10792;
    assign in10792_1 = {c8327};
    assign in10792_2 = {c8328};
    Full_Adder FA_10792(s10792, c10792, in10792_1, in10792_2, c8326);
    wire[0:0] s10793, in10793_1, in10793_2;
    wire c10793;
    assign in10793_1 = {c8330};
    assign in10793_2 = {c8331};
    Full_Adder FA_10793(s10793, c10793, in10793_1, in10793_2, c8329);
    wire[0:0] s10794, in10794_1, in10794_2;
    wire c10794;
    assign in10794_1 = {c8333};
    assign in10794_2 = {c8334};
    Full_Adder FA_10794(s10794, c10794, in10794_1, in10794_2, c8332);
    wire[0:0] s10795, in10795_1, in10795_2;
    wire c10795;
    assign in10795_1 = {s8336[0]};
    assign in10795_2 = {s8337[0]};
    Full_Adder FA_10795(s10795, c10795, in10795_1, in10795_2, c8335);
    wire[0:0] s10796, in10796_1, in10796_2;
    wire c10796;
    assign in10796_1 = {s8339[0]};
    assign in10796_2 = {s8340[0]};
    Full_Adder FA_10796(s10796, c10796, in10796_1, in10796_2, s8338[0]);
    wire[0:0] s10797, in10797_1, in10797_2;
    wire c10797;
    assign in10797_1 = {s8342[0]};
    assign in10797_2 = {s8343[0]};
    Full_Adder FA_10797(s10797, c10797, in10797_1, in10797_2, s8341[0]);
    wire[0:0] s10798, in10798_1, in10798_2;
    wire c10798;
    assign in10798_1 = {s8345[0]};
    assign in10798_2 = {s8346[0]};
    Full_Adder FA_10798(s10798, c10798, in10798_1, in10798_2, s8344[0]);
    wire[0:0] s10799, in10799_1, in10799_2;
    wire c10799;
    assign in10799_1 = {c8337};
    assign in10799_2 = {c8338};
    Full_Adder FA_10799(s10799, c10799, in10799_1, in10799_2, c8336);
    wire[0:0] s10800, in10800_1, in10800_2;
    wire c10800;
    assign in10800_1 = {c8340};
    assign in10800_2 = {c8341};
    Full_Adder FA_10800(s10800, c10800, in10800_1, in10800_2, c8339);
    wire[0:0] s10801, in10801_1, in10801_2;
    wire c10801;
    assign in10801_1 = {c8343};
    assign in10801_2 = {c8344};
    Full_Adder FA_10801(s10801, c10801, in10801_1, in10801_2, c8342);
    wire[0:0] s10802, in10802_1, in10802_2;
    wire c10802;
    assign in10802_1 = {c8346};
    assign in10802_2 = {c8347};
    Full_Adder FA_10802(s10802, c10802, in10802_1, in10802_2, c8345);
    wire[0:0] s10803, in10803_1, in10803_2;
    wire c10803;
    assign in10803_1 = {s8349[0]};
    assign in10803_2 = {s8350[0]};
    Full_Adder FA_10803(s10803, c10803, in10803_1, in10803_2, c8348);
    wire[0:0] s10804, in10804_1, in10804_2;
    wire c10804;
    assign in10804_1 = {s8352[0]};
    assign in10804_2 = {s8353[0]};
    Full_Adder FA_10804(s10804, c10804, in10804_1, in10804_2, s8351[0]);
    wire[0:0] s10805, in10805_1, in10805_2;
    wire c10805;
    assign in10805_1 = {s8355[0]};
    assign in10805_2 = {s8356[0]};
    Full_Adder FA_10805(s10805, c10805, in10805_1, in10805_2, s8354[0]);
    wire[0:0] s10806, in10806_1, in10806_2;
    wire c10806;
    assign in10806_1 = {s8358[0]};
    assign in10806_2 = {s8359[0]};
    Full_Adder FA_10806(s10806, c10806, in10806_1, in10806_2, s8357[0]);
    wire[0:0] s10807, in10807_1, in10807_2;
    wire c10807;
    assign in10807_1 = {c8350};
    assign in10807_2 = {c8351};
    Full_Adder FA_10807(s10807, c10807, in10807_1, in10807_2, c8349);
    wire[0:0] s10808, in10808_1, in10808_2;
    wire c10808;
    assign in10808_1 = {c8353};
    assign in10808_2 = {c8354};
    Full_Adder FA_10808(s10808, c10808, in10808_1, in10808_2, c8352);
    wire[0:0] s10809, in10809_1, in10809_2;
    wire c10809;
    assign in10809_1 = {c8356};
    assign in10809_2 = {c8357};
    Full_Adder FA_10809(s10809, c10809, in10809_1, in10809_2, c8355);
    wire[0:0] s10810, in10810_1, in10810_2;
    wire c10810;
    assign in10810_1 = {c8359};
    assign in10810_2 = {c8360};
    Full_Adder FA_10810(s10810, c10810, in10810_1, in10810_2, c8358);
    wire[0:0] s10811, in10811_1, in10811_2;
    wire c10811;
    assign in10811_1 = {s8362[0]};
    assign in10811_2 = {s8363[0]};
    Full_Adder FA_10811(s10811, c10811, in10811_1, in10811_2, c8361);
    wire[0:0] s10812, in10812_1, in10812_2;
    wire c10812;
    assign in10812_1 = {s8365[0]};
    assign in10812_2 = {s8366[0]};
    Full_Adder FA_10812(s10812, c10812, in10812_1, in10812_2, s8364[0]);
    wire[0:0] s10813, in10813_1, in10813_2;
    wire c10813;
    assign in10813_1 = {s8368[0]};
    assign in10813_2 = {s8369[0]};
    Full_Adder FA_10813(s10813, c10813, in10813_1, in10813_2, s8367[0]);
    wire[0:0] s10814, in10814_1, in10814_2;
    wire c10814;
    assign in10814_1 = {s8371[0]};
    assign in10814_2 = {s8372[0]};
    Full_Adder FA_10814(s10814, c10814, in10814_1, in10814_2, s8370[0]);
    wire[0:0] s10815, in10815_1, in10815_2;
    wire c10815;
    assign in10815_1 = {c8363};
    assign in10815_2 = {c8364};
    Full_Adder FA_10815(s10815, c10815, in10815_1, in10815_2, c8362);
    wire[0:0] s10816, in10816_1, in10816_2;
    wire c10816;
    assign in10816_1 = {c8366};
    assign in10816_2 = {c8367};
    Full_Adder FA_10816(s10816, c10816, in10816_1, in10816_2, c8365);
    wire[0:0] s10817, in10817_1, in10817_2;
    wire c10817;
    assign in10817_1 = {c8369};
    assign in10817_2 = {c8370};
    Full_Adder FA_10817(s10817, c10817, in10817_1, in10817_2, c8368);
    wire[0:0] s10818, in10818_1, in10818_2;
    wire c10818;
    assign in10818_1 = {c8372};
    assign in10818_2 = {c8373};
    Full_Adder FA_10818(s10818, c10818, in10818_1, in10818_2, c8371);
    wire[0:0] s10819, in10819_1, in10819_2;
    wire c10819;
    assign in10819_1 = {s8375[0]};
    assign in10819_2 = {s8376[0]};
    Full_Adder FA_10819(s10819, c10819, in10819_1, in10819_2, c8374);
    wire[0:0] s10820, in10820_1, in10820_2;
    wire c10820;
    assign in10820_1 = {s8378[0]};
    assign in10820_2 = {s8379[0]};
    Full_Adder FA_10820(s10820, c10820, in10820_1, in10820_2, s8377[0]);
    wire[0:0] s10821, in10821_1, in10821_2;
    wire c10821;
    assign in10821_1 = {s8381[0]};
    assign in10821_2 = {s8382[0]};
    Full_Adder FA_10821(s10821, c10821, in10821_1, in10821_2, s8380[0]);
    wire[0:0] s10822, in10822_1, in10822_2;
    wire c10822;
    assign in10822_1 = {s8384[0]};
    assign in10822_2 = {s8385[0]};
    Full_Adder FA_10822(s10822, c10822, in10822_1, in10822_2, s8383[0]);
    wire[0:0] s10823, in10823_1, in10823_2;
    wire c10823;
    assign in10823_1 = {c8376};
    assign in10823_2 = {c8377};
    Full_Adder FA_10823(s10823, c10823, in10823_1, in10823_2, c8375);
    wire[0:0] s10824, in10824_1, in10824_2;
    wire c10824;
    assign in10824_1 = {c8379};
    assign in10824_2 = {c8380};
    Full_Adder FA_10824(s10824, c10824, in10824_1, in10824_2, c8378);
    wire[0:0] s10825, in10825_1, in10825_2;
    wire c10825;
    assign in10825_1 = {c8382};
    assign in10825_2 = {c8383};
    Full_Adder FA_10825(s10825, c10825, in10825_1, in10825_2, c8381);
    wire[0:0] s10826, in10826_1, in10826_2;
    wire c10826;
    assign in10826_1 = {c8385};
    assign in10826_2 = {c8386};
    Full_Adder FA_10826(s10826, c10826, in10826_1, in10826_2, c8384);
    wire[0:0] s10827, in10827_1, in10827_2;
    wire c10827;
    assign in10827_1 = {s8388[0]};
    assign in10827_2 = {s8389[0]};
    Full_Adder FA_10827(s10827, c10827, in10827_1, in10827_2, c8387);
    wire[0:0] s10828, in10828_1, in10828_2;
    wire c10828;
    assign in10828_1 = {s8391[0]};
    assign in10828_2 = {s8392[0]};
    Full_Adder FA_10828(s10828, c10828, in10828_1, in10828_2, s8390[0]);
    wire[0:0] s10829, in10829_1, in10829_2;
    wire c10829;
    assign in10829_1 = {s8394[0]};
    assign in10829_2 = {s8395[0]};
    Full_Adder FA_10829(s10829, c10829, in10829_1, in10829_2, s8393[0]);
    wire[0:0] s10830, in10830_1, in10830_2;
    wire c10830;
    assign in10830_1 = {s8397[0]};
    assign in10830_2 = {s8398[0]};
    Full_Adder FA_10830(s10830, c10830, in10830_1, in10830_2, s8396[0]);
    wire[0:0] s10831, in10831_1, in10831_2;
    wire c10831;
    assign in10831_1 = {c8389};
    assign in10831_2 = {c8390};
    Full_Adder FA_10831(s10831, c10831, in10831_1, in10831_2, c8388);
    wire[0:0] s10832, in10832_1, in10832_2;
    wire c10832;
    assign in10832_1 = {c8392};
    assign in10832_2 = {c8393};
    Full_Adder FA_10832(s10832, c10832, in10832_1, in10832_2, c8391);
    wire[0:0] s10833, in10833_1, in10833_2;
    wire c10833;
    assign in10833_1 = {c8395};
    assign in10833_2 = {c8396};
    Full_Adder FA_10833(s10833, c10833, in10833_1, in10833_2, c8394);
    wire[0:0] s10834, in10834_1, in10834_2;
    wire c10834;
    assign in10834_1 = {c8398};
    assign in10834_2 = {c8399};
    Full_Adder FA_10834(s10834, c10834, in10834_1, in10834_2, c8397);
    wire[0:0] s10835, in10835_1, in10835_2;
    wire c10835;
    assign in10835_1 = {s8401[0]};
    assign in10835_2 = {s8402[0]};
    Full_Adder FA_10835(s10835, c10835, in10835_1, in10835_2, c8400);
    wire[0:0] s10836, in10836_1, in10836_2;
    wire c10836;
    assign in10836_1 = {s8404[0]};
    assign in10836_2 = {s8405[0]};
    Full_Adder FA_10836(s10836, c10836, in10836_1, in10836_2, s8403[0]);
    wire[0:0] s10837, in10837_1, in10837_2;
    wire c10837;
    assign in10837_1 = {s8407[0]};
    assign in10837_2 = {s8408[0]};
    Full_Adder FA_10837(s10837, c10837, in10837_1, in10837_2, s8406[0]);
    wire[0:0] s10838, in10838_1, in10838_2;
    wire c10838;
    assign in10838_1 = {s8410[0]};
    assign in10838_2 = {s8411[0]};
    Full_Adder FA_10838(s10838, c10838, in10838_1, in10838_2, s8409[0]);
    wire[0:0] s10839, in10839_1, in10839_2;
    wire c10839;
    assign in10839_1 = {c8402};
    assign in10839_2 = {c8403};
    Full_Adder FA_10839(s10839, c10839, in10839_1, in10839_2, c8401);
    wire[0:0] s10840, in10840_1, in10840_2;
    wire c10840;
    assign in10840_1 = {c8405};
    assign in10840_2 = {c8406};
    Full_Adder FA_10840(s10840, c10840, in10840_1, in10840_2, c8404);
    wire[0:0] s10841, in10841_1, in10841_2;
    wire c10841;
    assign in10841_1 = {c8408};
    assign in10841_2 = {c8409};
    Full_Adder FA_10841(s10841, c10841, in10841_1, in10841_2, c8407);
    wire[0:0] s10842, in10842_1, in10842_2;
    wire c10842;
    assign in10842_1 = {c8411};
    assign in10842_2 = {c8412};
    Full_Adder FA_10842(s10842, c10842, in10842_1, in10842_2, c8410);
    wire[0:0] s10843, in10843_1, in10843_2;
    wire c10843;
    assign in10843_1 = {s8414[0]};
    assign in10843_2 = {s8415[0]};
    Full_Adder FA_10843(s10843, c10843, in10843_1, in10843_2, c8413);
    wire[0:0] s10844, in10844_1, in10844_2;
    wire c10844;
    assign in10844_1 = {s8417[0]};
    assign in10844_2 = {s8418[0]};
    Full_Adder FA_10844(s10844, c10844, in10844_1, in10844_2, s8416[0]);
    wire[0:0] s10845, in10845_1, in10845_2;
    wire c10845;
    assign in10845_1 = {s8420[0]};
    assign in10845_2 = {s8421[0]};
    Full_Adder FA_10845(s10845, c10845, in10845_1, in10845_2, s8419[0]);
    wire[0:0] s10846, in10846_1, in10846_2;
    wire c10846;
    assign in10846_1 = {s8423[0]};
    assign in10846_2 = {s8424[0]};
    Full_Adder FA_10846(s10846, c10846, in10846_1, in10846_2, s8422[0]);
    wire[0:0] s10847, in10847_1, in10847_2;
    wire c10847;
    assign in10847_1 = {c8415};
    assign in10847_2 = {c8416};
    Full_Adder FA_10847(s10847, c10847, in10847_1, in10847_2, c8414);
    wire[0:0] s10848, in10848_1, in10848_2;
    wire c10848;
    assign in10848_1 = {c8418};
    assign in10848_2 = {c8419};
    Full_Adder FA_10848(s10848, c10848, in10848_1, in10848_2, c8417);
    wire[0:0] s10849, in10849_1, in10849_2;
    wire c10849;
    assign in10849_1 = {c8421};
    assign in10849_2 = {c8422};
    Full_Adder FA_10849(s10849, c10849, in10849_1, in10849_2, c8420);
    wire[0:0] s10850, in10850_1, in10850_2;
    wire c10850;
    assign in10850_1 = {c8424};
    assign in10850_2 = {c8425};
    Full_Adder FA_10850(s10850, c10850, in10850_1, in10850_2, c8423);
    wire[0:0] s10851, in10851_1, in10851_2;
    wire c10851;
    assign in10851_1 = {s8427[0]};
    assign in10851_2 = {s8428[0]};
    Full_Adder FA_10851(s10851, c10851, in10851_1, in10851_2, c8426);
    wire[0:0] s10852, in10852_1, in10852_2;
    wire c10852;
    assign in10852_1 = {s8430[0]};
    assign in10852_2 = {s8431[0]};
    Full_Adder FA_10852(s10852, c10852, in10852_1, in10852_2, s8429[0]);
    wire[0:0] s10853, in10853_1, in10853_2;
    wire c10853;
    assign in10853_1 = {s8433[0]};
    assign in10853_2 = {s8434[0]};
    Full_Adder FA_10853(s10853, c10853, in10853_1, in10853_2, s8432[0]);
    wire[0:0] s10854, in10854_1, in10854_2;
    wire c10854;
    assign in10854_1 = {s8436[0]};
    assign in10854_2 = {s8437[0]};
    Full_Adder FA_10854(s10854, c10854, in10854_1, in10854_2, s8435[0]);
    wire[0:0] s10855, in10855_1, in10855_2;
    wire c10855;
    assign in10855_1 = {c8428};
    assign in10855_2 = {c8429};
    Full_Adder FA_10855(s10855, c10855, in10855_1, in10855_2, c8427);
    wire[0:0] s10856, in10856_1, in10856_2;
    wire c10856;
    assign in10856_1 = {c8431};
    assign in10856_2 = {c8432};
    Full_Adder FA_10856(s10856, c10856, in10856_1, in10856_2, c8430);
    wire[0:0] s10857, in10857_1, in10857_2;
    wire c10857;
    assign in10857_1 = {c8434};
    assign in10857_2 = {c8435};
    Full_Adder FA_10857(s10857, c10857, in10857_1, in10857_2, c8433);
    wire[0:0] s10858, in10858_1, in10858_2;
    wire c10858;
    assign in10858_1 = {c8437};
    assign in10858_2 = {c8438};
    Full_Adder FA_10858(s10858, c10858, in10858_1, in10858_2, c8436);
    wire[0:0] s10859, in10859_1, in10859_2;
    wire c10859;
    assign in10859_1 = {s8440[0]};
    assign in10859_2 = {s8441[0]};
    Full_Adder FA_10859(s10859, c10859, in10859_1, in10859_2, c8439);
    wire[0:0] s10860, in10860_1, in10860_2;
    wire c10860;
    assign in10860_1 = {s8443[0]};
    assign in10860_2 = {s8444[0]};
    Full_Adder FA_10860(s10860, c10860, in10860_1, in10860_2, s8442[0]);
    wire[0:0] s10861, in10861_1, in10861_2;
    wire c10861;
    assign in10861_1 = {s8446[0]};
    assign in10861_2 = {s8447[0]};
    Full_Adder FA_10861(s10861, c10861, in10861_1, in10861_2, s8445[0]);
    wire[0:0] s10862, in10862_1, in10862_2;
    wire c10862;
    assign in10862_1 = {s8449[0]};
    assign in10862_2 = {s8450[0]};
    Full_Adder FA_10862(s10862, c10862, in10862_1, in10862_2, s8448[0]);
    wire[0:0] s10863, in10863_1, in10863_2;
    wire c10863;
    assign in10863_1 = {c8441};
    assign in10863_2 = {c8442};
    Full_Adder FA_10863(s10863, c10863, in10863_1, in10863_2, c8440);
    wire[0:0] s10864, in10864_1, in10864_2;
    wire c10864;
    assign in10864_1 = {c8444};
    assign in10864_2 = {c8445};
    Full_Adder FA_10864(s10864, c10864, in10864_1, in10864_2, c8443);
    wire[0:0] s10865, in10865_1, in10865_2;
    wire c10865;
    assign in10865_1 = {c8447};
    assign in10865_2 = {c8448};
    Full_Adder FA_10865(s10865, c10865, in10865_1, in10865_2, c8446);
    wire[0:0] s10866, in10866_1, in10866_2;
    wire c10866;
    assign in10866_1 = {c8450};
    assign in10866_2 = {c8451};
    Full_Adder FA_10866(s10866, c10866, in10866_1, in10866_2, c8449);
    wire[0:0] s10867, in10867_1, in10867_2;
    wire c10867;
    assign in10867_1 = {s8453[0]};
    assign in10867_2 = {s8454[0]};
    Full_Adder FA_10867(s10867, c10867, in10867_1, in10867_2, c8452);
    wire[0:0] s10868, in10868_1, in10868_2;
    wire c10868;
    assign in10868_1 = {s8456[0]};
    assign in10868_2 = {s8457[0]};
    Full_Adder FA_10868(s10868, c10868, in10868_1, in10868_2, s8455[0]);
    wire[0:0] s10869, in10869_1, in10869_2;
    wire c10869;
    assign in10869_1 = {s8459[0]};
    assign in10869_2 = {s8460[0]};
    Full_Adder FA_10869(s10869, c10869, in10869_1, in10869_2, s8458[0]);
    wire[0:0] s10870, in10870_1, in10870_2;
    wire c10870;
    assign in10870_1 = {s8462[0]};
    assign in10870_2 = {s8463[0]};
    Full_Adder FA_10870(s10870, c10870, in10870_1, in10870_2, s8461[0]);
    wire[0:0] s10871, in10871_1, in10871_2;
    wire c10871;
    assign in10871_1 = {c8454};
    assign in10871_2 = {c8455};
    Full_Adder FA_10871(s10871, c10871, in10871_1, in10871_2, c8453);
    wire[0:0] s10872, in10872_1, in10872_2;
    wire c10872;
    assign in10872_1 = {c8457};
    assign in10872_2 = {c8458};
    Full_Adder FA_10872(s10872, c10872, in10872_1, in10872_2, c8456);
    wire[0:0] s10873, in10873_1, in10873_2;
    wire c10873;
    assign in10873_1 = {c8460};
    assign in10873_2 = {c8461};
    Full_Adder FA_10873(s10873, c10873, in10873_1, in10873_2, c8459);
    wire[0:0] s10874, in10874_1, in10874_2;
    wire c10874;
    assign in10874_1 = {c8463};
    assign in10874_2 = {c8464};
    Full_Adder FA_10874(s10874, c10874, in10874_1, in10874_2, c8462);
    wire[0:0] s10875, in10875_1, in10875_2;
    wire c10875;
    assign in10875_1 = {s8466[0]};
    assign in10875_2 = {s8467[0]};
    Full_Adder FA_10875(s10875, c10875, in10875_1, in10875_2, c8465);
    wire[0:0] s10876, in10876_1, in10876_2;
    wire c10876;
    assign in10876_1 = {s8469[0]};
    assign in10876_2 = {s8470[0]};
    Full_Adder FA_10876(s10876, c10876, in10876_1, in10876_2, s8468[0]);
    wire[0:0] s10877, in10877_1, in10877_2;
    wire c10877;
    assign in10877_1 = {s8472[0]};
    assign in10877_2 = {s8473[0]};
    Full_Adder FA_10877(s10877, c10877, in10877_1, in10877_2, s8471[0]);
    wire[0:0] s10878, in10878_1, in10878_2;
    wire c10878;
    assign in10878_1 = {s8475[0]};
    assign in10878_2 = {s8476[0]};
    Full_Adder FA_10878(s10878, c10878, in10878_1, in10878_2, s8474[0]);
    wire[0:0] s10879, in10879_1, in10879_2;
    wire c10879;
    assign in10879_1 = {c8467};
    assign in10879_2 = {c8468};
    Full_Adder FA_10879(s10879, c10879, in10879_1, in10879_2, c8466);
    wire[0:0] s10880, in10880_1, in10880_2;
    wire c10880;
    assign in10880_1 = {c8470};
    assign in10880_2 = {c8471};
    Full_Adder FA_10880(s10880, c10880, in10880_1, in10880_2, c8469);
    wire[0:0] s10881, in10881_1, in10881_2;
    wire c10881;
    assign in10881_1 = {c8473};
    assign in10881_2 = {c8474};
    Full_Adder FA_10881(s10881, c10881, in10881_1, in10881_2, c8472);
    wire[0:0] s10882, in10882_1, in10882_2;
    wire c10882;
    assign in10882_1 = {c8476};
    assign in10882_2 = {c8477};
    Full_Adder FA_10882(s10882, c10882, in10882_1, in10882_2, c8475);
    wire[0:0] s10883, in10883_1, in10883_2;
    wire c10883;
    assign in10883_1 = {s8479[0]};
    assign in10883_2 = {s8480[0]};
    Full_Adder FA_10883(s10883, c10883, in10883_1, in10883_2, c8478);
    wire[0:0] s10884, in10884_1, in10884_2;
    wire c10884;
    assign in10884_1 = {s8482[0]};
    assign in10884_2 = {s8483[0]};
    Full_Adder FA_10884(s10884, c10884, in10884_1, in10884_2, s8481[0]);
    wire[0:0] s10885, in10885_1, in10885_2;
    wire c10885;
    assign in10885_1 = {s8485[0]};
    assign in10885_2 = {s8486[0]};
    Full_Adder FA_10885(s10885, c10885, in10885_1, in10885_2, s8484[0]);
    wire[0:0] s10886, in10886_1, in10886_2;
    wire c10886;
    assign in10886_1 = {s8488[0]};
    assign in10886_2 = {s8489[0]};
    Full_Adder FA_10886(s10886, c10886, in10886_1, in10886_2, s8487[0]);
    wire[0:0] s10887, in10887_1, in10887_2;
    wire c10887;
    assign in10887_1 = {c8480};
    assign in10887_2 = {c8481};
    Full_Adder FA_10887(s10887, c10887, in10887_1, in10887_2, c8479);
    wire[0:0] s10888, in10888_1, in10888_2;
    wire c10888;
    assign in10888_1 = {c8483};
    assign in10888_2 = {c8484};
    Full_Adder FA_10888(s10888, c10888, in10888_1, in10888_2, c8482);
    wire[0:0] s10889, in10889_1, in10889_2;
    wire c10889;
    assign in10889_1 = {c8486};
    assign in10889_2 = {c8487};
    Full_Adder FA_10889(s10889, c10889, in10889_1, in10889_2, c8485);
    wire[0:0] s10890, in10890_1, in10890_2;
    wire c10890;
    assign in10890_1 = {c8489};
    assign in10890_2 = {c8490};
    Full_Adder FA_10890(s10890, c10890, in10890_1, in10890_2, c8488);
    wire[0:0] s10891, in10891_1, in10891_2;
    wire c10891;
    assign in10891_1 = {s8492[0]};
    assign in10891_2 = {s8493[0]};
    Full_Adder FA_10891(s10891, c10891, in10891_1, in10891_2, c8491);
    wire[0:0] s10892, in10892_1, in10892_2;
    wire c10892;
    assign in10892_1 = {s8495[0]};
    assign in10892_2 = {s8496[0]};
    Full_Adder FA_10892(s10892, c10892, in10892_1, in10892_2, s8494[0]);
    wire[0:0] s10893, in10893_1, in10893_2;
    wire c10893;
    assign in10893_1 = {s8498[0]};
    assign in10893_2 = {s8499[0]};
    Full_Adder FA_10893(s10893, c10893, in10893_1, in10893_2, s8497[0]);
    wire[0:0] s10894, in10894_1, in10894_2;
    wire c10894;
    assign in10894_1 = {s8501[0]};
    assign in10894_2 = {s8502[0]};
    Full_Adder FA_10894(s10894, c10894, in10894_1, in10894_2, s8500[0]);
    wire[0:0] s10895, in10895_1, in10895_2;
    wire c10895;
    assign in10895_1 = {c8493};
    assign in10895_2 = {c8494};
    Full_Adder FA_10895(s10895, c10895, in10895_1, in10895_2, c8492);
    wire[0:0] s10896, in10896_1, in10896_2;
    wire c10896;
    assign in10896_1 = {c8496};
    assign in10896_2 = {c8497};
    Full_Adder FA_10896(s10896, c10896, in10896_1, in10896_2, c8495);
    wire[0:0] s10897, in10897_1, in10897_2;
    wire c10897;
    assign in10897_1 = {c8499};
    assign in10897_2 = {c8500};
    Full_Adder FA_10897(s10897, c10897, in10897_1, in10897_2, c8498);
    wire[0:0] s10898, in10898_1, in10898_2;
    wire c10898;
    assign in10898_1 = {c8502};
    assign in10898_2 = {c8503};
    Full_Adder FA_10898(s10898, c10898, in10898_1, in10898_2, c8501);
    wire[0:0] s10899, in10899_1, in10899_2;
    wire c10899;
    assign in10899_1 = {s8505[0]};
    assign in10899_2 = {s8506[0]};
    Full_Adder FA_10899(s10899, c10899, in10899_1, in10899_2, c8504);
    wire[0:0] s10900, in10900_1, in10900_2;
    wire c10900;
    assign in10900_1 = {s8508[0]};
    assign in10900_2 = {s8509[0]};
    Full_Adder FA_10900(s10900, c10900, in10900_1, in10900_2, s8507[0]);
    wire[0:0] s10901, in10901_1, in10901_2;
    wire c10901;
    assign in10901_1 = {s8511[0]};
    assign in10901_2 = {s8512[0]};
    Full_Adder FA_10901(s10901, c10901, in10901_1, in10901_2, s8510[0]);
    wire[0:0] s10902, in10902_1, in10902_2;
    wire c10902;
    assign in10902_1 = {s8514[0]};
    assign in10902_2 = {s8515[0]};
    Full_Adder FA_10902(s10902, c10902, in10902_1, in10902_2, s8513[0]);
    wire[0:0] s10903, in10903_1, in10903_2;
    wire c10903;
    assign in10903_1 = {c8506};
    assign in10903_2 = {c8507};
    Full_Adder FA_10903(s10903, c10903, in10903_1, in10903_2, c8505);
    wire[0:0] s10904, in10904_1, in10904_2;
    wire c10904;
    assign in10904_1 = {c8509};
    assign in10904_2 = {c8510};
    Full_Adder FA_10904(s10904, c10904, in10904_1, in10904_2, c8508);
    wire[0:0] s10905, in10905_1, in10905_2;
    wire c10905;
    assign in10905_1 = {c8512};
    assign in10905_2 = {c8513};
    Full_Adder FA_10905(s10905, c10905, in10905_1, in10905_2, c8511);
    wire[0:0] s10906, in10906_1, in10906_2;
    wire c10906;
    assign in10906_1 = {c8515};
    assign in10906_2 = {c8516};
    Full_Adder FA_10906(s10906, c10906, in10906_1, in10906_2, c8514);
    wire[0:0] s10907, in10907_1, in10907_2;
    wire c10907;
    assign in10907_1 = {s8518[0]};
    assign in10907_2 = {s8519[0]};
    Full_Adder FA_10907(s10907, c10907, in10907_1, in10907_2, c8517);
    wire[0:0] s10908, in10908_1, in10908_2;
    wire c10908;
    assign in10908_1 = {s8521[0]};
    assign in10908_2 = {s8522[0]};
    Full_Adder FA_10908(s10908, c10908, in10908_1, in10908_2, s8520[0]);
    wire[0:0] s10909, in10909_1, in10909_2;
    wire c10909;
    assign in10909_1 = {s8524[0]};
    assign in10909_2 = {s8525[0]};
    Full_Adder FA_10909(s10909, c10909, in10909_1, in10909_2, s8523[0]);
    wire[0:0] s10910, in10910_1, in10910_2;
    wire c10910;
    assign in10910_1 = {s8527[0]};
    assign in10910_2 = {s8528[0]};
    Full_Adder FA_10910(s10910, c10910, in10910_1, in10910_2, s8526[0]);
    wire[0:0] s10911, in10911_1, in10911_2;
    wire c10911;
    assign in10911_1 = {c8519};
    assign in10911_2 = {c8520};
    Full_Adder FA_10911(s10911, c10911, in10911_1, in10911_2, c8518);
    wire[0:0] s10912, in10912_1, in10912_2;
    wire c10912;
    assign in10912_1 = {c8522};
    assign in10912_2 = {c8523};
    Full_Adder FA_10912(s10912, c10912, in10912_1, in10912_2, c8521);
    wire[0:0] s10913, in10913_1, in10913_2;
    wire c10913;
    assign in10913_1 = {c8525};
    assign in10913_2 = {c8526};
    Full_Adder FA_10913(s10913, c10913, in10913_1, in10913_2, c8524);
    wire[0:0] s10914, in10914_1, in10914_2;
    wire c10914;
    assign in10914_1 = {c8528};
    assign in10914_2 = {c8529};
    Full_Adder FA_10914(s10914, c10914, in10914_1, in10914_2, c8527);
    wire[0:0] s10915, in10915_1, in10915_2;
    wire c10915;
    assign in10915_1 = {s8531[0]};
    assign in10915_2 = {s8532[0]};
    Full_Adder FA_10915(s10915, c10915, in10915_1, in10915_2, c8530);
    wire[0:0] s10916, in10916_1, in10916_2;
    wire c10916;
    assign in10916_1 = {s8534[0]};
    assign in10916_2 = {s8535[0]};
    Full_Adder FA_10916(s10916, c10916, in10916_1, in10916_2, s8533[0]);
    wire[0:0] s10917, in10917_1, in10917_2;
    wire c10917;
    assign in10917_1 = {s8537[0]};
    assign in10917_2 = {s8538[0]};
    Full_Adder FA_10917(s10917, c10917, in10917_1, in10917_2, s8536[0]);
    wire[0:0] s10918, in10918_1, in10918_2;
    wire c10918;
    assign in10918_1 = {s8540[0]};
    assign in10918_2 = {s8541[0]};
    Full_Adder FA_10918(s10918, c10918, in10918_1, in10918_2, s8539[0]);
    wire[0:0] s10919, in10919_1, in10919_2;
    wire c10919;
    assign in10919_1 = {c8532};
    assign in10919_2 = {c8533};
    Full_Adder FA_10919(s10919, c10919, in10919_1, in10919_2, c8531);
    wire[0:0] s10920, in10920_1, in10920_2;
    wire c10920;
    assign in10920_1 = {c8535};
    assign in10920_2 = {c8536};
    Full_Adder FA_10920(s10920, c10920, in10920_1, in10920_2, c8534);
    wire[0:0] s10921, in10921_1, in10921_2;
    wire c10921;
    assign in10921_1 = {c8538};
    assign in10921_2 = {c8539};
    Full_Adder FA_10921(s10921, c10921, in10921_1, in10921_2, c8537);
    wire[0:0] s10922, in10922_1, in10922_2;
    wire c10922;
    assign in10922_1 = {c8541};
    assign in10922_2 = {c8542};
    Full_Adder FA_10922(s10922, c10922, in10922_1, in10922_2, c8540);
    wire[0:0] s10923, in10923_1, in10923_2;
    wire c10923;
    assign in10923_1 = {s8544[0]};
    assign in10923_2 = {s8545[0]};
    Full_Adder FA_10923(s10923, c10923, in10923_1, in10923_2, c8543);
    wire[0:0] s10924, in10924_1, in10924_2;
    wire c10924;
    assign in10924_1 = {s8547[0]};
    assign in10924_2 = {s8548[0]};
    Full_Adder FA_10924(s10924, c10924, in10924_1, in10924_2, s8546[0]);
    wire[0:0] s10925, in10925_1, in10925_2;
    wire c10925;
    assign in10925_1 = {s8550[0]};
    assign in10925_2 = {s8551[0]};
    Full_Adder FA_10925(s10925, c10925, in10925_1, in10925_2, s8549[0]);
    wire[0:0] s10926, in10926_1, in10926_2;
    wire c10926;
    assign in10926_1 = {s8553[0]};
    assign in10926_2 = {s8554[0]};
    Full_Adder FA_10926(s10926, c10926, in10926_1, in10926_2, s8552[0]);
    wire[0:0] s10927, in10927_1, in10927_2;
    wire c10927;
    assign in10927_1 = {c8545};
    assign in10927_2 = {c8546};
    Full_Adder FA_10927(s10927, c10927, in10927_1, in10927_2, c8544);
    wire[0:0] s10928, in10928_1, in10928_2;
    wire c10928;
    assign in10928_1 = {c8548};
    assign in10928_2 = {c8549};
    Full_Adder FA_10928(s10928, c10928, in10928_1, in10928_2, c8547);
    wire[0:0] s10929, in10929_1, in10929_2;
    wire c10929;
    assign in10929_1 = {c8551};
    assign in10929_2 = {c8552};
    Full_Adder FA_10929(s10929, c10929, in10929_1, in10929_2, c8550);
    wire[0:0] s10930, in10930_1, in10930_2;
    wire c10930;
    assign in10930_1 = {c8554};
    assign in10930_2 = {c8555};
    Full_Adder FA_10930(s10930, c10930, in10930_1, in10930_2, c8553);
    wire[0:0] s10931, in10931_1, in10931_2;
    wire c10931;
    assign in10931_1 = {s8557[0]};
    assign in10931_2 = {s8558[0]};
    Full_Adder FA_10931(s10931, c10931, in10931_1, in10931_2, c8556);
    wire[0:0] s10932, in10932_1, in10932_2;
    wire c10932;
    assign in10932_1 = {s8560[0]};
    assign in10932_2 = {s8561[0]};
    Full_Adder FA_10932(s10932, c10932, in10932_1, in10932_2, s8559[0]);
    wire[0:0] s10933, in10933_1, in10933_2;
    wire c10933;
    assign in10933_1 = {s8563[0]};
    assign in10933_2 = {s8564[0]};
    Full_Adder FA_10933(s10933, c10933, in10933_1, in10933_2, s8562[0]);
    wire[0:0] s10934, in10934_1, in10934_2;
    wire c10934;
    assign in10934_1 = {s8566[0]};
    assign in10934_2 = {s8567[0]};
    Full_Adder FA_10934(s10934, c10934, in10934_1, in10934_2, s8565[0]);
    wire[0:0] s10935, in10935_1, in10935_2;
    wire c10935;
    assign in10935_1 = {c8558};
    assign in10935_2 = {c8559};
    Full_Adder FA_10935(s10935, c10935, in10935_1, in10935_2, c8557);
    wire[0:0] s10936, in10936_1, in10936_2;
    wire c10936;
    assign in10936_1 = {c8561};
    assign in10936_2 = {c8562};
    Full_Adder FA_10936(s10936, c10936, in10936_1, in10936_2, c8560);
    wire[0:0] s10937, in10937_1, in10937_2;
    wire c10937;
    assign in10937_1 = {c8564};
    assign in10937_2 = {c8565};
    Full_Adder FA_10937(s10937, c10937, in10937_1, in10937_2, c8563);
    wire[0:0] s10938, in10938_1, in10938_2;
    wire c10938;
    assign in10938_1 = {c8567};
    assign in10938_2 = {c8568};
    Full_Adder FA_10938(s10938, c10938, in10938_1, in10938_2, c8566);
    wire[0:0] s10939, in10939_1, in10939_2;
    wire c10939;
    assign in10939_1 = {s8570[0]};
    assign in10939_2 = {s8571[0]};
    Full_Adder FA_10939(s10939, c10939, in10939_1, in10939_2, c8569);
    wire[0:0] s10940, in10940_1, in10940_2;
    wire c10940;
    assign in10940_1 = {s8573[0]};
    assign in10940_2 = {s8574[0]};
    Full_Adder FA_10940(s10940, c10940, in10940_1, in10940_2, s8572[0]);
    wire[0:0] s10941, in10941_1, in10941_2;
    wire c10941;
    assign in10941_1 = {s8576[0]};
    assign in10941_2 = {s8577[0]};
    Full_Adder FA_10941(s10941, c10941, in10941_1, in10941_2, s8575[0]);
    wire[0:0] s10942, in10942_1, in10942_2;
    wire c10942;
    assign in10942_1 = {s8579[0]};
    assign in10942_2 = {s8580[0]};
    Full_Adder FA_10942(s10942, c10942, in10942_1, in10942_2, s8578[0]);
    wire[0:0] s10943, in10943_1, in10943_2;
    wire c10943;
    assign in10943_1 = {c8571};
    assign in10943_2 = {c8572};
    Full_Adder FA_10943(s10943, c10943, in10943_1, in10943_2, c8570);
    wire[0:0] s10944, in10944_1, in10944_2;
    wire c10944;
    assign in10944_1 = {c8574};
    assign in10944_2 = {c8575};
    Full_Adder FA_10944(s10944, c10944, in10944_1, in10944_2, c8573);
    wire[0:0] s10945, in10945_1, in10945_2;
    wire c10945;
    assign in10945_1 = {c8577};
    assign in10945_2 = {c8578};
    Full_Adder FA_10945(s10945, c10945, in10945_1, in10945_2, c8576);
    wire[0:0] s10946, in10946_1, in10946_2;
    wire c10946;
    assign in10946_1 = {c8580};
    assign in10946_2 = {c8581};
    Full_Adder FA_10946(s10946, c10946, in10946_1, in10946_2, c8579);
    wire[0:0] s10947, in10947_1, in10947_2;
    wire c10947;
    assign in10947_1 = {s8583[0]};
    assign in10947_2 = {s8584[0]};
    Full_Adder FA_10947(s10947, c10947, in10947_1, in10947_2, c8582);
    wire[0:0] s10948, in10948_1, in10948_2;
    wire c10948;
    assign in10948_1 = {s8586[0]};
    assign in10948_2 = {s8587[0]};
    Full_Adder FA_10948(s10948, c10948, in10948_1, in10948_2, s8585[0]);
    wire[0:0] s10949, in10949_1, in10949_2;
    wire c10949;
    assign in10949_1 = {s8589[0]};
    assign in10949_2 = {s8590[0]};
    Full_Adder FA_10949(s10949, c10949, in10949_1, in10949_2, s8588[0]);
    wire[0:0] s10950, in10950_1, in10950_2;
    wire c10950;
    assign in10950_1 = {s8592[0]};
    assign in10950_2 = {s8593[0]};
    Full_Adder FA_10950(s10950, c10950, in10950_1, in10950_2, s8591[0]);
    wire[0:0] s10951, in10951_1, in10951_2;
    wire c10951;
    assign in10951_1 = {c8584};
    assign in10951_2 = {c8585};
    Full_Adder FA_10951(s10951, c10951, in10951_1, in10951_2, c8583);
    wire[0:0] s10952, in10952_1, in10952_2;
    wire c10952;
    assign in10952_1 = {c8587};
    assign in10952_2 = {c8588};
    Full_Adder FA_10952(s10952, c10952, in10952_1, in10952_2, c8586);
    wire[0:0] s10953, in10953_1, in10953_2;
    wire c10953;
    assign in10953_1 = {c8590};
    assign in10953_2 = {c8591};
    Full_Adder FA_10953(s10953, c10953, in10953_1, in10953_2, c8589);
    wire[0:0] s10954, in10954_1, in10954_2;
    wire c10954;
    assign in10954_1 = {c8593};
    assign in10954_2 = {c8594};
    Full_Adder FA_10954(s10954, c10954, in10954_1, in10954_2, c8592);
    wire[0:0] s10955, in10955_1, in10955_2;
    wire c10955;
    assign in10955_1 = {s8596[0]};
    assign in10955_2 = {s8597[0]};
    Full_Adder FA_10955(s10955, c10955, in10955_1, in10955_2, c8595);
    wire[0:0] s10956, in10956_1, in10956_2;
    wire c10956;
    assign in10956_1 = {s8599[0]};
    assign in10956_2 = {s8600[0]};
    Full_Adder FA_10956(s10956, c10956, in10956_1, in10956_2, s8598[0]);
    wire[0:0] s10957, in10957_1, in10957_2;
    wire c10957;
    assign in10957_1 = {s8602[0]};
    assign in10957_2 = {s8603[0]};
    Full_Adder FA_10957(s10957, c10957, in10957_1, in10957_2, s8601[0]);
    wire[0:0] s10958, in10958_1, in10958_2;
    wire c10958;
    assign in10958_1 = {s8605[0]};
    assign in10958_2 = {s8606[0]};
    Full_Adder FA_10958(s10958, c10958, in10958_1, in10958_2, s8604[0]);
    wire[0:0] s10959, in10959_1, in10959_2;
    wire c10959;
    assign in10959_1 = {c8597};
    assign in10959_2 = {c8598};
    Full_Adder FA_10959(s10959, c10959, in10959_1, in10959_2, c8596);
    wire[0:0] s10960, in10960_1, in10960_2;
    wire c10960;
    assign in10960_1 = {c8600};
    assign in10960_2 = {c8601};
    Full_Adder FA_10960(s10960, c10960, in10960_1, in10960_2, c8599);
    wire[0:0] s10961, in10961_1, in10961_2;
    wire c10961;
    assign in10961_1 = {c8603};
    assign in10961_2 = {c8604};
    Full_Adder FA_10961(s10961, c10961, in10961_1, in10961_2, c8602);
    wire[0:0] s10962, in10962_1, in10962_2;
    wire c10962;
    assign in10962_1 = {c8606};
    assign in10962_2 = {c8607};
    Full_Adder FA_10962(s10962, c10962, in10962_1, in10962_2, c8605);
    wire[0:0] s10963, in10963_1, in10963_2;
    wire c10963;
    assign in10963_1 = {s8609[0]};
    assign in10963_2 = {s8610[0]};
    Full_Adder FA_10963(s10963, c10963, in10963_1, in10963_2, c8608);
    wire[0:0] s10964, in10964_1, in10964_2;
    wire c10964;
    assign in10964_1 = {s8612[0]};
    assign in10964_2 = {s8613[0]};
    Full_Adder FA_10964(s10964, c10964, in10964_1, in10964_2, s8611[0]);
    wire[0:0] s10965, in10965_1, in10965_2;
    wire c10965;
    assign in10965_1 = {s8615[0]};
    assign in10965_2 = {s8616[0]};
    Full_Adder FA_10965(s10965, c10965, in10965_1, in10965_2, s8614[0]);
    wire[0:0] s10966, in10966_1, in10966_2;
    wire c10966;
    assign in10966_1 = {s8618[0]};
    assign in10966_2 = {s8619[0]};
    Full_Adder FA_10966(s10966, c10966, in10966_1, in10966_2, s8617[0]);
    wire[0:0] s10967, in10967_1, in10967_2;
    wire c10967;
    assign in10967_1 = {c8610};
    assign in10967_2 = {c8611};
    Full_Adder FA_10967(s10967, c10967, in10967_1, in10967_2, c8609);
    wire[0:0] s10968, in10968_1, in10968_2;
    wire c10968;
    assign in10968_1 = {c8613};
    assign in10968_2 = {c8614};
    Full_Adder FA_10968(s10968, c10968, in10968_1, in10968_2, c8612);
    wire[0:0] s10969, in10969_1, in10969_2;
    wire c10969;
    assign in10969_1 = {c8616};
    assign in10969_2 = {c8617};
    Full_Adder FA_10969(s10969, c10969, in10969_1, in10969_2, c8615);
    wire[0:0] s10970, in10970_1, in10970_2;
    wire c10970;
    assign in10970_1 = {c8619};
    assign in10970_2 = {c8620};
    Full_Adder FA_10970(s10970, c10970, in10970_1, in10970_2, c8618);
    wire[0:0] s10971, in10971_1, in10971_2;
    wire c10971;
    assign in10971_1 = {s8622[0]};
    assign in10971_2 = {s8623[0]};
    Full_Adder FA_10971(s10971, c10971, in10971_1, in10971_2, c8621);
    wire[0:0] s10972, in10972_1, in10972_2;
    wire c10972;
    assign in10972_1 = {s8625[0]};
    assign in10972_2 = {s8626[0]};
    Full_Adder FA_10972(s10972, c10972, in10972_1, in10972_2, s8624[0]);
    wire[0:0] s10973, in10973_1, in10973_2;
    wire c10973;
    assign in10973_1 = {s8628[0]};
    assign in10973_2 = {s8629[0]};
    Full_Adder FA_10973(s10973, c10973, in10973_1, in10973_2, s8627[0]);
    wire[0:0] s10974, in10974_1, in10974_2;
    wire c10974;
    assign in10974_1 = {s8631[0]};
    assign in10974_2 = {s8632[0]};
    Full_Adder FA_10974(s10974, c10974, in10974_1, in10974_2, s8630[0]);
    wire[0:0] s10975, in10975_1, in10975_2;
    wire c10975;
    assign in10975_1 = {c8623};
    assign in10975_2 = {c8624};
    Full_Adder FA_10975(s10975, c10975, in10975_1, in10975_2, c8622);
    wire[0:0] s10976, in10976_1, in10976_2;
    wire c10976;
    assign in10976_1 = {c8626};
    assign in10976_2 = {c8627};
    Full_Adder FA_10976(s10976, c10976, in10976_1, in10976_2, c8625);
    wire[0:0] s10977, in10977_1, in10977_2;
    wire c10977;
    assign in10977_1 = {c8629};
    assign in10977_2 = {c8630};
    Full_Adder FA_10977(s10977, c10977, in10977_1, in10977_2, c8628);
    wire[0:0] s10978, in10978_1, in10978_2;
    wire c10978;
    assign in10978_1 = {c8632};
    assign in10978_2 = {c8633};
    Full_Adder FA_10978(s10978, c10978, in10978_1, in10978_2, c8631);
    wire[0:0] s10979, in10979_1, in10979_2;
    wire c10979;
    assign in10979_1 = {s8635[0]};
    assign in10979_2 = {s8636[0]};
    Full_Adder FA_10979(s10979, c10979, in10979_1, in10979_2, c8634);
    wire[0:0] s10980, in10980_1, in10980_2;
    wire c10980;
    assign in10980_1 = {s8638[0]};
    assign in10980_2 = {s8639[0]};
    Full_Adder FA_10980(s10980, c10980, in10980_1, in10980_2, s8637[0]);
    wire[0:0] s10981, in10981_1, in10981_2;
    wire c10981;
    assign in10981_1 = {s8641[0]};
    assign in10981_2 = {s8642[0]};
    Full_Adder FA_10981(s10981, c10981, in10981_1, in10981_2, s8640[0]);
    wire[0:0] s10982, in10982_1, in10982_2;
    wire c10982;
    assign in10982_1 = {s8644[0]};
    assign in10982_2 = {s8645[0]};
    Full_Adder FA_10982(s10982, c10982, in10982_1, in10982_2, s8643[0]);
    wire[0:0] s10983, in10983_1, in10983_2;
    wire c10983;
    assign in10983_1 = {c8636};
    assign in10983_2 = {c8637};
    Full_Adder FA_10983(s10983, c10983, in10983_1, in10983_2, c8635);
    wire[0:0] s10984, in10984_1, in10984_2;
    wire c10984;
    assign in10984_1 = {c8639};
    assign in10984_2 = {c8640};
    Full_Adder FA_10984(s10984, c10984, in10984_1, in10984_2, c8638);
    wire[0:0] s10985, in10985_1, in10985_2;
    wire c10985;
    assign in10985_1 = {c8642};
    assign in10985_2 = {c8643};
    Full_Adder FA_10985(s10985, c10985, in10985_1, in10985_2, c8641);
    wire[0:0] s10986, in10986_1, in10986_2;
    wire c10986;
    assign in10986_1 = {c8645};
    assign in10986_2 = {c8646};
    Full_Adder FA_10986(s10986, c10986, in10986_1, in10986_2, c8644);
    wire[0:0] s10987, in10987_1, in10987_2;
    wire c10987;
    assign in10987_1 = {s8648[0]};
    assign in10987_2 = {s8649[0]};
    Full_Adder FA_10987(s10987, c10987, in10987_1, in10987_2, c8647);
    wire[0:0] s10988, in10988_1, in10988_2;
    wire c10988;
    assign in10988_1 = {s8651[0]};
    assign in10988_2 = {s8652[0]};
    Full_Adder FA_10988(s10988, c10988, in10988_1, in10988_2, s8650[0]);
    wire[0:0] s10989, in10989_1, in10989_2;
    wire c10989;
    assign in10989_1 = {s8654[0]};
    assign in10989_2 = {s8655[0]};
    Full_Adder FA_10989(s10989, c10989, in10989_1, in10989_2, s8653[0]);
    wire[0:0] s10990, in10990_1, in10990_2;
    wire c10990;
    assign in10990_1 = {s8657[0]};
    assign in10990_2 = {s8658[0]};
    Full_Adder FA_10990(s10990, c10990, in10990_1, in10990_2, s8656[0]);
    wire[0:0] s10991, in10991_1, in10991_2;
    wire c10991;
    assign in10991_1 = {c8649};
    assign in10991_2 = {c8650};
    Full_Adder FA_10991(s10991, c10991, in10991_1, in10991_2, c8648);
    wire[0:0] s10992, in10992_1, in10992_2;
    wire c10992;
    assign in10992_1 = {c8652};
    assign in10992_2 = {c8653};
    Full_Adder FA_10992(s10992, c10992, in10992_1, in10992_2, c8651);
    wire[0:0] s10993, in10993_1, in10993_2;
    wire c10993;
    assign in10993_1 = {c8655};
    assign in10993_2 = {c8656};
    Full_Adder FA_10993(s10993, c10993, in10993_1, in10993_2, c8654);
    wire[0:0] s10994, in10994_1, in10994_2;
    wire c10994;
    assign in10994_1 = {c8658};
    assign in10994_2 = {c8659};
    Full_Adder FA_10994(s10994, c10994, in10994_1, in10994_2, c8657);
    wire[0:0] s10995, in10995_1, in10995_2;
    wire c10995;
    assign in10995_1 = {s8661[0]};
    assign in10995_2 = {s8662[0]};
    Full_Adder FA_10995(s10995, c10995, in10995_1, in10995_2, c8660);
    wire[0:0] s10996, in10996_1, in10996_2;
    wire c10996;
    assign in10996_1 = {s8664[0]};
    assign in10996_2 = {s8665[0]};
    Full_Adder FA_10996(s10996, c10996, in10996_1, in10996_2, s8663[0]);
    wire[0:0] s10997, in10997_1, in10997_2;
    wire c10997;
    assign in10997_1 = {s8667[0]};
    assign in10997_2 = {s8668[0]};
    Full_Adder FA_10997(s10997, c10997, in10997_1, in10997_2, s8666[0]);
    wire[0:0] s10998, in10998_1, in10998_2;
    wire c10998;
    assign in10998_1 = {s8670[0]};
    assign in10998_2 = {s8671[0]};
    Full_Adder FA_10998(s10998, c10998, in10998_1, in10998_2, s8669[0]);
    wire[0:0] s10999, in10999_1, in10999_2;
    wire c10999;
    assign in10999_1 = {c8662};
    assign in10999_2 = {c8663};
    Full_Adder FA_10999(s10999, c10999, in10999_1, in10999_2, c8661);
    wire[0:0] s11000, in11000_1, in11000_2;
    wire c11000;
    assign in11000_1 = {c8665};
    assign in11000_2 = {c8666};
    Full_Adder FA_11000(s11000, c11000, in11000_1, in11000_2, c8664);
    wire[0:0] s11001, in11001_1, in11001_2;
    wire c11001;
    assign in11001_1 = {c8668};
    assign in11001_2 = {c8669};
    Full_Adder FA_11001(s11001, c11001, in11001_1, in11001_2, c8667);
    wire[0:0] s11002, in11002_1, in11002_2;
    wire c11002;
    assign in11002_1 = {c8671};
    assign in11002_2 = {c8672};
    Full_Adder FA_11002(s11002, c11002, in11002_1, in11002_2, c8670);
    wire[0:0] s11003, in11003_1, in11003_2;
    wire c11003;
    assign in11003_1 = {s8674[0]};
    assign in11003_2 = {s8675[0]};
    Full_Adder FA_11003(s11003, c11003, in11003_1, in11003_2, c8673);
    wire[0:0] s11004, in11004_1, in11004_2;
    wire c11004;
    assign in11004_1 = {s8677[0]};
    assign in11004_2 = {s8678[0]};
    Full_Adder FA_11004(s11004, c11004, in11004_1, in11004_2, s8676[0]);
    wire[0:0] s11005, in11005_1, in11005_2;
    wire c11005;
    assign in11005_1 = {s8680[0]};
    assign in11005_2 = {s8681[0]};
    Full_Adder FA_11005(s11005, c11005, in11005_1, in11005_2, s8679[0]);
    wire[0:0] s11006, in11006_1, in11006_2;
    wire c11006;
    assign in11006_1 = {s8683[0]};
    assign in11006_2 = {s8684[0]};
    Full_Adder FA_11006(s11006, c11006, in11006_1, in11006_2, s8682[0]);
    wire[0:0] s11007, in11007_1, in11007_2;
    wire c11007;
    assign in11007_1 = {c8675};
    assign in11007_2 = {c8676};
    Full_Adder FA_11007(s11007, c11007, in11007_1, in11007_2, c8674);
    wire[0:0] s11008, in11008_1, in11008_2;
    wire c11008;
    assign in11008_1 = {c8678};
    assign in11008_2 = {c8679};
    Full_Adder FA_11008(s11008, c11008, in11008_1, in11008_2, c8677);
    wire[0:0] s11009, in11009_1, in11009_2;
    wire c11009;
    assign in11009_1 = {c8681};
    assign in11009_2 = {c8682};
    Full_Adder FA_11009(s11009, c11009, in11009_1, in11009_2, c8680);
    wire[0:0] s11010, in11010_1, in11010_2;
    wire c11010;
    assign in11010_1 = {c8684};
    assign in11010_2 = {c8685};
    Full_Adder FA_11010(s11010, c11010, in11010_1, in11010_2, c8683);
    wire[0:0] s11011, in11011_1, in11011_2;
    wire c11011;
    assign in11011_1 = {s8687[0]};
    assign in11011_2 = {s8688[0]};
    Full_Adder FA_11011(s11011, c11011, in11011_1, in11011_2, c8686);
    wire[0:0] s11012, in11012_1, in11012_2;
    wire c11012;
    assign in11012_1 = {s8690[0]};
    assign in11012_2 = {s8691[0]};
    Full_Adder FA_11012(s11012, c11012, in11012_1, in11012_2, s8689[0]);
    wire[0:0] s11013, in11013_1, in11013_2;
    wire c11013;
    assign in11013_1 = {s8693[0]};
    assign in11013_2 = {s8694[0]};
    Full_Adder FA_11013(s11013, c11013, in11013_1, in11013_2, s8692[0]);
    wire[0:0] s11014, in11014_1, in11014_2;
    wire c11014;
    assign in11014_1 = {s8696[0]};
    assign in11014_2 = {s8697[0]};
    Full_Adder FA_11014(s11014, c11014, in11014_1, in11014_2, s8695[0]);
    wire[0:0] s11015, in11015_1, in11015_2;
    wire c11015;
    assign in11015_1 = {c8688};
    assign in11015_2 = {c8689};
    Full_Adder FA_11015(s11015, c11015, in11015_1, in11015_2, c8687);
    wire[0:0] s11016, in11016_1, in11016_2;
    wire c11016;
    assign in11016_1 = {c8691};
    assign in11016_2 = {c8692};
    Full_Adder FA_11016(s11016, c11016, in11016_1, in11016_2, c8690);
    wire[0:0] s11017, in11017_1, in11017_2;
    wire c11017;
    assign in11017_1 = {c8694};
    assign in11017_2 = {c8695};
    Full_Adder FA_11017(s11017, c11017, in11017_1, in11017_2, c8693);
    wire[0:0] s11018, in11018_1, in11018_2;
    wire c11018;
    assign in11018_1 = {c8697};
    assign in11018_2 = {c8698};
    Full_Adder FA_11018(s11018, c11018, in11018_1, in11018_2, c8696);
    wire[0:0] s11019, in11019_1, in11019_2;
    wire c11019;
    assign in11019_1 = {s8700[0]};
    assign in11019_2 = {s8701[0]};
    Full_Adder FA_11019(s11019, c11019, in11019_1, in11019_2, c8699);
    wire[0:0] s11020, in11020_1, in11020_2;
    wire c11020;
    assign in11020_1 = {s8703[0]};
    assign in11020_2 = {s8704[0]};
    Full_Adder FA_11020(s11020, c11020, in11020_1, in11020_2, s8702[0]);
    wire[0:0] s11021, in11021_1, in11021_2;
    wire c11021;
    assign in11021_1 = {s8706[0]};
    assign in11021_2 = {s8707[0]};
    Full_Adder FA_11021(s11021, c11021, in11021_1, in11021_2, s8705[0]);
    wire[0:0] s11022, in11022_1, in11022_2;
    wire c11022;
    assign in11022_1 = {s8709[0]};
    assign in11022_2 = {s8710[0]};
    Full_Adder FA_11022(s11022, c11022, in11022_1, in11022_2, s8708[0]);
    wire[0:0] s11023, in11023_1, in11023_2;
    wire c11023;
    assign in11023_1 = {c8701};
    assign in11023_2 = {c8702};
    Full_Adder FA_11023(s11023, c11023, in11023_1, in11023_2, c8700);
    wire[0:0] s11024, in11024_1, in11024_2;
    wire c11024;
    assign in11024_1 = {c8704};
    assign in11024_2 = {c8705};
    Full_Adder FA_11024(s11024, c11024, in11024_1, in11024_2, c8703);
    wire[0:0] s11025, in11025_1, in11025_2;
    wire c11025;
    assign in11025_1 = {c8707};
    assign in11025_2 = {c8708};
    Full_Adder FA_11025(s11025, c11025, in11025_1, in11025_2, c8706);
    wire[0:0] s11026, in11026_1, in11026_2;
    wire c11026;
    assign in11026_1 = {c8710};
    assign in11026_2 = {c8711};
    Full_Adder FA_11026(s11026, c11026, in11026_1, in11026_2, c8709);
    wire[0:0] s11027, in11027_1, in11027_2;
    wire c11027;
    assign in11027_1 = {s8713[0]};
    assign in11027_2 = {s8714[0]};
    Full_Adder FA_11027(s11027, c11027, in11027_1, in11027_2, c8712);
    wire[0:0] s11028, in11028_1, in11028_2;
    wire c11028;
    assign in11028_1 = {s8716[0]};
    assign in11028_2 = {s8717[0]};
    Full_Adder FA_11028(s11028, c11028, in11028_1, in11028_2, s8715[0]);
    wire[0:0] s11029, in11029_1, in11029_2;
    wire c11029;
    assign in11029_1 = {s8719[0]};
    assign in11029_2 = {s8720[0]};
    Full_Adder FA_11029(s11029, c11029, in11029_1, in11029_2, s8718[0]);
    wire[0:0] s11030, in11030_1, in11030_2;
    wire c11030;
    assign in11030_1 = {s8722[0]};
    assign in11030_2 = {s8723[0]};
    Full_Adder FA_11030(s11030, c11030, in11030_1, in11030_2, s8721[0]);
    wire[0:0] s11031, in11031_1, in11031_2;
    wire c11031;
    assign in11031_1 = {c8714};
    assign in11031_2 = {c8715};
    Full_Adder FA_11031(s11031, c11031, in11031_1, in11031_2, c8713);
    wire[0:0] s11032, in11032_1, in11032_2;
    wire c11032;
    assign in11032_1 = {c8717};
    assign in11032_2 = {c8718};
    Full_Adder FA_11032(s11032, c11032, in11032_1, in11032_2, c8716);
    wire[0:0] s11033, in11033_1, in11033_2;
    wire c11033;
    assign in11033_1 = {c8720};
    assign in11033_2 = {c8721};
    Full_Adder FA_11033(s11033, c11033, in11033_1, in11033_2, c8719);
    wire[0:0] s11034, in11034_1, in11034_2;
    wire c11034;
    assign in11034_1 = {c8723};
    assign in11034_2 = {c8724};
    Full_Adder FA_11034(s11034, c11034, in11034_1, in11034_2, c8722);
    wire[0:0] s11035, in11035_1, in11035_2;
    wire c11035;
    assign in11035_1 = {s8726[0]};
    assign in11035_2 = {s8727[0]};
    Full_Adder FA_11035(s11035, c11035, in11035_1, in11035_2, c8725);
    wire[0:0] s11036, in11036_1, in11036_2;
    wire c11036;
    assign in11036_1 = {s8729[0]};
    assign in11036_2 = {s8730[0]};
    Full_Adder FA_11036(s11036, c11036, in11036_1, in11036_2, s8728[0]);
    wire[0:0] s11037, in11037_1, in11037_2;
    wire c11037;
    assign in11037_1 = {s8732[0]};
    assign in11037_2 = {s8733[0]};
    Full_Adder FA_11037(s11037, c11037, in11037_1, in11037_2, s8731[0]);
    wire[0:0] s11038, in11038_1, in11038_2;
    wire c11038;
    assign in11038_1 = {s8735[0]};
    assign in11038_2 = {s8736[0]};
    Full_Adder FA_11038(s11038, c11038, in11038_1, in11038_2, s8734[0]);
    wire[0:0] s11039, in11039_1, in11039_2;
    wire c11039;
    assign in11039_1 = {c8727};
    assign in11039_2 = {c8728};
    Full_Adder FA_11039(s11039, c11039, in11039_1, in11039_2, c8726);
    wire[0:0] s11040, in11040_1, in11040_2;
    wire c11040;
    assign in11040_1 = {c8730};
    assign in11040_2 = {c8731};
    Full_Adder FA_11040(s11040, c11040, in11040_1, in11040_2, c8729);
    wire[0:0] s11041, in11041_1, in11041_2;
    wire c11041;
    assign in11041_1 = {c8733};
    assign in11041_2 = {c8734};
    Full_Adder FA_11041(s11041, c11041, in11041_1, in11041_2, c8732);
    wire[0:0] s11042, in11042_1, in11042_2;
    wire c11042;
    assign in11042_1 = {c8736};
    assign in11042_2 = {c8737};
    Full_Adder FA_11042(s11042, c11042, in11042_1, in11042_2, c8735);
    wire[0:0] s11043, in11043_1, in11043_2;
    wire c11043;
    assign in11043_1 = {s8739[0]};
    assign in11043_2 = {s8740[0]};
    Full_Adder FA_11043(s11043, c11043, in11043_1, in11043_2, c8738);
    wire[0:0] s11044, in11044_1, in11044_2;
    wire c11044;
    assign in11044_1 = {s8742[0]};
    assign in11044_2 = {s8743[0]};
    Full_Adder FA_11044(s11044, c11044, in11044_1, in11044_2, s8741[0]);
    wire[0:0] s11045, in11045_1, in11045_2;
    wire c11045;
    assign in11045_1 = {s8745[0]};
    assign in11045_2 = {s8746[0]};
    Full_Adder FA_11045(s11045, c11045, in11045_1, in11045_2, s8744[0]);
    wire[0:0] s11046, in11046_1, in11046_2;
    wire c11046;
    assign in11046_1 = {s8748[0]};
    assign in11046_2 = {s8749[0]};
    Full_Adder FA_11046(s11046, c11046, in11046_1, in11046_2, s8747[0]);
    wire[0:0] s11047, in11047_1, in11047_2;
    wire c11047;
    assign in11047_1 = {c8740};
    assign in11047_2 = {c8741};
    Full_Adder FA_11047(s11047, c11047, in11047_1, in11047_2, c8739);
    wire[0:0] s11048, in11048_1, in11048_2;
    wire c11048;
    assign in11048_1 = {c8743};
    assign in11048_2 = {c8744};
    Full_Adder FA_11048(s11048, c11048, in11048_1, in11048_2, c8742);
    wire[0:0] s11049, in11049_1, in11049_2;
    wire c11049;
    assign in11049_1 = {c8746};
    assign in11049_2 = {c8747};
    Full_Adder FA_11049(s11049, c11049, in11049_1, in11049_2, c8745);
    wire[0:0] s11050, in11050_1, in11050_2;
    wire c11050;
    assign in11050_1 = {c8749};
    assign in11050_2 = {c8750};
    Full_Adder FA_11050(s11050, c11050, in11050_1, in11050_2, c8748);
    wire[0:0] s11051, in11051_1, in11051_2;
    wire c11051;
    assign in11051_1 = {s8752[0]};
    assign in11051_2 = {s8753[0]};
    Full_Adder FA_11051(s11051, c11051, in11051_1, in11051_2, c8751);
    wire[0:0] s11052, in11052_1, in11052_2;
    wire c11052;
    assign in11052_1 = {s8755[0]};
    assign in11052_2 = {s8756[0]};
    Full_Adder FA_11052(s11052, c11052, in11052_1, in11052_2, s8754[0]);
    wire[0:0] s11053, in11053_1, in11053_2;
    wire c11053;
    assign in11053_1 = {s8758[0]};
    assign in11053_2 = {s8759[0]};
    Full_Adder FA_11053(s11053, c11053, in11053_1, in11053_2, s8757[0]);
    wire[0:0] s11054, in11054_1, in11054_2;
    wire c11054;
    assign in11054_1 = {s8761[0]};
    assign in11054_2 = {s8762[0]};
    Full_Adder FA_11054(s11054, c11054, in11054_1, in11054_2, s8760[0]);
    wire[0:0] s11055, in11055_1, in11055_2;
    wire c11055;
    assign in11055_1 = {c8753};
    assign in11055_2 = {c8754};
    Full_Adder FA_11055(s11055, c11055, in11055_1, in11055_2, c8752);
    wire[0:0] s11056, in11056_1, in11056_2;
    wire c11056;
    assign in11056_1 = {c8756};
    assign in11056_2 = {c8757};
    Full_Adder FA_11056(s11056, c11056, in11056_1, in11056_2, c8755);
    wire[0:0] s11057, in11057_1, in11057_2;
    wire c11057;
    assign in11057_1 = {c8759};
    assign in11057_2 = {c8760};
    Full_Adder FA_11057(s11057, c11057, in11057_1, in11057_2, c8758);
    wire[0:0] s11058, in11058_1, in11058_2;
    wire c11058;
    assign in11058_1 = {c8762};
    assign in11058_2 = {c8763};
    Full_Adder FA_11058(s11058, c11058, in11058_1, in11058_2, c8761);
    wire[0:0] s11059, in11059_1, in11059_2;
    wire c11059;
    assign in11059_1 = {s8765[0]};
    assign in11059_2 = {s8766[0]};
    Full_Adder FA_11059(s11059, c11059, in11059_1, in11059_2, c8764);
    wire[0:0] s11060, in11060_1, in11060_2;
    wire c11060;
    assign in11060_1 = {s8768[0]};
    assign in11060_2 = {s8769[0]};
    Full_Adder FA_11060(s11060, c11060, in11060_1, in11060_2, s8767[0]);
    wire[0:0] s11061, in11061_1, in11061_2;
    wire c11061;
    assign in11061_1 = {s8771[0]};
    assign in11061_2 = {s8772[0]};
    Full_Adder FA_11061(s11061, c11061, in11061_1, in11061_2, s8770[0]);
    wire[0:0] s11062, in11062_1, in11062_2;
    wire c11062;
    assign in11062_1 = {s8774[0]};
    assign in11062_2 = {s8775[0]};
    Full_Adder FA_11062(s11062, c11062, in11062_1, in11062_2, s8773[0]);
    wire[0:0] s11063, in11063_1, in11063_2;
    wire c11063;
    assign in11063_1 = {c8766};
    assign in11063_2 = {c8767};
    Full_Adder FA_11063(s11063, c11063, in11063_1, in11063_2, c8765);
    wire[0:0] s11064, in11064_1, in11064_2;
    wire c11064;
    assign in11064_1 = {c8769};
    assign in11064_2 = {c8770};
    Full_Adder FA_11064(s11064, c11064, in11064_1, in11064_2, c8768);
    wire[0:0] s11065, in11065_1, in11065_2;
    wire c11065;
    assign in11065_1 = {c8772};
    assign in11065_2 = {c8773};
    Full_Adder FA_11065(s11065, c11065, in11065_1, in11065_2, c8771);
    wire[0:0] s11066, in11066_1, in11066_2;
    wire c11066;
    assign in11066_1 = {c8775};
    assign in11066_2 = {c8776};
    Full_Adder FA_11066(s11066, c11066, in11066_1, in11066_2, c8774);
    wire[0:0] s11067, in11067_1, in11067_2;
    wire c11067;
    assign in11067_1 = {s8778[0]};
    assign in11067_2 = {s8779[0]};
    Full_Adder FA_11067(s11067, c11067, in11067_1, in11067_2, c8777);
    wire[0:0] s11068, in11068_1, in11068_2;
    wire c11068;
    assign in11068_1 = {s8781[0]};
    assign in11068_2 = {s8782[0]};
    Full_Adder FA_11068(s11068, c11068, in11068_1, in11068_2, s8780[0]);
    wire[0:0] s11069, in11069_1, in11069_2;
    wire c11069;
    assign in11069_1 = {s8784[0]};
    assign in11069_2 = {s8785[0]};
    Full_Adder FA_11069(s11069, c11069, in11069_1, in11069_2, s8783[0]);
    wire[0:0] s11070, in11070_1, in11070_2;
    wire c11070;
    assign in11070_1 = {s8787[0]};
    assign in11070_2 = {s8788[0]};
    Full_Adder FA_11070(s11070, c11070, in11070_1, in11070_2, s8786[0]);
    wire[0:0] s11071, in11071_1, in11071_2;
    wire c11071;
    assign in11071_1 = {c8779};
    assign in11071_2 = {c8780};
    Full_Adder FA_11071(s11071, c11071, in11071_1, in11071_2, c8778);
    wire[0:0] s11072, in11072_1, in11072_2;
    wire c11072;
    assign in11072_1 = {c8782};
    assign in11072_2 = {c8783};
    Full_Adder FA_11072(s11072, c11072, in11072_1, in11072_2, c8781);
    wire[0:0] s11073, in11073_1, in11073_2;
    wire c11073;
    assign in11073_1 = {c8785};
    assign in11073_2 = {c8786};
    Full_Adder FA_11073(s11073, c11073, in11073_1, in11073_2, c8784);
    wire[0:0] s11074, in11074_1, in11074_2;
    wire c11074;
    assign in11074_1 = {c8788};
    assign in11074_2 = {c8789};
    Full_Adder FA_11074(s11074, c11074, in11074_1, in11074_2, c8787);
    wire[0:0] s11075, in11075_1, in11075_2;
    wire c11075;
    assign in11075_1 = {s8791[0]};
    assign in11075_2 = {s8792[0]};
    Full_Adder FA_11075(s11075, c11075, in11075_1, in11075_2, c8790);
    wire[0:0] s11076, in11076_1, in11076_2;
    wire c11076;
    assign in11076_1 = {s8794[0]};
    assign in11076_2 = {s8795[0]};
    Full_Adder FA_11076(s11076, c11076, in11076_1, in11076_2, s8793[0]);
    wire[0:0] s11077, in11077_1, in11077_2;
    wire c11077;
    assign in11077_1 = {s8797[0]};
    assign in11077_2 = {s8798[0]};
    Full_Adder FA_11077(s11077, c11077, in11077_1, in11077_2, s8796[0]);
    wire[0:0] s11078, in11078_1, in11078_2;
    wire c11078;
    assign in11078_1 = {s8800[0]};
    assign in11078_2 = {s8801[0]};
    Full_Adder FA_11078(s11078, c11078, in11078_1, in11078_2, s8799[0]);
    wire[0:0] s11079, in11079_1, in11079_2;
    wire c11079;
    assign in11079_1 = {c8792};
    assign in11079_2 = {c8793};
    Full_Adder FA_11079(s11079, c11079, in11079_1, in11079_2, c8791);
    wire[0:0] s11080, in11080_1, in11080_2;
    wire c11080;
    assign in11080_1 = {c8795};
    assign in11080_2 = {c8796};
    Full_Adder FA_11080(s11080, c11080, in11080_1, in11080_2, c8794);
    wire[0:0] s11081, in11081_1, in11081_2;
    wire c11081;
    assign in11081_1 = {c8798};
    assign in11081_2 = {c8799};
    Full_Adder FA_11081(s11081, c11081, in11081_1, in11081_2, c8797);
    wire[0:0] s11082, in11082_1, in11082_2;
    wire c11082;
    assign in11082_1 = {c8801};
    assign in11082_2 = {c8802};
    Full_Adder FA_11082(s11082, c11082, in11082_1, in11082_2, c8800);
    wire[0:0] s11083, in11083_1, in11083_2;
    wire c11083;
    assign in11083_1 = {s8804[0]};
    assign in11083_2 = {s8805[0]};
    Full_Adder FA_11083(s11083, c11083, in11083_1, in11083_2, c8803);
    wire[0:0] s11084, in11084_1, in11084_2;
    wire c11084;
    assign in11084_1 = {s8807[0]};
    assign in11084_2 = {s8808[0]};
    Full_Adder FA_11084(s11084, c11084, in11084_1, in11084_2, s8806[0]);
    wire[0:0] s11085, in11085_1, in11085_2;
    wire c11085;
    assign in11085_1 = {s8810[0]};
    assign in11085_2 = {s8811[0]};
    Full_Adder FA_11085(s11085, c11085, in11085_1, in11085_2, s8809[0]);
    wire[0:0] s11086, in11086_1, in11086_2;
    wire c11086;
    assign in11086_1 = {s8813[0]};
    assign in11086_2 = {s8814[0]};
    Full_Adder FA_11086(s11086, c11086, in11086_1, in11086_2, s8812[0]);
    wire[0:0] s11087, in11087_1, in11087_2;
    wire c11087;
    assign in11087_1 = {c8805};
    assign in11087_2 = {c8806};
    Full_Adder FA_11087(s11087, c11087, in11087_1, in11087_2, c8804);
    wire[0:0] s11088, in11088_1, in11088_2;
    wire c11088;
    assign in11088_1 = {c8808};
    assign in11088_2 = {c8809};
    Full_Adder FA_11088(s11088, c11088, in11088_1, in11088_2, c8807);
    wire[0:0] s11089, in11089_1, in11089_2;
    wire c11089;
    assign in11089_1 = {c8811};
    assign in11089_2 = {c8812};
    Full_Adder FA_11089(s11089, c11089, in11089_1, in11089_2, c8810);
    wire[0:0] s11090, in11090_1, in11090_2;
    wire c11090;
    assign in11090_1 = {c8814};
    assign in11090_2 = {c8815};
    Full_Adder FA_11090(s11090, c11090, in11090_1, in11090_2, c8813);
    wire[0:0] s11091, in11091_1, in11091_2;
    wire c11091;
    assign in11091_1 = {s8817[0]};
    assign in11091_2 = {s8818[0]};
    Full_Adder FA_11091(s11091, c11091, in11091_1, in11091_2, c8816);
    wire[0:0] s11092, in11092_1, in11092_2;
    wire c11092;
    assign in11092_1 = {s8820[0]};
    assign in11092_2 = {s8821[0]};
    Full_Adder FA_11092(s11092, c11092, in11092_1, in11092_2, s8819[0]);
    wire[0:0] s11093, in11093_1, in11093_2;
    wire c11093;
    assign in11093_1 = {s8823[0]};
    assign in11093_2 = {s8824[0]};
    Full_Adder FA_11093(s11093, c11093, in11093_1, in11093_2, s8822[0]);
    wire[0:0] s11094, in11094_1, in11094_2;
    wire c11094;
    assign in11094_1 = {s8826[0]};
    assign in11094_2 = {s8827[0]};
    Full_Adder FA_11094(s11094, c11094, in11094_1, in11094_2, s8825[0]);
    wire[0:0] s11095, in11095_1, in11095_2;
    wire c11095;
    assign in11095_1 = {c8818};
    assign in11095_2 = {c8819};
    Full_Adder FA_11095(s11095, c11095, in11095_1, in11095_2, c8817);
    wire[0:0] s11096, in11096_1, in11096_2;
    wire c11096;
    assign in11096_1 = {c8821};
    assign in11096_2 = {c8822};
    Full_Adder FA_11096(s11096, c11096, in11096_1, in11096_2, c8820);
    wire[0:0] s11097, in11097_1, in11097_2;
    wire c11097;
    assign in11097_1 = {c8824};
    assign in11097_2 = {c8825};
    Full_Adder FA_11097(s11097, c11097, in11097_1, in11097_2, c8823);
    wire[0:0] s11098, in11098_1, in11098_2;
    wire c11098;
    assign in11098_1 = {c8827};
    assign in11098_2 = {c8828};
    Full_Adder FA_11098(s11098, c11098, in11098_1, in11098_2, c8826);
    wire[0:0] s11099, in11099_1, in11099_2;
    wire c11099;
    assign in11099_1 = {s8830[0]};
    assign in11099_2 = {s8831[0]};
    Full_Adder FA_11099(s11099, c11099, in11099_1, in11099_2, c8829);
    wire[0:0] s11100, in11100_1, in11100_2;
    wire c11100;
    assign in11100_1 = {s8833[0]};
    assign in11100_2 = {s8834[0]};
    Full_Adder FA_11100(s11100, c11100, in11100_1, in11100_2, s8832[0]);
    wire[0:0] s11101, in11101_1, in11101_2;
    wire c11101;
    assign in11101_1 = {s8836[0]};
    assign in11101_2 = {s8837[0]};
    Full_Adder FA_11101(s11101, c11101, in11101_1, in11101_2, s8835[0]);
    wire[0:0] s11102, in11102_1, in11102_2;
    wire c11102;
    assign in11102_1 = {s8839[0]};
    assign in11102_2 = {s8840[0]};
    Full_Adder FA_11102(s11102, c11102, in11102_1, in11102_2, s8838[0]);
    wire[0:0] s11103, in11103_1, in11103_2;
    wire c11103;
    assign in11103_1 = {c8831};
    assign in11103_2 = {c8832};
    Full_Adder FA_11103(s11103, c11103, in11103_1, in11103_2, c8830);
    wire[0:0] s11104, in11104_1, in11104_2;
    wire c11104;
    assign in11104_1 = {c8834};
    assign in11104_2 = {c8835};
    Full_Adder FA_11104(s11104, c11104, in11104_1, in11104_2, c8833);
    wire[0:0] s11105, in11105_1, in11105_2;
    wire c11105;
    assign in11105_1 = {c8837};
    assign in11105_2 = {c8838};
    Full_Adder FA_11105(s11105, c11105, in11105_1, in11105_2, c8836);
    wire[0:0] s11106, in11106_1, in11106_2;
    wire c11106;
    assign in11106_1 = {c8840};
    assign in11106_2 = {c8841};
    Full_Adder FA_11106(s11106, c11106, in11106_1, in11106_2, c8839);
    wire[0:0] s11107, in11107_1, in11107_2;
    wire c11107;
    assign in11107_1 = {s8843[0]};
    assign in11107_2 = {s8844[0]};
    Full_Adder FA_11107(s11107, c11107, in11107_1, in11107_2, c8842);
    wire[0:0] s11108, in11108_1, in11108_2;
    wire c11108;
    assign in11108_1 = {s8846[0]};
    assign in11108_2 = {s8847[0]};
    Full_Adder FA_11108(s11108, c11108, in11108_1, in11108_2, s8845[0]);
    wire[0:0] s11109, in11109_1, in11109_2;
    wire c11109;
    assign in11109_1 = {s8849[0]};
    assign in11109_2 = {s8850[0]};
    Full_Adder FA_11109(s11109, c11109, in11109_1, in11109_2, s8848[0]);
    wire[0:0] s11110, in11110_1, in11110_2;
    wire c11110;
    assign in11110_1 = {s8852[0]};
    assign in11110_2 = {s8853[0]};
    Full_Adder FA_11110(s11110, c11110, in11110_1, in11110_2, s8851[0]);
    wire[0:0] s11111, in11111_1, in11111_2;
    wire c11111;
    assign in11111_1 = {c8844};
    assign in11111_2 = {c8845};
    Full_Adder FA_11111(s11111, c11111, in11111_1, in11111_2, c8843);
    wire[0:0] s11112, in11112_1, in11112_2;
    wire c11112;
    assign in11112_1 = {c8847};
    assign in11112_2 = {c8848};
    Full_Adder FA_11112(s11112, c11112, in11112_1, in11112_2, c8846);
    wire[0:0] s11113, in11113_1, in11113_2;
    wire c11113;
    assign in11113_1 = {c8850};
    assign in11113_2 = {c8851};
    Full_Adder FA_11113(s11113, c11113, in11113_1, in11113_2, c8849);
    wire[0:0] s11114, in11114_1, in11114_2;
    wire c11114;
    assign in11114_1 = {c8853};
    assign in11114_2 = {c8854};
    Full_Adder FA_11114(s11114, c11114, in11114_1, in11114_2, c8852);
    wire[0:0] s11115, in11115_1, in11115_2;
    wire c11115;
    assign in11115_1 = {s8856[0]};
    assign in11115_2 = {s8857[0]};
    Full_Adder FA_11115(s11115, c11115, in11115_1, in11115_2, c8855);
    wire[0:0] s11116, in11116_1, in11116_2;
    wire c11116;
    assign in11116_1 = {s8859[0]};
    assign in11116_2 = {s8860[0]};
    Full_Adder FA_11116(s11116, c11116, in11116_1, in11116_2, s8858[0]);
    wire[0:0] s11117, in11117_1, in11117_2;
    wire c11117;
    assign in11117_1 = {s8862[0]};
    assign in11117_2 = {s8863[0]};
    Full_Adder FA_11117(s11117, c11117, in11117_1, in11117_2, s8861[0]);
    wire[0:0] s11118, in11118_1, in11118_2;
    wire c11118;
    assign in11118_1 = {s8865[0]};
    assign in11118_2 = {s8866[0]};
    Full_Adder FA_11118(s11118, c11118, in11118_1, in11118_2, s8864[0]);
    wire[0:0] s11119, in11119_1, in11119_2;
    wire c11119;
    assign in11119_1 = {c8857};
    assign in11119_2 = {c8858};
    Full_Adder FA_11119(s11119, c11119, in11119_1, in11119_2, c8856);
    wire[0:0] s11120, in11120_1, in11120_2;
    wire c11120;
    assign in11120_1 = {c8860};
    assign in11120_2 = {c8861};
    Full_Adder FA_11120(s11120, c11120, in11120_1, in11120_2, c8859);
    wire[0:0] s11121, in11121_1, in11121_2;
    wire c11121;
    assign in11121_1 = {c8863};
    assign in11121_2 = {c8864};
    Full_Adder FA_11121(s11121, c11121, in11121_1, in11121_2, c8862);
    wire[0:0] s11122, in11122_1, in11122_2;
    wire c11122;
    assign in11122_1 = {c8866};
    assign in11122_2 = {c8867};
    Full_Adder FA_11122(s11122, c11122, in11122_1, in11122_2, c8865);
    wire[0:0] s11123, in11123_1, in11123_2;
    wire c11123;
    assign in11123_1 = {s8869[0]};
    assign in11123_2 = {s8870[0]};
    Full_Adder FA_11123(s11123, c11123, in11123_1, in11123_2, c8868);
    wire[0:0] s11124, in11124_1, in11124_2;
    wire c11124;
    assign in11124_1 = {s8872[0]};
    assign in11124_2 = {s8873[0]};
    Full_Adder FA_11124(s11124, c11124, in11124_1, in11124_2, s8871[0]);
    wire[0:0] s11125, in11125_1, in11125_2;
    wire c11125;
    assign in11125_1 = {s8875[0]};
    assign in11125_2 = {s8876[0]};
    Full_Adder FA_11125(s11125, c11125, in11125_1, in11125_2, s8874[0]);
    wire[0:0] s11126, in11126_1, in11126_2;
    wire c11126;
    assign in11126_1 = {s8878[0]};
    assign in11126_2 = {s8879[0]};
    Full_Adder FA_11126(s11126, c11126, in11126_1, in11126_2, s8877[0]);
    wire[0:0] s11127, in11127_1, in11127_2;
    wire c11127;
    assign in11127_1 = {c8870};
    assign in11127_2 = {c8871};
    Full_Adder FA_11127(s11127, c11127, in11127_1, in11127_2, c8869);
    wire[0:0] s11128, in11128_1, in11128_2;
    wire c11128;
    assign in11128_1 = {c8873};
    assign in11128_2 = {c8874};
    Full_Adder FA_11128(s11128, c11128, in11128_1, in11128_2, c8872);
    wire[0:0] s11129, in11129_1, in11129_2;
    wire c11129;
    assign in11129_1 = {c8876};
    assign in11129_2 = {c8877};
    Full_Adder FA_11129(s11129, c11129, in11129_1, in11129_2, c8875);
    wire[0:0] s11130, in11130_1, in11130_2;
    wire c11130;
    assign in11130_1 = {c8879};
    assign in11130_2 = {c8880};
    Full_Adder FA_11130(s11130, c11130, in11130_1, in11130_2, c8878);
    wire[0:0] s11131, in11131_1, in11131_2;
    wire c11131;
    assign in11131_1 = {s8882[0]};
    assign in11131_2 = {s8883[0]};
    Full_Adder FA_11131(s11131, c11131, in11131_1, in11131_2, c8881);
    wire[0:0] s11132, in11132_1, in11132_2;
    wire c11132;
    assign in11132_1 = {s8885[0]};
    assign in11132_2 = {s8886[0]};
    Full_Adder FA_11132(s11132, c11132, in11132_1, in11132_2, s8884[0]);
    wire[0:0] s11133, in11133_1, in11133_2;
    wire c11133;
    assign in11133_1 = {s8888[0]};
    assign in11133_2 = {s8889[0]};
    Full_Adder FA_11133(s11133, c11133, in11133_1, in11133_2, s8887[0]);
    wire[0:0] s11134, in11134_1, in11134_2;
    wire c11134;
    assign in11134_1 = {s8891[0]};
    assign in11134_2 = {s8892[0]};
    Full_Adder FA_11134(s11134, c11134, in11134_1, in11134_2, s8890[0]);
    wire[0:0] s11135, in11135_1, in11135_2;
    wire c11135;
    assign in11135_1 = {c8883};
    assign in11135_2 = {c8884};
    Full_Adder FA_11135(s11135, c11135, in11135_1, in11135_2, c8882);
    wire[0:0] s11136, in11136_1, in11136_2;
    wire c11136;
    assign in11136_1 = {c8886};
    assign in11136_2 = {c8887};
    Full_Adder FA_11136(s11136, c11136, in11136_1, in11136_2, c8885);
    wire[0:0] s11137, in11137_1, in11137_2;
    wire c11137;
    assign in11137_1 = {c8889};
    assign in11137_2 = {c8890};
    Full_Adder FA_11137(s11137, c11137, in11137_1, in11137_2, c8888);
    wire[0:0] s11138, in11138_1, in11138_2;
    wire c11138;
    assign in11138_1 = {c8892};
    assign in11138_2 = {c8893};
    Full_Adder FA_11138(s11138, c11138, in11138_1, in11138_2, c8891);
    wire[0:0] s11139, in11139_1, in11139_2;
    wire c11139;
    assign in11139_1 = {s8895[0]};
    assign in11139_2 = {s8896[0]};
    Full_Adder FA_11139(s11139, c11139, in11139_1, in11139_2, c8894);
    wire[0:0] s11140, in11140_1, in11140_2;
    wire c11140;
    assign in11140_1 = {s8898[0]};
    assign in11140_2 = {s8899[0]};
    Full_Adder FA_11140(s11140, c11140, in11140_1, in11140_2, s8897[0]);
    wire[0:0] s11141, in11141_1, in11141_2;
    wire c11141;
    assign in11141_1 = {s8901[0]};
    assign in11141_2 = {s8902[0]};
    Full_Adder FA_11141(s11141, c11141, in11141_1, in11141_2, s8900[0]);
    wire[0:0] s11142, in11142_1, in11142_2;
    wire c11142;
    assign in11142_1 = {s8904[0]};
    assign in11142_2 = {s8905[0]};
    Full_Adder FA_11142(s11142, c11142, in11142_1, in11142_2, s8903[0]);
    wire[0:0] s11143, in11143_1, in11143_2;
    wire c11143;
    assign in11143_1 = {c8896};
    assign in11143_2 = {c8897};
    Full_Adder FA_11143(s11143, c11143, in11143_1, in11143_2, c8895);
    wire[0:0] s11144, in11144_1, in11144_2;
    wire c11144;
    assign in11144_1 = {c8899};
    assign in11144_2 = {c8900};
    Full_Adder FA_11144(s11144, c11144, in11144_1, in11144_2, c8898);
    wire[0:0] s11145, in11145_1, in11145_2;
    wire c11145;
    assign in11145_1 = {c8902};
    assign in11145_2 = {c8903};
    Full_Adder FA_11145(s11145, c11145, in11145_1, in11145_2, c8901);
    wire[0:0] s11146, in11146_1, in11146_2;
    wire c11146;
    assign in11146_1 = {c8905};
    assign in11146_2 = {c8906};
    Full_Adder FA_11146(s11146, c11146, in11146_1, in11146_2, c8904);
    wire[0:0] s11147, in11147_1, in11147_2;
    wire c11147;
    assign in11147_1 = {s8908[0]};
    assign in11147_2 = {s8909[0]};
    Full_Adder FA_11147(s11147, c11147, in11147_1, in11147_2, c8907);
    wire[0:0] s11148, in11148_1, in11148_2;
    wire c11148;
    assign in11148_1 = {s8911[0]};
    assign in11148_2 = {s8912[0]};
    Full_Adder FA_11148(s11148, c11148, in11148_1, in11148_2, s8910[0]);
    wire[0:0] s11149, in11149_1, in11149_2;
    wire c11149;
    assign in11149_1 = {s8914[0]};
    assign in11149_2 = {s8915[0]};
    Full_Adder FA_11149(s11149, c11149, in11149_1, in11149_2, s8913[0]);
    wire[0:0] s11150, in11150_1, in11150_2;
    wire c11150;
    assign in11150_1 = {s8917[0]};
    assign in11150_2 = {s8918[0]};
    Full_Adder FA_11150(s11150, c11150, in11150_1, in11150_2, s8916[0]);
    wire[0:0] s11151, in11151_1, in11151_2;
    wire c11151;
    assign in11151_1 = {c8909};
    assign in11151_2 = {c8910};
    Full_Adder FA_11151(s11151, c11151, in11151_1, in11151_2, c8908);
    wire[0:0] s11152, in11152_1, in11152_2;
    wire c11152;
    assign in11152_1 = {c8912};
    assign in11152_2 = {c8913};
    Full_Adder FA_11152(s11152, c11152, in11152_1, in11152_2, c8911);
    wire[0:0] s11153, in11153_1, in11153_2;
    wire c11153;
    assign in11153_1 = {c8915};
    assign in11153_2 = {c8916};
    Full_Adder FA_11153(s11153, c11153, in11153_1, in11153_2, c8914);
    wire[0:0] s11154, in11154_1, in11154_2;
    wire c11154;
    assign in11154_1 = {c8918};
    assign in11154_2 = {c8919};
    Full_Adder FA_11154(s11154, c11154, in11154_1, in11154_2, c8917);
    wire[0:0] s11155, in11155_1, in11155_2;
    wire c11155;
    assign in11155_1 = {s8921[0]};
    assign in11155_2 = {s8922[0]};
    Full_Adder FA_11155(s11155, c11155, in11155_1, in11155_2, c8920);
    wire[0:0] s11156, in11156_1, in11156_2;
    wire c11156;
    assign in11156_1 = {s8924[0]};
    assign in11156_2 = {s8925[0]};
    Full_Adder FA_11156(s11156, c11156, in11156_1, in11156_2, s8923[0]);
    wire[0:0] s11157, in11157_1, in11157_2;
    wire c11157;
    assign in11157_1 = {s8927[0]};
    assign in11157_2 = {s8928[0]};
    Full_Adder FA_11157(s11157, c11157, in11157_1, in11157_2, s8926[0]);
    wire[0:0] s11158, in11158_1, in11158_2;
    wire c11158;
    assign in11158_1 = {s8930[0]};
    assign in11158_2 = {s8931[0]};
    Full_Adder FA_11158(s11158, c11158, in11158_1, in11158_2, s8929[0]);
    wire[0:0] s11159, in11159_1, in11159_2;
    wire c11159;
    assign in11159_1 = {c8922};
    assign in11159_2 = {c8923};
    Full_Adder FA_11159(s11159, c11159, in11159_1, in11159_2, c8921);
    wire[0:0] s11160, in11160_1, in11160_2;
    wire c11160;
    assign in11160_1 = {c8925};
    assign in11160_2 = {c8926};
    Full_Adder FA_11160(s11160, c11160, in11160_1, in11160_2, c8924);
    wire[0:0] s11161, in11161_1, in11161_2;
    wire c11161;
    assign in11161_1 = {c8928};
    assign in11161_2 = {c8929};
    Full_Adder FA_11161(s11161, c11161, in11161_1, in11161_2, c8927);
    wire[0:0] s11162, in11162_1, in11162_2;
    wire c11162;
    assign in11162_1 = {c8931};
    assign in11162_2 = {c8932};
    Full_Adder FA_11162(s11162, c11162, in11162_1, in11162_2, c8930);
    wire[0:0] s11163, in11163_1, in11163_2;
    wire c11163;
    assign in11163_1 = {s8934[0]};
    assign in11163_2 = {s8935[0]};
    Full_Adder FA_11163(s11163, c11163, in11163_1, in11163_2, c8933);
    wire[0:0] s11164, in11164_1, in11164_2;
    wire c11164;
    assign in11164_1 = {s8937[0]};
    assign in11164_2 = {s8938[0]};
    Full_Adder FA_11164(s11164, c11164, in11164_1, in11164_2, s8936[0]);
    wire[0:0] s11165, in11165_1, in11165_2;
    wire c11165;
    assign in11165_1 = {s8940[0]};
    assign in11165_2 = {s8941[0]};
    Full_Adder FA_11165(s11165, c11165, in11165_1, in11165_2, s8939[0]);
    wire[0:0] s11166, in11166_1, in11166_2;
    wire c11166;
    assign in11166_1 = {s8943[0]};
    assign in11166_2 = {s8944[0]};
    Full_Adder FA_11166(s11166, c11166, in11166_1, in11166_2, s8942[0]);
    wire[0:0] s11167, in11167_1, in11167_2;
    wire c11167;
    assign in11167_1 = {c8935};
    assign in11167_2 = {c8936};
    Full_Adder FA_11167(s11167, c11167, in11167_1, in11167_2, c8934);
    wire[0:0] s11168, in11168_1, in11168_2;
    wire c11168;
    assign in11168_1 = {c8938};
    assign in11168_2 = {c8939};
    Full_Adder FA_11168(s11168, c11168, in11168_1, in11168_2, c8937);
    wire[0:0] s11169, in11169_1, in11169_2;
    wire c11169;
    assign in11169_1 = {c8941};
    assign in11169_2 = {c8942};
    Full_Adder FA_11169(s11169, c11169, in11169_1, in11169_2, c8940);
    wire[0:0] s11170, in11170_1, in11170_2;
    wire c11170;
    assign in11170_1 = {c8944};
    assign in11170_2 = {c8945};
    Full_Adder FA_11170(s11170, c11170, in11170_1, in11170_2, c8943);
    wire[0:0] s11171, in11171_1, in11171_2;
    wire c11171;
    assign in11171_1 = {s8947[0]};
    assign in11171_2 = {s8948[0]};
    Full_Adder FA_11171(s11171, c11171, in11171_1, in11171_2, c8946);
    wire[0:0] s11172, in11172_1, in11172_2;
    wire c11172;
    assign in11172_1 = {s8950[0]};
    assign in11172_2 = {s8951[0]};
    Full_Adder FA_11172(s11172, c11172, in11172_1, in11172_2, s8949[0]);
    wire[0:0] s11173, in11173_1, in11173_2;
    wire c11173;
    assign in11173_1 = {s8953[0]};
    assign in11173_2 = {s8954[0]};
    Full_Adder FA_11173(s11173, c11173, in11173_1, in11173_2, s8952[0]);
    wire[0:0] s11174, in11174_1, in11174_2;
    wire c11174;
    assign in11174_1 = {s8956[0]};
    assign in11174_2 = {s8957[0]};
    Full_Adder FA_11174(s11174, c11174, in11174_1, in11174_2, s8955[0]);
    wire[0:0] s11175, in11175_1, in11175_2;
    wire c11175;
    assign in11175_1 = {c8948};
    assign in11175_2 = {c8949};
    Full_Adder FA_11175(s11175, c11175, in11175_1, in11175_2, c8947);
    wire[0:0] s11176, in11176_1, in11176_2;
    wire c11176;
    assign in11176_1 = {c8951};
    assign in11176_2 = {c8952};
    Full_Adder FA_11176(s11176, c11176, in11176_1, in11176_2, c8950);
    wire[0:0] s11177, in11177_1, in11177_2;
    wire c11177;
    assign in11177_1 = {c8954};
    assign in11177_2 = {c8955};
    Full_Adder FA_11177(s11177, c11177, in11177_1, in11177_2, c8953);
    wire[0:0] s11178, in11178_1, in11178_2;
    wire c11178;
    assign in11178_1 = {c8957};
    assign in11178_2 = {c8958};
    Full_Adder FA_11178(s11178, c11178, in11178_1, in11178_2, c8956);
    wire[0:0] s11179, in11179_1, in11179_2;
    wire c11179;
    assign in11179_1 = {s8960[0]};
    assign in11179_2 = {s8961[0]};
    Full_Adder FA_11179(s11179, c11179, in11179_1, in11179_2, c8959);
    wire[0:0] s11180, in11180_1, in11180_2;
    wire c11180;
    assign in11180_1 = {s8963[0]};
    assign in11180_2 = {s8964[0]};
    Full_Adder FA_11180(s11180, c11180, in11180_1, in11180_2, s8962[0]);
    wire[0:0] s11181, in11181_1, in11181_2;
    wire c11181;
    assign in11181_1 = {s8966[0]};
    assign in11181_2 = {s8967[0]};
    Full_Adder FA_11181(s11181, c11181, in11181_1, in11181_2, s8965[0]);
    wire[0:0] s11182, in11182_1, in11182_2;
    wire c11182;
    assign in11182_1 = {s8969[0]};
    assign in11182_2 = {s8970[0]};
    Full_Adder FA_11182(s11182, c11182, in11182_1, in11182_2, s8968[0]);
    wire[0:0] s11183, in11183_1, in11183_2;
    wire c11183;
    assign in11183_1 = {c8961};
    assign in11183_2 = {c8962};
    Full_Adder FA_11183(s11183, c11183, in11183_1, in11183_2, c8960);
    wire[0:0] s11184, in11184_1, in11184_2;
    wire c11184;
    assign in11184_1 = {c8964};
    assign in11184_2 = {c8965};
    Full_Adder FA_11184(s11184, c11184, in11184_1, in11184_2, c8963);
    wire[0:0] s11185, in11185_1, in11185_2;
    wire c11185;
    assign in11185_1 = {c8967};
    assign in11185_2 = {c8968};
    Full_Adder FA_11185(s11185, c11185, in11185_1, in11185_2, c8966);
    wire[0:0] s11186, in11186_1, in11186_2;
    wire c11186;
    assign in11186_1 = {c8970};
    assign in11186_2 = {c8971};
    Full_Adder FA_11186(s11186, c11186, in11186_1, in11186_2, c8969);
    wire[0:0] s11187, in11187_1, in11187_2;
    wire c11187;
    assign in11187_1 = {s8973[0]};
    assign in11187_2 = {s8974[0]};
    Full_Adder FA_11187(s11187, c11187, in11187_1, in11187_2, c8972);
    wire[0:0] s11188, in11188_1, in11188_2;
    wire c11188;
    assign in11188_1 = {s8976[0]};
    assign in11188_2 = {s8977[0]};
    Full_Adder FA_11188(s11188, c11188, in11188_1, in11188_2, s8975[0]);
    wire[0:0] s11189, in11189_1, in11189_2;
    wire c11189;
    assign in11189_1 = {s8979[0]};
    assign in11189_2 = {s8980[0]};
    Full_Adder FA_11189(s11189, c11189, in11189_1, in11189_2, s8978[0]);
    wire[0:0] s11190, in11190_1, in11190_2;
    wire c11190;
    assign in11190_1 = {s8982[0]};
    assign in11190_2 = {s8983[0]};
    Full_Adder FA_11190(s11190, c11190, in11190_1, in11190_2, s8981[0]);
    wire[0:0] s11191, in11191_1, in11191_2;
    wire c11191;
    assign in11191_1 = {c8974};
    assign in11191_2 = {c8975};
    Full_Adder FA_11191(s11191, c11191, in11191_1, in11191_2, c8973);
    wire[0:0] s11192, in11192_1, in11192_2;
    wire c11192;
    assign in11192_1 = {c8977};
    assign in11192_2 = {c8978};
    Full_Adder FA_11192(s11192, c11192, in11192_1, in11192_2, c8976);
    wire[0:0] s11193, in11193_1, in11193_2;
    wire c11193;
    assign in11193_1 = {c8980};
    assign in11193_2 = {c8981};
    Full_Adder FA_11193(s11193, c11193, in11193_1, in11193_2, c8979);
    wire[0:0] s11194, in11194_1, in11194_2;
    wire c11194;
    assign in11194_1 = {c8983};
    assign in11194_2 = {c8984};
    Full_Adder FA_11194(s11194, c11194, in11194_1, in11194_2, c8982);
    wire[0:0] s11195, in11195_1, in11195_2;
    wire c11195;
    assign in11195_1 = {s8986[0]};
    assign in11195_2 = {s8987[0]};
    Full_Adder FA_11195(s11195, c11195, in11195_1, in11195_2, c8985);
    wire[0:0] s11196, in11196_1, in11196_2;
    wire c11196;
    assign in11196_1 = {s8989[0]};
    assign in11196_2 = {s8990[0]};
    Full_Adder FA_11196(s11196, c11196, in11196_1, in11196_2, s8988[0]);
    wire[0:0] s11197, in11197_1, in11197_2;
    wire c11197;
    assign in11197_1 = {s8992[0]};
    assign in11197_2 = {s8993[0]};
    Full_Adder FA_11197(s11197, c11197, in11197_1, in11197_2, s8991[0]);
    wire[0:0] s11198, in11198_1, in11198_2;
    wire c11198;
    assign in11198_1 = {s8995[0]};
    assign in11198_2 = {s8996[0]};
    Full_Adder FA_11198(s11198, c11198, in11198_1, in11198_2, s8994[0]);
    wire[0:0] s11199, in11199_1, in11199_2;
    wire c11199;
    assign in11199_1 = {c8987};
    assign in11199_2 = {c8988};
    Full_Adder FA_11199(s11199, c11199, in11199_1, in11199_2, c8986);
    wire[0:0] s11200, in11200_1, in11200_2;
    wire c11200;
    assign in11200_1 = {c8990};
    assign in11200_2 = {c8991};
    Full_Adder FA_11200(s11200, c11200, in11200_1, in11200_2, c8989);
    wire[0:0] s11201, in11201_1, in11201_2;
    wire c11201;
    assign in11201_1 = {c8993};
    assign in11201_2 = {c8994};
    Full_Adder FA_11201(s11201, c11201, in11201_1, in11201_2, c8992);
    wire[0:0] s11202, in11202_1, in11202_2;
    wire c11202;
    assign in11202_1 = {c8996};
    assign in11202_2 = {c8997};
    Full_Adder FA_11202(s11202, c11202, in11202_1, in11202_2, c8995);
    wire[0:0] s11203, in11203_1, in11203_2;
    wire c11203;
    assign in11203_1 = {s8999[0]};
    assign in11203_2 = {s9000[0]};
    Full_Adder FA_11203(s11203, c11203, in11203_1, in11203_2, c8998);
    wire[0:0] s11204, in11204_1, in11204_2;
    wire c11204;
    assign in11204_1 = {s9002[0]};
    assign in11204_2 = {s9003[0]};
    Full_Adder FA_11204(s11204, c11204, in11204_1, in11204_2, s9001[0]);
    wire[0:0] s11205, in11205_1, in11205_2;
    wire c11205;
    assign in11205_1 = {s9005[0]};
    assign in11205_2 = {s9006[0]};
    Full_Adder FA_11205(s11205, c11205, in11205_1, in11205_2, s9004[0]);
    wire[0:0] s11206, in11206_1, in11206_2;
    wire c11206;
    assign in11206_1 = {s9008[0]};
    assign in11206_2 = {s9009[0]};
    Full_Adder FA_11206(s11206, c11206, in11206_1, in11206_2, s9007[0]);
    wire[0:0] s11207, in11207_1, in11207_2;
    wire c11207;
    assign in11207_1 = {c9000};
    assign in11207_2 = {c9001};
    Full_Adder FA_11207(s11207, c11207, in11207_1, in11207_2, c8999);
    wire[0:0] s11208, in11208_1, in11208_2;
    wire c11208;
    assign in11208_1 = {c9003};
    assign in11208_2 = {c9004};
    Full_Adder FA_11208(s11208, c11208, in11208_1, in11208_2, c9002);
    wire[0:0] s11209, in11209_1, in11209_2;
    wire c11209;
    assign in11209_1 = {c9006};
    assign in11209_2 = {c9007};
    Full_Adder FA_11209(s11209, c11209, in11209_1, in11209_2, c9005);
    wire[0:0] s11210, in11210_1, in11210_2;
    wire c11210;
    assign in11210_1 = {c9009};
    assign in11210_2 = {c9010};
    Full_Adder FA_11210(s11210, c11210, in11210_1, in11210_2, c9008);
    wire[0:0] s11211, in11211_1, in11211_2;
    wire c11211;
    assign in11211_1 = {s9012[0]};
    assign in11211_2 = {s9013[0]};
    Full_Adder FA_11211(s11211, c11211, in11211_1, in11211_2, c9011);
    wire[0:0] s11212, in11212_1, in11212_2;
    wire c11212;
    assign in11212_1 = {s9015[0]};
    assign in11212_2 = {s9016[0]};
    Full_Adder FA_11212(s11212, c11212, in11212_1, in11212_2, s9014[0]);
    wire[0:0] s11213, in11213_1, in11213_2;
    wire c11213;
    assign in11213_1 = {s9018[0]};
    assign in11213_2 = {s9019[0]};
    Full_Adder FA_11213(s11213, c11213, in11213_1, in11213_2, s9017[0]);
    wire[0:0] s11214, in11214_1, in11214_2;
    wire c11214;
    assign in11214_1 = {s9021[0]};
    assign in11214_2 = {s9022[0]};
    Full_Adder FA_11214(s11214, c11214, in11214_1, in11214_2, s9020[0]);
    wire[0:0] s11215, in11215_1, in11215_2;
    wire c11215;
    assign in11215_1 = {c9013};
    assign in11215_2 = {c9014};
    Full_Adder FA_11215(s11215, c11215, in11215_1, in11215_2, c9012);
    wire[0:0] s11216, in11216_1, in11216_2;
    wire c11216;
    assign in11216_1 = {c9016};
    assign in11216_2 = {c9017};
    Full_Adder FA_11216(s11216, c11216, in11216_1, in11216_2, c9015);
    wire[0:0] s11217, in11217_1, in11217_2;
    wire c11217;
    assign in11217_1 = {c9019};
    assign in11217_2 = {c9020};
    Full_Adder FA_11217(s11217, c11217, in11217_1, in11217_2, c9018);
    wire[0:0] s11218, in11218_1, in11218_2;
    wire c11218;
    assign in11218_1 = {c9022};
    assign in11218_2 = {c9023};
    Full_Adder FA_11218(s11218, c11218, in11218_1, in11218_2, c9021);
    wire[0:0] s11219, in11219_1, in11219_2;
    wire c11219;
    assign in11219_1 = {s9025[0]};
    assign in11219_2 = {s9026[0]};
    Full_Adder FA_11219(s11219, c11219, in11219_1, in11219_2, c9024);
    wire[0:0] s11220, in11220_1, in11220_2;
    wire c11220;
    assign in11220_1 = {s9028[0]};
    assign in11220_2 = {s9029[0]};
    Full_Adder FA_11220(s11220, c11220, in11220_1, in11220_2, s9027[0]);
    wire[0:0] s11221, in11221_1, in11221_2;
    wire c11221;
    assign in11221_1 = {s9031[0]};
    assign in11221_2 = {s9032[0]};
    Full_Adder FA_11221(s11221, c11221, in11221_1, in11221_2, s9030[0]);
    wire[0:0] s11222, in11222_1, in11222_2;
    wire c11222;
    assign in11222_1 = {s9034[0]};
    assign in11222_2 = {s9035[0]};
    Full_Adder FA_11222(s11222, c11222, in11222_1, in11222_2, s9033[0]);
    wire[0:0] s11223, in11223_1, in11223_2;
    wire c11223;
    assign in11223_1 = {c9026};
    assign in11223_2 = {c9027};
    Full_Adder FA_11223(s11223, c11223, in11223_1, in11223_2, c9025);
    wire[0:0] s11224, in11224_1, in11224_2;
    wire c11224;
    assign in11224_1 = {c9029};
    assign in11224_2 = {c9030};
    Full_Adder FA_11224(s11224, c11224, in11224_1, in11224_2, c9028);
    wire[0:0] s11225, in11225_1, in11225_2;
    wire c11225;
    assign in11225_1 = {c9032};
    assign in11225_2 = {c9033};
    Full_Adder FA_11225(s11225, c11225, in11225_1, in11225_2, c9031);
    wire[0:0] s11226, in11226_1, in11226_2;
    wire c11226;
    assign in11226_1 = {c9035};
    assign in11226_2 = {c9036};
    Full_Adder FA_11226(s11226, c11226, in11226_1, in11226_2, c9034);
    wire[0:0] s11227, in11227_1, in11227_2;
    wire c11227;
    assign in11227_1 = {s9038[0]};
    assign in11227_2 = {s9039[0]};
    Full_Adder FA_11227(s11227, c11227, in11227_1, in11227_2, c9037);
    wire[0:0] s11228, in11228_1, in11228_2;
    wire c11228;
    assign in11228_1 = {s9041[0]};
    assign in11228_2 = {s9042[0]};
    Full_Adder FA_11228(s11228, c11228, in11228_1, in11228_2, s9040[0]);
    wire[0:0] s11229, in11229_1, in11229_2;
    wire c11229;
    assign in11229_1 = {s9044[0]};
    assign in11229_2 = {s9045[0]};
    Full_Adder FA_11229(s11229, c11229, in11229_1, in11229_2, s9043[0]);
    wire[0:0] s11230, in11230_1, in11230_2;
    wire c11230;
    assign in11230_1 = {s9047[0]};
    assign in11230_2 = {s9048[0]};
    Full_Adder FA_11230(s11230, c11230, in11230_1, in11230_2, s9046[0]);
    wire[0:0] s11231, in11231_1, in11231_2;
    wire c11231;
    assign in11231_1 = {c9039};
    assign in11231_2 = {c9040};
    Full_Adder FA_11231(s11231, c11231, in11231_1, in11231_2, c9038);
    wire[0:0] s11232, in11232_1, in11232_2;
    wire c11232;
    assign in11232_1 = {c9042};
    assign in11232_2 = {c9043};
    Full_Adder FA_11232(s11232, c11232, in11232_1, in11232_2, c9041);
    wire[0:0] s11233, in11233_1, in11233_2;
    wire c11233;
    assign in11233_1 = {c9045};
    assign in11233_2 = {c9046};
    Full_Adder FA_11233(s11233, c11233, in11233_1, in11233_2, c9044);
    wire[0:0] s11234, in11234_1, in11234_2;
    wire c11234;
    assign in11234_1 = {c9048};
    assign in11234_2 = {c9049};
    Full_Adder FA_11234(s11234, c11234, in11234_1, in11234_2, c9047);
    wire[0:0] s11235, in11235_1, in11235_2;
    wire c11235;
    assign in11235_1 = {s9051[0]};
    assign in11235_2 = {s9052[0]};
    Full_Adder FA_11235(s11235, c11235, in11235_1, in11235_2, c9050);
    wire[0:0] s11236, in11236_1, in11236_2;
    wire c11236;
    assign in11236_1 = {s9054[0]};
    assign in11236_2 = {s9055[0]};
    Full_Adder FA_11236(s11236, c11236, in11236_1, in11236_2, s9053[0]);
    wire[0:0] s11237, in11237_1, in11237_2;
    wire c11237;
    assign in11237_1 = {s9057[0]};
    assign in11237_2 = {s9058[0]};
    Full_Adder FA_11237(s11237, c11237, in11237_1, in11237_2, s9056[0]);
    wire[0:0] s11238, in11238_1, in11238_2;
    wire c11238;
    assign in11238_1 = {s9060[0]};
    assign in11238_2 = {s9061[0]};
    Full_Adder FA_11238(s11238, c11238, in11238_1, in11238_2, s9059[0]);
    wire[0:0] s11239, in11239_1, in11239_2;
    wire c11239;
    assign in11239_1 = {c9052};
    assign in11239_2 = {c9053};
    Full_Adder FA_11239(s11239, c11239, in11239_1, in11239_2, c9051);
    wire[0:0] s11240, in11240_1, in11240_2;
    wire c11240;
    assign in11240_1 = {c9055};
    assign in11240_2 = {c9056};
    Full_Adder FA_11240(s11240, c11240, in11240_1, in11240_2, c9054);
    wire[0:0] s11241, in11241_1, in11241_2;
    wire c11241;
    assign in11241_1 = {c9058};
    assign in11241_2 = {c9059};
    Full_Adder FA_11241(s11241, c11241, in11241_1, in11241_2, c9057);
    wire[0:0] s11242, in11242_1, in11242_2;
    wire c11242;
    assign in11242_1 = {c9061};
    assign in11242_2 = {c9062};
    Full_Adder FA_11242(s11242, c11242, in11242_1, in11242_2, c9060);
    wire[0:0] s11243, in11243_1, in11243_2;
    wire c11243;
    assign in11243_1 = {s9064[0]};
    assign in11243_2 = {s9065[0]};
    Full_Adder FA_11243(s11243, c11243, in11243_1, in11243_2, c9063);
    wire[0:0] s11244, in11244_1, in11244_2;
    wire c11244;
    assign in11244_1 = {s9067[0]};
    assign in11244_2 = {s9068[0]};
    Full_Adder FA_11244(s11244, c11244, in11244_1, in11244_2, s9066[0]);
    wire[0:0] s11245, in11245_1, in11245_2;
    wire c11245;
    assign in11245_1 = {s9070[0]};
    assign in11245_2 = {s9071[0]};
    Full_Adder FA_11245(s11245, c11245, in11245_1, in11245_2, s9069[0]);
    wire[0:0] s11246, in11246_1, in11246_2;
    wire c11246;
    assign in11246_1 = {s9073[0]};
    assign in11246_2 = {s9074[0]};
    Full_Adder FA_11246(s11246, c11246, in11246_1, in11246_2, s9072[0]);
    wire[0:0] s11247, in11247_1, in11247_2;
    wire c11247;
    assign in11247_1 = {c9065};
    assign in11247_2 = {c9066};
    Full_Adder FA_11247(s11247, c11247, in11247_1, in11247_2, c9064);
    wire[0:0] s11248, in11248_1, in11248_2;
    wire c11248;
    assign in11248_1 = {c9068};
    assign in11248_2 = {c9069};
    Full_Adder FA_11248(s11248, c11248, in11248_1, in11248_2, c9067);
    wire[0:0] s11249, in11249_1, in11249_2;
    wire c11249;
    assign in11249_1 = {c9071};
    assign in11249_2 = {c9072};
    Full_Adder FA_11249(s11249, c11249, in11249_1, in11249_2, c9070);
    wire[0:0] s11250, in11250_1, in11250_2;
    wire c11250;
    assign in11250_1 = {c9074};
    assign in11250_2 = {c9075};
    Full_Adder FA_11250(s11250, c11250, in11250_1, in11250_2, c9073);
    wire[0:0] s11251, in11251_1, in11251_2;
    wire c11251;
    assign in11251_1 = {s9077[0]};
    assign in11251_2 = {s9078[0]};
    Full_Adder FA_11251(s11251, c11251, in11251_1, in11251_2, c9076);
    wire[0:0] s11252, in11252_1, in11252_2;
    wire c11252;
    assign in11252_1 = {s9080[0]};
    assign in11252_2 = {s9081[0]};
    Full_Adder FA_11252(s11252, c11252, in11252_1, in11252_2, s9079[0]);
    wire[0:0] s11253, in11253_1, in11253_2;
    wire c11253;
    assign in11253_1 = {s9083[0]};
    assign in11253_2 = {s9084[0]};
    Full_Adder FA_11253(s11253, c11253, in11253_1, in11253_2, s9082[0]);
    wire[0:0] s11254, in11254_1, in11254_2;
    wire c11254;
    assign in11254_1 = {s9086[0]};
    assign in11254_2 = {s9087[0]};
    Full_Adder FA_11254(s11254, c11254, in11254_1, in11254_2, s9085[0]);
    wire[0:0] s11255, in11255_1, in11255_2;
    wire c11255;
    assign in11255_1 = {c9078};
    assign in11255_2 = {c9079};
    Full_Adder FA_11255(s11255, c11255, in11255_1, in11255_2, c9077);
    wire[0:0] s11256, in11256_1, in11256_2;
    wire c11256;
    assign in11256_1 = {c9081};
    assign in11256_2 = {c9082};
    Full_Adder FA_11256(s11256, c11256, in11256_1, in11256_2, c9080);
    wire[0:0] s11257, in11257_1, in11257_2;
    wire c11257;
    assign in11257_1 = {c9084};
    assign in11257_2 = {c9085};
    Full_Adder FA_11257(s11257, c11257, in11257_1, in11257_2, c9083);
    wire[0:0] s11258, in11258_1, in11258_2;
    wire c11258;
    assign in11258_1 = {c9087};
    assign in11258_2 = {c9088};
    Full_Adder FA_11258(s11258, c11258, in11258_1, in11258_2, c9086);
    wire[0:0] s11259, in11259_1, in11259_2;
    wire c11259;
    assign in11259_1 = {s9090[0]};
    assign in11259_2 = {s9091[0]};
    Full_Adder FA_11259(s11259, c11259, in11259_1, in11259_2, c9089);
    wire[0:0] s11260, in11260_1, in11260_2;
    wire c11260;
    assign in11260_1 = {s9093[0]};
    assign in11260_2 = {s9094[0]};
    Full_Adder FA_11260(s11260, c11260, in11260_1, in11260_2, s9092[0]);
    wire[0:0] s11261, in11261_1, in11261_2;
    wire c11261;
    assign in11261_1 = {s9096[0]};
    assign in11261_2 = {s9097[0]};
    Full_Adder FA_11261(s11261, c11261, in11261_1, in11261_2, s9095[0]);
    wire[0:0] s11262, in11262_1, in11262_2;
    wire c11262;
    assign in11262_1 = {s9099[0]};
    assign in11262_2 = {s9100[0]};
    Full_Adder FA_11262(s11262, c11262, in11262_1, in11262_2, s9098[0]);
    wire[0:0] s11263, in11263_1, in11263_2;
    wire c11263;
    assign in11263_1 = {c9091};
    assign in11263_2 = {c9092};
    Full_Adder FA_11263(s11263, c11263, in11263_1, in11263_2, c9090);
    wire[0:0] s11264, in11264_1, in11264_2;
    wire c11264;
    assign in11264_1 = {c9094};
    assign in11264_2 = {c9095};
    Full_Adder FA_11264(s11264, c11264, in11264_1, in11264_2, c9093);
    wire[0:0] s11265, in11265_1, in11265_2;
    wire c11265;
    assign in11265_1 = {c9097};
    assign in11265_2 = {c9098};
    Full_Adder FA_11265(s11265, c11265, in11265_1, in11265_2, c9096);
    wire[0:0] s11266, in11266_1, in11266_2;
    wire c11266;
    assign in11266_1 = {c9100};
    assign in11266_2 = {c9101};
    Full_Adder FA_11266(s11266, c11266, in11266_1, in11266_2, c9099);
    wire[0:0] s11267, in11267_1, in11267_2;
    wire c11267;
    assign in11267_1 = {s9103[0]};
    assign in11267_2 = {s9104[0]};
    Full_Adder FA_11267(s11267, c11267, in11267_1, in11267_2, c9102);
    wire[0:0] s11268, in11268_1, in11268_2;
    wire c11268;
    assign in11268_1 = {s9106[0]};
    assign in11268_2 = {s9107[0]};
    Full_Adder FA_11268(s11268, c11268, in11268_1, in11268_2, s9105[0]);
    wire[0:0] s11269, in11269_1, in11269_2;
    wire c11269;
    assign in11269_1 = {s9109[0]};
    assign in11269_2 = {s9110[0]};
    Full_Adder FA_11269(s11269, c11269, in11269_1, in11269_2, s9108[0]);
    wire[0:0] s11270, in11270_1, in11270_2;
    wire c11270;
    assign in11270_1 = {s9112[0]};
    assign in11270_2 = {s9113[0]};
    Full_Adder FA_11270(s11270, c11270, in11270_1, in11270_2, s9111[0]);
    wire[0:0] s11271, in11271_1, in11271_2;
    wire c11271;
    assign in11271_1 = {c9104};
    assign in11271_2 = {c9105};
    Full_Adder FA_11271(s11271, c11271, in11271_1, in11271_2, c9103);
    wire[0:0] s11272, in11272_1, in11272_2;
    wire c11272;
    assign in11272_1 = {c9107};
    assign in11272_2 = {c9108};
    Full_Adder FA_11272(s11272, c11272, in11272_1, in11272_2, c9106);
    wire[0:0] s11273, in11273_1, in11273_2;
    wire c11273;
    assign in11273_1 = {c9110};
    assign in11273_2 = {c9111};
    Full_Adder FA_11273(s11273, c11273, in11273_1, in11273_2, c9109);
    wire[0:0] s11274, in11274_1, in11274_2;
    wire c11274;
    assign in11274_1 = {c9113};
    assign in11274_2 = {c9114};
    Full_Adder FA_11274(s11274, c11274, in11274_1, in11274_2, c9112);
    wire[0:0] s11275, in11275_1, in11275_2;
    wire c11275;
    assign in11275_1 = {s9116[0]};
    assign in11275_2 = {s9117[0]};
    Full_Adder FA_11275(s11275, c11275, in11275_1, in11275_2, c9115);
    wire[0:0] s11276, in11276_1, in11276_2;
    wire c11276;
    assign in11276_1 = {s9119[0]};
    assign in11276_2 = {s9120[0]};
    Full_Adder FA_11276(s11276, c11276, in11276_1, in11276_2, s9118[0]);
    wire[0:0] s11277, in11277_1, in11277_2;
    wire c11277;
    assign in11277_1 = {s9122[0]};
    assign in11277_2 = {s9123[0]};
    Full_Adder FA_11277(s11277, c11277, in11277_1, in11277_2, s9121[0]);
    wire[0:0] s11278, in11278_1, in11278_2;
    wire c11278;
    assign in11278_1 = {s9125[0]};
    assign in11278_2 = {s9126[0]};
    Full_Adder FA_11278(s11278, c11278, in11278_1, in11278_2, s9124[0]);
    wire[0:0] s11279, in11279_1, in11279_2;
    wire c11279;
    assign in11279_1 = {c9117};
    assign in11279_2 = {c9118};
    Full_Adder FA_11279(s11279, c11279, in11279_1, in11279_2, c9116);
    wire[0:0] s11280, in11280_1, in11280_2;
    wire c11280;
    assign in11280_1 = {c9120};
    assign in11280_2 = {c9121};
    Full_Adder FA_11280(s11280, c11280, in11280_1, in11280_2, c9119);
    wire[0:0] s11281, in11281_1, in11281_2;
    wire c11281;
    assign in11281_1 = {c9123};
    assign in11281_2 = {c9124};
    Full_Adder FA_11281(s11281, c11281, in11281_1, in11281_2, c9122);
    wire[0:0] s11282, in11282_1, in11282_2;
    wire c11282;
    assign in11282_1 = {c9126};
    assign in11282_2 = {c9127};
    Full_Adder FA_11282(s11282, c11282, in11282_1, in11282_2, c9125);
    wire[0:0] s11283, in11283_1, in11283_2;
    wire c11283;
    assign in11283_1 = {s9129[0]};
    assign in11283_2 = {s9130[0]};
    Full_Adder FA_11283(s11283, c11283, in11283_1, in11283_2, c9128);
    wire[0:0] s11284, in11284_1, in11284_2;
    wire c11284;
    assign in11284_1 = {s9132[0]};
    assign in11284_2 = {s9133[0]};
    Full_Adder FA_11284(s11284, c11284, in11284_1, in11284_2, s9131[0]);
    wire[0:0] s11285, in11285_1, in11285_2;
    wire c11285;
    assign in11285_1 = {s9135[0]};
    assign in11285_2 = {s9136[0]};
    Full_Adder FA_11285(s11285, c11285, in11285_1, in11285_2, s9134[0]);
    wire[0:0] s11286, in11286_1, in11286_2;
    wire c11286;
    assign in11286_1 = {s9138[0]};
    assign in11286_2 = {s9139[0]};
    Full_Adder FA_11286(s11286, c11286, in11286_1, in11286_2, s9137[0]);
    wire[0:0] s11287, in11287_1, in11287_2;
    wire c11287;
    assign in11287_1 = {c9130};
    assign in11287_2 = {c9131};
    Full_Adder FA_11287(s11287, c11287, in11287_1, in11287_2, c9129);
    wire[0:0] s11288, in11288_1, in11288_2;
    wire c11288;
    assign in11288_1 = {c9133};
    assign in11288_2 = {c9134};
    Full_Adder FA_11288(s11288, c11288, in11288_1, in11288_2, c9132);
    wire[0:0] s11289, in11289_1, in11289_2;
    wire c11289;
    assign in11289_1 = {c9136};
    assign in11289_2 = {c9137};
    Full_Adder FA_11289(s11289, c11289, in11289_1, in11289_2, c9135);
    wire[0:0] s11290, in11290_1, in11290_2;
    wire c11290;
    assign in11290_1 = {c9139};
    assign in11290_2 = {c9140};
    Full_Adder FA_11290(s11290, c11290, in11290_1, in11290_2, c9138);
    wire[0:0] s11291, in11291_1, in11291_2;
    wire c11291;
    assign in11291_1 = {s9142[0]};
    assign in11291_2 = {s9143[0]};
    Full_Adder FA_11291(s11291, c11291, in11291_1, in11291_2, c9141);
    wire[0:0] s11292, in11292_1, in11292_2;
    wire c11292;
    assign in11292_1 = {s9145[0]};
    assign in11292_2 = {s9146[0]};
    Full_Adder FA_11292(s11292, c11292, in11292_1, in11292_2, s9144[0]);
    wire[0:0] s11293, in11293_1, in11293_2;
    wire c11293;
    assign in11293_1 = {s9148[0]};
    assign in11293_2 = {s9149[0]};
    Full_Adder FA_11293(s11293, c11293, in11293_1, in11293_2, s9147[0]);
    wire[0:0] s11294, in11294_1, in11294_2;
    wire c11294;
    assign in11294_1 = {s9151[0]};
    assign in11294_2 = {s9152[0]};
    Full_Adder FA_11294(s11294, c11294, in11294_1, in11294_2, s9150[0]);
    wire[0:0] s11295, in11295_1, in11295_2;
    wire c11295;
    assign in11295_1 = {c9143};
    assign in11295_2 = {c9144};
    Full_Adder FA_11295(s11295, c11295, in11295_1, in11295_2, c9142);
    wire[0:0] s11296, in11296_1, in11296_2;
    wire c11296;
    assign in11296_1 = {c9146};
    assign in11296_2 = {c9147};
    Full_Adder FA_11296(s11296, c11296, in11296_1, in11296_2, c9145);
    wire[0:0] s11297, in11297_1, in11297_2;
    wire c11297;
    assign in11297_1 = {c9149};
    assign in11297_2 = {c9150};
    Full_Adder FA_11297(s11297, c11297, in11297_1, in11297_2, c9148);
    wire[0:0] s11298, in11298_1, in11298_2;
    wire c11298;
    assign in11298_1 = {c9152};
    assign in11298_2 = {c9153};
    Full_Adder FA_11298(s11298, c11298, in11298_1, in11298_2, c9151);
    wire[0:0] s11299, in11299_1, in11299_2;
    wire c11299;
    assign in11299_1 = {s9155[0]};
    assign in11299_2 = {s9156[0]};
    Full_Adder FA_11299(s11299, c11299, in11299_1, in11299_2, c9154);
    wire[0:0] s11300, in11300_1, in11300_2;
    wire c11300;
    assign in11300_1 = {s9158[0]};
    assign in11300_2 = {s9159[0]};
    Full_Adder FA_11300(s11300, c11300, in11300_1, in11300_2, s9157[0]);
    wire[0:0] s11301, in11301_1, in11301_2;
    wire c11301;
    assign in11301_1 = {s9161[0]};
    assign in11301_2 = {s9162[0]};
    Full_Adder FA_11301(s11301, c11301, in11301_1, in11301_2, s9160[0]);
    wire[0:0] s11302, in11302_1, in11302_2;
    wire c11302;
    assign in11302_1 = {s9164[0]};
    assign in11302_2 = {s9165[0]};
    Full_Adder FA_11302(s11302, c11302, in11302_1, in11302_2, s9163[0]);
    wire[0:0] s11303, in11303_1, in11303_2;
    wire c11303;
    assign in11303_1 = {c9156};
    assign in11303_2 = {c9157};
    Full_Adder FA_11303(s11303, c11303, in11303_1, in11303_2, c9155);
    wire[0:0] s11304, in11304_1, in11304_2;
    wire c11304;
    assign in11304_1 = {c9159};
    assign in11304_2 = {c9160};
    Full_Adder FA_11304(s11304, c11304, in11304_1, in11304_2, c9158);
    wire[0:0] s11305, in11305_1, in11305_2;
    wire c11305;
    assign in11305_1 = {c9162};
    assign in11305_2 = {c9163};
    Full_Adder FA_11305(s11305, c11305, in11305_1, in11305_2, c9161);
    wire[0:0] s11306, in11306_1, in11306_2;
    wire c11306;
    assign in11306_1 = {c9165};
    assign in11306_2 = {c9166};
    Full_Adder FA_11306(s11306, c11306, in11306_1, in11306_2, c9164);
    wire[0:0] s11307, in11307_1, in11307_2;
    wire c11307;
    assign in11307_1 = {s9168[0]};
    assign in11307_2 = {s9169[0]};
    Full_Adder FA_11307(s11307, c11307, in11307_1, in11307_2, c9167);
    wire[0:0] s11308, in11308_1, in11308_2;
    wire c11308;
    assign in11308_1 = {s9171[0]};
    assign in11308_2 = {s9172[0]};
    Full_Adder FA_11308(s11308, c11308, in11308_1, in11308_2, s9170[0]);
    wire[0:0] s11309, in11309_1, in11309_2;
    wire c11309;
    assign in11309_1 = {s9174[0]};
    assign in11309_2 = {s9175[0]};
    Full_Adder FA_11309(s11309, c11309, in11309_1, in11309_2, s9173[0]);
    wire[0:0] s11310, in11310_1, in11310_2;
    wire c11310;
    assign in11310_1 = {s9177[0]};
    assign in11310_2 = {s9178[0]};
    Full_Adder FA_11310(s11310, c11310, in11310_1, in11310_2, s9176[0]);
    wire[0:0] s11311, in11311_1, in11311_2;
    wire c11311;
    assign in11311_1 = {c9169};
    assign in11311_2 = {c9170};
    Full_Adder FA_11311(s11311, c11311, in11311_1, in11311_2, c9168);
    wire[0:0] s11312, in11312_1, in11312_2;
    wire c11312;
    assign in11312_1 = {c9172};
    assign in11312_2 = {c9173};
    Full_Adder FA_11312(s11312, c11312, in11312_1, in11312_2, c9171);
    wire[0:0] s11313, in11313_1, in11313_2;
    wire c11313;
    assign in11313_1 = {c9175};
    assign in11313_2 = {c9176};
    Full_Adder FA_11313(s11313, c11313, in11313_1, in11313_2, c9174);
    wire[0:0] s11314, in11314_1, in11314_2;
    wire c11314;
    assign in11314_1 = {c9178};
    assign in11314_2 = {c9179};
    Full_Adder FA_11314(s11314, c11314, in11314_1, in11314_2, c9177);
    wire[0:0] s11315, in11315_1, in11315_2;
    wire c11315;
    assign in11315_1 = {s9181[0]};
    assign in11315_2 = {s9182[0]};
    Full_Adder FA_11315(s11315, c11315, in11315_1, in11315_2, c9180);
    wire[0:0] s11316, in11316_1, in11316_2;
    wire c11316;
    assign in11316_1 = {s9184[0]};
    assign in11316_2 = {s9185[0]};
    Full_Adder FA_11316(s11316, c11316, in11316_1, in11316_2, s9183[0]);
    wire[0:0] s11317, in11317_1, in11317_2;
    wire c11317;
    assign in11317_1 = {s9187[0]};
    assign in11317_2 = {s9188[0]};
    Full_Adder FA_11317(s11317, c11317, in11317_1, in11317_2, s9186[0]);
    wire[0:0] s11318, in11318_1, in11318_2;
    wire c11318;
    assign in11318_1 = {s9190[0]};
    assign in11318_2 = {s9191[0]};
    Full_Adder FA_11318(s11318, c11318, in11318_1, in11318_2, s9189[0]);
    wire[0:0] s11319, in11319_1, in11319_2;
    wire c11319;
    assign in11319_1 = {c9182};
    assign in11319_2 = {c9183};
    Full_Adder FA_11319(s11319, c11319, in11319_1, in11319_2, c9181);
    wire[0:0] s11320, in11320_1, in11320_2;
    wire c11320;
    assign in11320_1 = {c9185};
    assign in11320_2 = {c9186};
    Full_Adder FA_11320(s11320, c11320, in11320_1, in11320_2, c9184);
    wire[0:0] s11321, in11321_1, in11321_2;
    wire c11321;
    assign in11321_1 = {c9188};
    assign in11321_2 = {c9189};
    Full_Adder FA_11321(s11321, c11321, in11321_1, in11321_2, c9187);
    wire[0:0] s11322, in11322_1, in11322_2;
    wire c11322;
    assign in11322_1 = {c9191};
    assign in11322_2 = {c9192};
    Full_Adder FA_11322(s11322, c11322, in11322_1, in11322_2, c9190);
    wire[0:0] s11323, in11323_1, in11323_2;
    wire c11323;
    assign in11323_1 = {s9194[0]};
    assign in11323_2 = {s9195[0]};
    Full_Adder FA_11323(s11323, c11323, in11323_1, in11323_2, c9193);
    wire[0:0] s11324, in11324_1, in11324_2;
    wire c11324;
    assign in11324_1 = {s9197[0]};
    assign in11324_2 = {s9198[0]};
    Full_Adder FA_11324(s11324, c11324, in11324_1, in11324_2, s9196[0]);
    wire[0:0] s11325, in11325_1, in11325_2;
    wire c11325;
    assign in11325_1 = {s9200[0]};
    assign in11325_2 = {s9201[0]};
    Full_Adder FA_11325(s11325, c11325, in11325_1, in11325_2, s9199[0]);
    wire[0:0] s11326, in11326_1, in11326_2;
    wire c11326;
    assign in11326_1 = {s9203[0]};
    assign in11326_2 = {s9204[0]};
    Full_Adder FA_11326(s11326, c11326, in11326_1, in11326_2, s9202[0]);
    wire[0:0] s11327, in11327_1, in11327_2;
    wire c11327;
    assign in11327_1 = {c9195};
    assign in11327_2 = {c9196};
    Full_Adder FA_11327(s11327, c11327, in11327_1, in11327_2, c9194);
    wire[0:0] s11328, in11328_1, in11328_2;
    wire c11328;
    assign in11328_1 = {c9198};
    assign in11328_2 = {c9199};
    Full_Adder FA_11328(s11328, c11328, in11328_1, in11328_2, c9197);
    wire[0:0] s11329, in11329_1, in11329_2;
    wire c11329;
    assign in11329_1 = {c9201};
    assign in11329_2 = {c9202};
    Full_Adder FA_11329(s11329, c11329, in11329_1, in11329_2, c9200);
    wire[0:0] s11330, in11330_1, in11330_2;
    wire c11330;
    assign in11330_1 = {c9204};
    assign in11330_2 = {c9205};
    Full_Adder FA_11330(s11330, c11330, in11330_1, in11330_2, c9203);
    wire[0:0] s11331, in11331_1, in11331_2;
    wire c11331;
    assign in11331_1 = {s9207[0]};
    assign in11331_2 = {s9208[0]};
    Full_Adder FA_11331(s11331, c11331, in11331_1, in11331_2, c9206);
    wire[0:0] s11332, in11332_1, in11332_2;
    wire c11332;
    assign in11332_1 = {s9210[0]};
    assign in11332_2 = {s9211[0]};
    Full_Adder FA_11332(s11332, c11332, in11332_1, in11332_2, s9209[0]);
    wire[0:0] s11333, in11333_1, in11333_2;
    wire c11333;
    assign in11333_1 = {s9213[0]};
    assign in11333_2 = {s9214[0]};
    Full_Adder FA_11333(s11333, c11333, in11333_1, in11333_2, s9212[0]);
    wire[0:0] s11334, in11334_1, in11334_2;
    wire c11334;
    assign in11334_1 = {s9216[0]};
    assign in11334_2 = {s9217[0]};
    Full_Adder FA_11334(s11334, c11334, in11334_1, in11334_2, s9215[0]);
    wire[0:0] s11335, in11335_1, in11335_2;
    wire c11335;
    assign in11335_1 = {c9208};
    assign in11335_2 = {c9209};
    Full_Adder FA_11335(s11335, c11335, in11335_1, in11335_2, c9207);
    wire[0:0] s11336, in11336_1, in11336_2;
    wire c11336;
    assign in11336_1 = {c9211};
    assign in11336_2 = {c9212};
    Full_Adder FA_11336(s11336, c11336, in11336_1, in11336_2, c9210);
    wire[0:0] s11337, in11337_1, in11337_2;
    wire c11337;
    assign in11337_1 = {c9214};
    assign in11337_2 = {c9215};
    Full_Adder FA_11337(s11337, c11337, in11337_1, in11337_2, c9213);
    wire[0:0] s11338, in11338_1, in11338_2;
    wire c11338;
    assign in11338_1 = {c9217};
    assign in11338_2 = {c9218};
    Full_Adder FA_11338(s11338, c11338, in11338_1, in11338_2, c9216);
    wire[0:0] s11339, in11339_1, in11339_2;
    wire c11339;
    assign in11339_1 = {s9220[0]};
    assign in11339_2 = {s9221[0]};
    Full_Adder FA_11339(s11339, c11339, in11339_1, in11339_2, c9219);
    wire[0:0] s11340, in11340_1, in11340_2;
    wire c11340;
    assign in11340_1 = {s9223[0]};
    assign in11340_2 = {s9224[0]};
    Full_Adder FA_11340(s11340, c11340, in11340_1, in11340_2, s9222[0]);
    wire[0:0] s11341, in11341_1, in11341_2;
    wire c11341;
    assign in11341_1 = {s9226[0]};
    assign in11341_2 = {s9227[0]};
    Full_Adder FA_11341(s11341, c11341, in11341_1, in11341_2, s9225[0]);
    wire[0:0] s11342, in11342_1, in11342_2;
    wire c11342;
    assign in11342_1 = {s9229[0]};
    assign in11342_2 = {s9230[0]};
    Full_Adder FA_11342(s11342, c11342, in11342_1, in11342_2, s9228[0]);
    wire[0:0] s11343, in11343_1, in11343_2;
    wire c11343;
    assign in11343_1 = {c9221};
    assign in11343_2 = {c9222};
    Full_Adder FA_11343(s11343, c11343, in11343_1, in11343_2, c9220);
    wire[0:0] s11344, in11344_1, in11344_2;
    wire c11344;
    assign in11344_1 = {c9224};
    assign in11344_2 = {c9225};
    Full_Adder FA_11344(s11344, c11344, in11344_1, in11344_2, c9223);
    wire[0:0] s11345, in11345_1, in11345_2;
    wire c11345;
    assign in11345_1 = {c9227};
    assign in11345_2 = {c9228};
    Full_Adder FA_11345(s11345, c11345, in11345_1, in11345_2, c9226);
    wire[0:0] s11346, in11346_1, in11346_2;
    wire c11346;
    assign in11346_1 = {c9230};
    assign in11346_2 = {c9231};
    Full_Adder FA_11346(s11346, c11346, in11346_1, in11346_2, c9229);
    wire[0:0] s11347, in11347_1, in11347_2;
    wire c11347;
    assign in11347_1 = {s9233[0]};
    assign in11347_2 = {s9234[0]};
    Full_Adder FA_11347(s11347, c11347, in11347_1, in11347_2, c9232);
    wire[0:0] s11348, in11348_1, in11348_2;
    wire c11348;
    assign in11348_1 = {s9236[0]};
    assign in11348_2 = {s9237[0]};
    Full_Adder FA_11348(s11348, c11348, in11348_1, in11348_2, s9235[0]);
    wire[0:0] s11349, in11349_1, in11349_2;
    wire c11349;
    assign in11349_1 = {s9239[0]};
    assign in11349_2 = {s9240[0]};
    Full_Adder FA_11349(s11349, c11349, in11349_1, in11349_2, s9238[0]);
    wire[0:0] s11350, in11350_1, in11350_2;
    wire c11350;
    assign in11350_1 = {s9242[0]};
    assign in11350_2 = {s9243[0]};
    Full_Adder FA_11350(s11350, c11350, in11350_1, in11350_2, s9241[0]);
    wire[0:0] s11351, in11351_1, in11351_2;
    wire c11351;
    assign in11351_1 = {c9234};
    assign in11351_2 = {c9235};
    Full_Adder FA_11351(s11351, c11351, in11351_1, in11351_2, c9233);
    wire[0:0] s11352, in11352_1, in11352_2;
    wire c11352;
    assign in11352_1 = {c9237};
    assign in11352_2 = {c9238};
    Full_Adder FA_11352(s11352, c11352, in11352_1, in11352_2, c9236);
    wire[0:0] s11353, in11353_1, in11353_2;
    wire c11353;
    assign in11353_1 = {c9240};
    assign in11353_2 = {c9241};
    Full_Adder FA_11353(s11353, c11353, in11353_1, in11353_2, c9239);
    wire[0:0] s11354, in11354_1, in11354_2;
    wire c11354;
    assign in11354_1 = {c9243};
    assign in11354_2 = {c9244};
    Full_Adder FA_11354(s11354, c11354, in11354_1, in11354_2, c9242);
    wire[0:0] s11355, in11355_1, in11355_2;
    wire c11355;
    assign in11355_1 = {s9246[0]};
    assign in11355_2 = {s9247[0]};
    Full_Adder FA_11355(s11355, c11355, in11355_1, in11355_2, c9245);
    wire[0:0] s11356, in11356_1, in11356_2;
    wire c11356;
    assign in11356_1 = {s9249[0]};
    assign in11356_2 = {s9250[0]};
    Full_Adder FA_11356(s11356, c11356, in11356_1, in11356_2, s9248[0]);
    wire[0:0] s11357, in11357_1, in11357_2;
    wire c11357;
    assign in11357_1 = {s9252[0]};
    assign in11357_2 = {s9253[0]};
    Full_Adder FA_11357(s11357, c11357, in11357_1, in11357_2, s9251[0]);
    wire[0:0] s11358, in11358_1, in11358_2;
    wire c11358;
    assign in11358_1 = {s9255[0]};
    assign in11358_2 = {s9256[0]};
    Full_Adder FA_11358(s11358, c11358, in11358_1, in11358_2, s9254[0]);
    wire[0:0] s11359, in11359_1, in11359_2;
    wire c11359;
    assign in11359_1 = {c9247};
    assign in11359_2 = {c9248};
    Full_Adder FA_11359(s11359, c11359, in11359_1, in11359_2, c9246);
    wire[0:0] s11360, in11360_1, in11360_2;
    wire c11360;
    assign in11360_1 = {c9250};
    assign in11360_2 = {c9251};
    Full_Adder FA_11360(s11360, c11360, in11360_1, in11360_2, c9249);
    wire[0:0] s11361, in11361_1, in11361_2;
    wire c11361;
    assign in11361_1 = {c9253};
    assign in11361_2 = {c9254};
    Full_Adder FA_11361(s11361, c11361, in11361_1, in11361_2, c9252);
    wire[0:0] s11362, in11362_1, in11362_2;
    wire c11362;
    assign in11362_1 = {c9256};
    assign in11362_2 = {c9257};
    Full_Adder FA_11362(s11362, c11362, in11362_1, in11362_2, c9255);
    wire[0:0] s11363, in11363_1, in11363_2;
    wire c11363;
    assign in11363_1 = {s9259[0]};
    assign in11363_2 = {s9260[0]};
    Full_Adder FA_11363(s11363, c11363, in11363_1, in11363_2, c9258);
    wire[0:0] s11364, in11364_1, in11364_2;
    wire c11364;
    assign in11364_1 = {s9262[0]};
    assign in11364_2 = {s9263[0]};
    Full_Adder FA_11364(s11364, c11364, in11364_1, in11364_2, s9261[0]);
    wire[0:0] s11365, in11365_1, in11365_2;
    wire c11365;
    assign in11365_1 = {s9265[0]};
    assign in11365_2 = {s9266[0]};
    Full_Adder FA_11365(s11365, c11365, in11365_1, in11365_2, s9264[0]);
    wire[0:0] s11366, in11366_1, in11366_2;
    wire c11366;
    assign in11366_1 = {s9268[0]};
    assign in11366_2 = {s9269[0]};
    Full_Adder FA_11366(s11366, c11366, in11366_1, in11366_2, s9267[0]);
    wire[0:0] s11367, in11367_1, in11367_2;
    wire c11367;
    assign in11367_1 = {c9260};
    assign in11367_2 = {c9261};
    Full_Adder FA_11367(s11367, c11367, in11367_1, in11367_2, c9259);
    wire[0:0] s11368, in11368_1, in11368_2;
    wire c11368;
    assign in11368_1 = {c9263};
    assign in11368_2 = {c9264};
    Full_Adder FA_11368(s11368, c11368, in11368_1, in11368_2, c9262);
    wire[0:0] s11369, in11369_1, in11369_2;
    wire c11369;
    assign in11369_1 = {c9266};
    assign in11369_2 = {c9267};
    Full_Adder FA_11369(s11369, c11369, in11369_1, in11369_2, c9265);
    wire[0:0] s11370, in11370_1, in11370_2;
    wire c11370;
    assign in11370_1 = {c9269};
    assign in11370_2 = {c9270};
    Full_Adder FA_11370(s11370, c11370, in11370_1, in11370_2, c9268);
    wire[0:0] s11371, in11371_1, in11371_2;
    wire c11371;
    assign in11371_1 = {s9272[0]};
    assign in11371_2 = {s9273[0]};
    Full_Adder FA_11371(s11371, c11371, in11371_1, in11371_2, c9271);
    wire[0:0] s11372, in11372_1, in11372_2;
    wire c11372;
    assign in11372_1 = {s9275[0]};
    assign in11372_2 = {s9276[0]};
    Full_Adder FA_11372(s11372, c11372, in11372_1, in11372_2, s9274[0]);
    wire[0:0] s11373, in11373_1, in11373_2;
    wire c11373;
    assign in11373_1 = {s9278[0]};
    assign in11373_2 = {s9279[0]};
    Full_Adder FA_11373(s11373, c11373, in11373_1, in11373_2, s9277[0]);
    wire[0:0] s11374, in11374_1, in11374_2;
    wire c11374;
    assign in11374_1 = {s9281[0]};
    assign in11374_2 = {s9282[0]};
    Full_Adder FA_11374(s11374, c11374, in11374_1, in11374_2, s9280[0]);
    wire[0:0] s11375, in11375_1, in11375_2;
    wire c11375;
    assign in11375_1 = {c9273};
    assign in11375_2 = {c9274};
    Full_Adder FA_11375(s11375, c11375, in11375_1, in11375_2, c9272);
    wire[0:0] s11376, in11376_1, in11376_2;
    wire c11376;
    assign in11376_1 = {c9276};
    assign in11376_2 = {c9277};
    Full_Adder FA_11376(s11376, c11376, in11376_1, in11376_2, c9275);
    wire[0:0] s11377, in11377_1, in11377_2;
    wire c11377;
    assign in11377_1 = {c9279};
    assign in11377_2 = {c9280};
    Full_Adder FA_11377(s11377, c11377, in11377_1, in11377_2, c9278);
    wire[0:0] s11378, in11378_1, in11378_2;
    wire c11378;
    assign in11378_1 = {c9282};
    assign in11378_2 = {c9283};
    Full_Adder FA_11378(s11378, c11378, in11378_1, in11378_2, c9281);
    wire[0:0] s11379, in11379_1, in11379_2;
    wire c11379;
    assign in11379_1 = {s9285[0]};
    assign in11379_2 = {s9286[0]};
    Full_Adder FA_11379(s11379, c11379, in11379_1, in11379_2, c9284);
    wire[0:0] s11380, in11380_1, in11380_2;
    wire c11380;
    assign in11380_1 = {s9288[0]};
    assign in11380_2 = {s9289[0]};
    Full_Adder FA_11380(s11380, c11380, in11380_1, in11380_2, s9287[0]);
    wire[0:0] s11381, in11381_1, in11381_2;
    wire c11381;
    assign in11381_1 = {s9291[0]};
    assign in11381_2 = {s9292[0]};
    Full_Adder FA_11381(s11381, c11381, in11381_1, in11381_2, s9290[0]);
    wire[0:0] s11382, in11382_1, in11382_2;
    wire c11382;
    assign in11382_1 = {s9294[0]};
    assign in11382_2 = {s9295[0]};
    Full_Adder FA_11382(s11382, c11382, in11382_1, in11382_2, s9293[0]);
    wire[0:0] s11383, in11383_1, in11383_2;
    wire c11383;
    assign in11383_1 = {c9286};
    assign in11383_2 = {c9287};
    Full_Adder FA_11383(s11383, c11383, in11383_1, in11383_2, c9285);
    wire[0:0] s11384, in11384_1, in11384_2;
    wire c11384;
    assign in11384_1 = {c9289};
    assign in11384_2 = {c9290};
    Full_Adder FA_11384(s11384, c11384, in11384_1, in11384_2, c9288);
    wire[0:0] s11385, in11385_1, in11385_2;
    wire c11385;
    assign in11385_1 = {c9292};
    assign in11385_2 = {c9293};
    Full_Adder FA_11385(s11385, c11385, in11385_1, in11385_2, c9291);
    wire[0:0] s11386, in11386_1, in11386_2;
    wire c11386;
    assign in11386_1 = {c9295};
    assign in11386_2 = {c9296};
    Full_Adder FA_11386(s11386, c11386, in11386_1, in11386_2, c9294);
    wire[0:0] s11387, in11387_1, in11387_2;
    wire c11387;
    assign in11387_1 = {s9298[0]};
    assign in11387_2 = {s9299[0]};
    Full_Adder FA_11387(s11387, c11387, in11387_1, in11387_2, c9297);
    wire[0:0] s11388, in11388_1, in11388_2;
    wire c11388;
    assign in11388_1 = {s9301[0]};
    assign in11388_2 = {s9302[0]};
    Full_Adder FA_11388(s11388, c11388, in11388_1, in11388_2, s9300[0]);
    wire[0:0] s11389, in11389_1, in11389_2;
    wire c11389;
    assign in11389_1 = {s9304[0]};
    assign in11389_2 = {s9305[0]};
    Full_Adder FA_11389(s11389, c11389, in11389_1, in11389_2, s9303[0]);
    wire[0:0] s11390, in11390_1, in11390_2;
    wire c11390;
    assign in11390_1 = {s9307[0]};
    assign in11390_2 = {s9308[0]};
    Full_Adder FA_11390(s11390, c11390, in11390_1, in11390_2, s9306[0]);
    wire[0:0] s11391, in11391_1, in11391_2;
    wire c11391;
    assign in11391_1 = {c9299};
    assign in11391_2 = {c9300};
    Full_Adder FA_11391(s11391, c11391, in11391_1, in11391_2, c9298);
    wire[0:0] s11392, in11392_1, in11392_2;
    wire c11392;
    assign in11392_1 = {c9302};
    assign in11392_2 = {c9303};
    Full_Adder FA_11392(s11392, c11392, in11392_1, in11392_2, c9301);
    wire[0:0] s11393, in11393_1, in11393_2;
    wire c11393;
    assign in11393_1 = {c9305};
    assign in11393_2 = {c9306};
    Full_Adder FA_11393(s11393, c11393, in11393_1, in11393_2, c9304);
    wire[0:0] s11394, in11394_1, in11394_2;
    wire c11394;
    assign in11394_1 = {c9308};
    assign in11394_2 = {c9309};
    Full_Adder FA_11394(s11394, c11394, in11394_1, in11394_2, c9307);
    wire[0:0] s11395, in11395_1, in11395_2;
    wire c11395;
    assign in11395_1 = {s9311[0]};
    assign in11395_2 = {s9312[0]};
    Full_Adder FA_11395(s11395, c11395, in11395_1, in11395_2, c9310);
    wire[0:0] s11396, in11396_1, in11396_2;
    wire c11396;
    assign in11396_1 = {s9314[0]};
    assign in11396_2 = {s9315[0]};
    Full_Adder FA_11396(s11396, c11396, in11396_1, in11396_2, s9313[0]);
    wire[0:0] s11397, in11397_1, in11397_2;
    wire c11397;
    assign in11397_1 = {s9317[0]};
    assign in11397_2 = {s9318[0]};
    Full_Adder FA_11397(s11397, c11397, in11397_1, in11397_2, s9316[0]);
    wire[0:0] s11398, in11398_1, in11398_2;
    wire c11398;
    assign in11398_1 = {s9320[0]};
    assign in11398_2 = {s9321[0]};
    Full_Adder FA_11398(s11398, c11398, in11398_1, in11398_2, s9319[0]);
    wire[0:0] s11399, in11399_1, in11399_2;
    wire c11399;
    assign in11399_1 = {c9312};
    assign in11399_2 = {c9313};
    Full_Adder FA_11399(s11399, c11399, in11399_1, in11399_2, c9311);
    wire[0:0] s11400, in11400_1, in11400_2;
    wire c11400;
    assign in11400_1 = {c9315};
    assign in11400_2 = {c9316};
    Full_Adder FA_11400(s11400, c11400, in11400_1, in11400_2, c9314);
    wire[0:0] s11401, in11401_1, in11401_2;
    wire c11401;
    assign in11401_1 = {c9318};
    assign in11401_2 = {c9319};
    Full_Adder FA_11401(s11401, c11401, in11401_1, in11401_2, c9317);
    wire[0:0] s11402, in11402_1, in11402_2;
    wire c11402;
    assign in11402_1 = {c9321};
    assign in11402_2 = {c9322};
    Full_Adder FA_11402(s11402, c11402, in11402_1, in11402_2, c9320);
    wire[0:0] s11403, in11403_1, in11403_2;
    wire c11403;
    assign in11403_1 = {s9324[0]};
    assign in11403_2 = {s9325[0]};
    Full_Adder FA_11403(s11403, c11403, in11403_1, in11403_2, c9323);
    wire[0:0] s11404, in11404_1, in11404_2;
    wire c11404;
    assign in11404_1 = {s9327[0]};
    assign in11404_2 = {s9328[0]};
    Full_Adder FA_11404(s11404, c11404, in11404_1, in11404_2, s9326[0]);
    wire[0:0] s11405, in11405_1, in11405_2;
    wire c11405;
    assign in11405_1 = {s9330[0]};
    assign in11405_2 = {s9331[0]};
    Full_Adder FA_11405(s11405, c11405, in11405_1, in11405_2, s9329[0]);
    wire[0:0] s11406, in11406_1, in11406_2;
    wire c11406;
    assign in11406_1 = {s9333[0]};
    assign in11406_2 = {s9334[0]};
    Full_Adder FA_11406(s11406, c11406, in11406_1, in11406_2, s9332[0]);
    wire[0:0] s11407, in11407_1, in11407_2;
    wire c11407;
    assign in11407_1 = {c9325};
    assign in11407_2 = {c9326};
    Full_Adder FA_11407(s11407, c11407, in11407_1, in11407_2, c9324);
    wire[0:0] s11408, in11408_1, in11408_2;
    wire c11408;
    assign in11408_1 = {c9328};
    assign in11408_2 = {c9329};
    Full_Adder FA_11408(s11408, c11408, in11408_1, in11408_2, c9327);
    wire[0:0] s11409, in11409_1, in11409_2;
    wire c11409;
    assign in11409_1 = {c9331};
    assign in11409_2 = {c9332};
    Full_Adder FA_11409(s11409, c11409, in11409_1, in11409_2, c9330);
    wire[0:0] s11410, in11410_1, in11410_2;
    wire c11410;
    assign in11410_1 = {c9334};
    assign in11410_2 = {c9335};
    Full_Adder FA_11410(s11410, c11410, in11410_1, in11410_2, c9333);
    wire[0:0] s11411, in11411_1, in11411_2;
    wire c11411;
    assign in11411_1 = {s9337[0]};
    assign in11411_2 = {s9338[0]};
    Full_Adder FA_11411(s11411, c11411, in11411_1, in11411_2, c9336);
    wire[0:0] s11412, in11412_1, in11412_2;
    wire c11412;
    assign in11412_1 = {s9340[0]};
    assign in11412_2 = {s9341[0]};
    Full_Adder FA_11412(s11412, c11412, in11412_1, in11412_2, s9339[0]);
    wire[0:0] s11413, in11413_1, in11413_2;
    wire c11413;
    assign in11413_1 = {s9343[0]};
    assign in11413_2 = {s9344[0]};
    Full_Adder FA_11413(s11413, c11413, in11413_1, in11413_2, s9342[0]);
    wire[0:0] s11414, in11414_1, in11414_2;
    wire c11414;
    assign in11414_1 = {s9346[0]};
    assign in11414_2 = {s9347[0]};
    Full_Adder FA_11414(s11414, c11414, in11414_1, in11414_2, s9345[0]);
    wire[0:0] s11415, in11415_1, in11415_2;
    wire c11415;
    assign in11415_1 = {c9338};
    assign in11415_2 = {c9339};
    Full_Adder FA_11415(s11415, c11415, in11415_1, in11415_2, c9337);
    wire[0:0] s11416, in11416_1, in11416_2;
    wire c11416;
    assign in11416_1 = {c9341};
    assign in11416_2 = {c9342};
    Full_Adder FA_11416(s11416, c11416, in11416_1, in11416_2, c9340);
    wire[0:0] s11417, in11417_1, in11417_2;
    wire c11417;
    assign in11417_1 = {c9344};
    assign in11417_2 = {c9345};
    Full_Adder FA_11417(s11417, c11417, in11417_1, in11417_2, c9343);
    wire[0:0] s11418, in11418_1, in11418_2;
    wire c11418;
    assign in11418_1 = {c9347};
    assign in11418_2 = {c9348};
    Full_Adder FA_11418(s11418, c11418, in11418_1, in11418_2, c9346);
    wire[0:0] s11419, in11419_1, in11419_2;
    wire c11419;
    assign in11419_1 = {s9350[0]};
    assign in11419_2 = {s9351[0]};
    Full_Adder FA_11419(s11419, c11419, in11419_1, in11419_2, c9349);
    wire[0:0] s11420, in11420_1, in11420_2;
    wire c11420;
    assign in11420_1 = {s9353[0]};
    assign in11420_2 = {s9354[0]};
    Full_Adder FA_11420(s11420, c11420, in11420_1, in11420_2, s9352[0]);
    wire[0:0] s11421, in11421_1, in11421_2;
    wire c11421;
    assign in11421_1 = {s9356[0]};
    assign in11421_2 = {s9357[0]};
    Full_Adder FA_11421(s11421, c11421, in11421_1, in11421_2, s9355[0]);
    wire[0:0] s11422, in11422_1, in11422_2;
    wire c11422;
    assign in11422_1 = {s9359[0]};
    assign in11422_2 = {s9360[0]};
    Full_Adder FA_11422(s11422, c11422, in11422_1, in11422_2, s9358[0]);
    wire[0:0] s11423, in11423_1, in11423_2;
    wire c11423;
    assign in11423_1 = {c9351};
    assign in11423_2 = {c9352};
    Full_Adder FA_11423(s11423, c11423, in11423_1, in11423_2, c9350);
    wire[0:0] s11424, in11424_1, in11424_2;
    wire c11424;
    assign in11424_1 = {c9354};
    assign in11424_2 = {c9355};
    Full_Adder FA_11424(s11424, c11424, in11424_1, in11424_2, c9353);
    wire[0:0] s11425, in11425_1, in11425_2;
    wire c11425;
    assign in11425_1 = {c9357};
    assign in11425_2 = {c9358};
    Full_Adder FA_11425(s11425, c11425, in11425_1, in11425_2, c9356);
    wire[0:0] s11426, in11426_1, in11426_2;
    wire c11426;
    assign in11426_1 = {c9360};
    assign in11426_2 = {c9361};
    Full_Adder FA_11426(s11426, c11426, in11426_1, in11426_2, c9359);
    wire[0:0] s11427, in11427_1, in11427_2;
    wire c11427;
    assign in11427_1 = {s9363[0]};
    assign in11427_2 = {s9364[0]};
    Full_Adder FA_11427(s11427, c11427, in11427_1, in11427_2, c9362);
    wire[0:0] s11428, in11428_1, in11428_2;
    wire c11428;
    assign in11428_1 = {s9366[0]};
    assign in11428_2 = {s9367[0]};
    Full_Adder FA_11428(s11428, c11428, in11428_1, in11428_2, s9365[0]);
    wire[0:0] s11429, in11429_1, in11429_2;
    wire c11429;
    assign in11429_1 = {s9369[0]};
    assign in11429_2 = {s9370[0]};
    Full_Adder FA_11429(s11429, c11429, in11429_1, in11429_2, s9368[0]);
    wire[0:0] s11430, in11430_1, in11430_2;
    wire c11430;
    assign in11430_1 = {s9372[0]};
    assign in11430_2 = {s9373[0]};
    Full_Adder FA_11430(s11430, c11430, in11430_1, in11430_2, s9371[0]);
    wire[0:0] s11431, in11431_1, in11431_2;
    wire c11431;
    assign in11431_1 = {c9364};
    assign in11431_2 = {c9365};
    Full_Adder FA_11431(s11431, c11431, in11431_1, in11431_2, c9363);
    wire[0:0] s11432, in11432_1, in11432_2;
    wire c11432;
    assign in11432_1 = {c9367};
    assign in11432_2 = {c9368};
    Full_Adder FA_11432(s11432, c11432, in11432_1, in11432_2, c9366);
    wire[0:0] s11433, in11433_1, in11433_2;
    wire c11433;
    assign in11433_1 = {c9370};
    assign in11433_2 = {c9371};
    Full_Adder FA_11433(s11433, c11433, in11433_1, in11433_2, c9369);
    wire[0:0] s11434, in11434_1, in11434_2;
    wire c11434;
    assign in11434_1 = {c9373};
    assign in11434_2 = {c9374};
    Full_Adder FA_11434(s11434, c11434, in11434_1, in11434_2, c9372);
    wire[0:0] s11435, in11435_1, in11435_2;
    wire c11435;
    assign in11435_1 = {s9376[0]};
    assign in11435_2 = {s9377[0]};
    Full_Adder FA_11435(s11435, c11435, in11435_1, in11435_2, c9375);
    wire[0:0] s11436, in11436_1, in11436_2;
    wire c11436;
    assign in11436_1 = {s9379[0]};
    assign in11436_2 = {s9380[0]};
    Full_Adder FA_11436(s11436, c11436, in11436_1, in11436_2, s9378[0]);
    wire[0:0] s11437, in11437_1, in11437_2;
    wire c11437;
    assign in11437_1 = {s9382[0]};
    assign in11437_2 = {s9383[0]};
    Full_Adder FA_11437(s11437, c11437, in11437_1, in11437_2, s9381[0]);
    wire[0:0] s11438, in11438_1, in11438_2;
    wire c11438;
    assign in11438_1 = {s9385[0]};
    assign in11438_2 = {s9386[0]};
    Full_Adder FA_11438(s11438, c11438, in11438_1, in11438_2, s9384[0]);
    wire[0:0] s11439, in11439_1, in11439_2;
    wire c11439;
    assign in11439_1 = {c9377};
    assign in11439_2 = {c9378};
    Full_Adder FA_11439(s11439, c11439, in11439_1, in11439_2, c9376);
    wire[0:0] s11440, in11440_1, in11440_2;
    wire c11440;
    assign in11440_1 = {c9380};
    assign in11440_2 = {c9381};
    Full_Adder FA_11440(s11440, c11440, in11440_1, in11440_2, c9379);
    wire[0:0] s11441, in11441_1, in11441_2;
    wire c11441;
    assign in11441_1 = {c9383};
    assign in11441_2 = {c9384};
    Full_Adder FA_11441(s11441, c11441, in11441_1, in11441_2, c9382);
    wire[0:0] s11442, in11442_1, in11442_2;
    wire c11442;
    assign in11442_1 = {c9386};
    assign in11442_2 = {c9387};
    Full_Adder FA_11442(s11442, c11442, in11442_1, in11442_2, c9385);
    wire[0:0] s11443, in11443_1, in11443_2;
    wire c11443;
    assign in11443_1 = {s9389[0]};
    assign in11443_2 = {s9390[0]};
    Full_Adder FA_11443(s11443, c11443, in11443_1, in11443_2, c9388);
    wire[0:0] s11444, in11444_1, in11444_2;
    wire c11444;
    assign in11444_1 = {s9392[0]};
    assign in11444_2 = {s9393[0]};
    Full_Adder FA_11444(s11444, c11444, in11444_1, in11444_2, s9391[0]);
    wire[0:0] s11445, in11445_1, in11445_2;
    wire c11445;
    assign in11445_1 = {s9395[0]};
    assign in11445_2 = {s9396[0]};
    Full_Adder FA_11445(s11445, c11445, in11445_1, in11445_2, s9394[0]);
    wire[0:0] s11446, in11446_1, in11446_2;
    wire c11446;
    assign in11446_1 = {s9398[0]};
    assign in11446_2 = {s9399[0]};
    Full_Adder FA_11446(s11446, c11446, in11446_1, in11446_2, s9397[0]);
    wire[0:0] s11447, in11447_1, in11447_2;
    wire c11447;
    assign in11447_1 = {c9390};
    assign in11447_2 = {c9391};
    Full_Adder FA_11447(s11447, c11447, in11447_1, in11447_2, c9389);
    wire[0:0] s11448, in11448_1, in11448_2;
    wire c11448;
    assign in11448_1 = {c9393};
    assign in11448_2 = {c9394};
    Full_Adder FA_11448(s11448, c11448, in11448_1, in11448_2, c9392);
    wire[0:0] s11449, in11449_1, in11449_2;
    wire c11449;
    assign in11449_1 = {c9396};
    assign in11449_2 = {c9397};
    Full_Adder FA_11449(s11449, c11449, in11449_1, in11449_2, c9395);
    wire[0:0] s11450, in11450_1, in11450_2;
    wire c11450;
    assign in11450_1 = {c9399};
    assign in11450_2 = {c9400};
    Full_Adder FA_11450(s11450, c11450, in11450_1, in11450_2, c9398);
    wire[0:0] s11451, in11451_1, in11451_2;
    wire c11451;
    assign in11451_1 = {s9402[0]};
    assign in11451_2 = {s9403[0]};
    Full_Adder FA_11451(s11451, c11451, in11451_1, in11451_2, c9401);
    wire[0:0] s11452, in11452_1, in11452_2;
    wire c11452;
    assign in11452_1 = {s9405[0]};
    assign in11452_2 = {s9406[0]};
    Full_Adder FA_11452(s11452, c11452, in11452_1, in11452_2, s9404[0]);
    wire[0:0] s11453, in11453_1, in11453_2;
    wire c11453;
    assign in11453_1 = {s9408[0]};
    assign in11453_2 = {s9409[0]};
    Full_Adder FA_11453(s11453, c11453, in11453_1, in11453_2, s9407[0]);
    wire[0:0] s11454, in11454_1, in11454_2;
    wire c11454;
    assign in11454_1 = {s9411[0]};
    assign in11454_2 = {s9412[0]};
    Full_Adder FA_11454(s11454, c11454, in11454_1, in11454_2, s9410[0]);
    wire[0:0] s11455, in11455_1, in11455_2;
    wire c11455;
    assign in11455_1 = {c9403};
    assign in11455_2 = {c9404};
    Full_Adder FA_11455(s11455, c11455, in11455_1, in11455_2, c9402);
    wire[0:0] s11456, in11456_1, in11456_2;
    wire c11456;
    assign in11456_1 = {c9406};
    assign in11456_2 = {c9407};
    Full_Adder FA_11456(s11456, c11456, in11456_1, in11456_2, c9405);
    wire[0:0] s11457, in11457_1, in11457_2;
    wire c11457;
    assign in11457_1 = {c9409};
    assign in11457_2 = {c9410};
    Full_Adder FA_11457(s11457, c11457, in11457_1, in11457_2, c9408);
    wire[0:0] s11458, in11458_1, in11458_2;
    wire c11458;
    assign in11458_1 = {c9412};
    assign in11458_2 = {c9413};
    Full_Adder FA_11458(s11458, c11458, in11458_1, in11458_2, c9411);
    wire[0:0] s11459, in11459_1, in11459_2;
    wire c11459;
    assign in11459_1 = {s9415[0]};
    assign in11459_2 = {s9416[0]};
    Full_Adder FA_11459(s11459, c11459, in11459_1, in11459_2, c9414);
    wire[0:0] s11460, in11460_1, in11460_2;
    wire c11460;
    assign in11460_1 = {s9418[0]};
    assign in11460_2 = {s9419[0]};
    Full_Adder FA_11460(s11460, c11460, in11460_1, in11460_2, s9417[0]);
    wire[0:0] s11461, in11461_1, in11461_2;
    wire c11461;
    assign in11461_1 = {s9421[0]};
    assign in11461_2 = {s9422[0]};
    Full_Adder FA_11461(s11461, c11461, in11461_1, in11461_2, s9420[0]);
    wire[0:0] s11462, in11462_1, in11462_2;
    wire c11462;
    assign in11462_1 = {s9424[0]};
    assign in11462_2 = {s9425[0]};
    Full_Adder FA_11462(s11462, c11462, in11462_1, in11462_2, s9423[0]);
    wire[0:0] s11463, in11463_1, in11463_2;
    wire c11463;
    assign in11463_1 = {c9416};
    assign in11463_2 = {c9417};
    Full_Adder FA_11463(s11463, c11463, in11463_1, in11463_2, c9415);
    wire[0:0] s11464, in11464_1, in11464_2;
    wire c11464;
    assign in11464_1 = {c9419};
    assign in11464_2 = {c9420};
    Full_Adder FA_11464(s11464, c11464, in11464_1, in11464_2, c9418);
    wire[0:0] s11465, in11465_1, in11465_2;
    wire c11465;
    assign in11465_1 = {c9422};
    assign in11465_2 = {c9423};
    Full_Adder FA_11465(s11465, c11465, in11465_1, in11465_2, c9421);
    wire[0:0] s11466, in11466_1, in11466_2;
    wire c11466;
    assign in11466_1 = {c9425};
    assign in11466_2 = {c9426};
    Full_Adder FA_11466(s11466, c11466, in11466_1, in11466_2, c9424);
    wire[0:0] s11467, in11467_1, in11467_2;
    wire c11467;
    assign in11467_1 = {s9428[0]};
    assign in11467_2 = {s9429[0]};
    Full_Adder FA_11467(s11467, c11467, in11467_1, in11467_2, c9427);
    wire[0:0] s11468, in11468_1, in11468_2;
    wire c11468;
    assign in11468_1 = {s9431[0]};
    assign in11468_2 = {s9432[0]};
    Full_Adder FA_11468(s11468, c11468, in11468_1, in11468_2, s9430[0]);
    wire[0:0] s11469, in11469_1, in11469_2;
    wire c11469;
    assign in11469_1 = {s9434[0]};
    assign in11469_2 = {s9435[0]};
    Full_Adder FA_11469(s11469, c11469, in11469_1, in11469_2, s9433[0]);
    wire[0:0] s11470, in11470_1, in11470_2;
    wire c11470;
    assign in11470_1 = {s9437[0]};
    assign in11470_2 = {s9438[0]};
    Full_Adder FA_11470(s11470, c11470, in11470_1, in11470_2, s9436[0]);
    wire[0:0] s11471, in11471_1, in11471_2;
    wire c11471;
    assign in11471_1 = {c9429};
    assign in11471_2 = {c9430};
    Full_Adder FA_11471(s11471, c11471, in11471_1, in11471_2, c9428);
    wire[0:0] s11472, in11472_1, in11472_2;
    wire c11472;
    assign in11472_1 = {c9432};
    assign in11472_2 = {c9433};
    Full_Adder FA_11472(s11472, c11472, in11472_1, in11472_2, c9431);
    wire[0:0] s11473, in11473_1, in11473_2;
    wire c11473;
    assign in11473_1 = {c9435};
    assign in11473_2 = {c9436};
    Full_Adder FA_11473(s11473, c11473, in11473_1, in11473_2, c9434);
    wire[0:0] s11474, in11474_1, in11474_2;
    wire c11474;
    assign in11474_1 = {c9438};
    assign in11474_2 = {c9439};
    Full_Adder FA_11474(s11474, c11474, in11474_1, in11474_2, c9437);
    wire[0:0] s11475, in11475_1, in11475_2;
    wire c11475;
    assign in11475_1 = {s9441[0]};
    assign in11475_2 = {s9442[0]};
    Full_Adder FA_11475(s11475, c11475, in11475_1, in11475_2, c9440);
    wire[0:0] s11476, in11476_1, in11476_2;
    wire c11476;
    assign in11476_1 = {s9444[0]};
    assign in11476_2 = {s9445[0]};
    Full_Adder FA_11476(s11476, c11476, in11476_1, in11476_2, s9443[0]);
    wire[0:0] s11477, in11477_1, in11477_2;
    wire c11477;
    assign in11477_1 = {s9447[0]};
    assign in11477_2 = {s9448[0]};
    Full_Adder FA_11477(s11477, c11477, in11477_1, in11477_2, s9446[0]);
    wire[0:0] s11478, in11478_1, in11478_2;
    wire c11478;
    assign in11478_1 = {s9450[0]};
    assign in11478_2 = {s9451[0]};
    Full_Adder FA_11478(s11478, c11478, in11478_1, in11478_2, s9449[0]);
    wire[0:0] s11479, in11479_1, in11479_2;
    wire c11479;
    assign in11479_1 = {c9442};
    assign in11479_2 = {c9443};
    Full_Adder FA_11479(s11479, c11479, in11479_1, in11479_2, c9441);
    wire[0:0] s11480, in11480_1, in11480_2;
    wire c11480;
    assign in11480_1 = {c9445};
    assign in11480_2 = {c9446};
    Full_Adder FA_11480(s11480, c11480, in11480_1, in11480_2, c9444);
    wire[0:0] s11481, in11481_1, in11481_2;
    wire c11481;
    assign in11481_1 = {c9448};
    assign in11481_2 = {c9449};
    Full_Adder FA_11481(s11481, c11481, in11481_1, in11481_2, c9447);
    wire[0:0] s11482, in11482_1, in11482_2;
    wire c11482;
    assign in11482_1 = {c9451};
    assign in11482_2 = {c9452};
    Full_Adder FA_11482(s11482, c11482, in11482_1, in11482_2, c9450);
    wire[0:0] s11483, in11483_1, in11483_2;
    wire c11483;
    assign in11483_1 = {s9454[0]};
    assign in11483_2 = {s9455[0]};
    Full_Adder FA_11483(s11483, c11483, in11483_1, in11483_2, c9453);
    wire[0:0] s11484, in11484_1, in11484_2;
    wire c11484;
    assign in11484_1 = {s9457[0]};
    assign in11484_2 = {s9458[0]};
    Full_Adder FA_11484(s11484, c11484, in11484_1, in11484_2, s9456[0]);
    wire[0:0] s11485, in11485_1, in11485_2;
    wire c11485;
    assign in11485_1 = {s9460[0]};
    assign in11485_2 = {s9461[0]};
    Full_Adder FA_11485(s11485, c11485, in11485_1, in11485_2, s9459[0]);
    wire[0:0] s11486, in11486_1, in11486_2;
    wire c11486;
    assign in11486_1 = {s9463[0]};
    assign in11486_2 = {s9464[0]};
    Full_Adder FA_11486(s11486, c11486, in11486_1, in11486_2, s9462[0]);
    wire[0:0] s11487, in11487_1, in11487_2;
    wire c11487;
    assign in11487_1 = {c9455};
    assign in11487_2 = {c9456};
    Full_Adder FA_11487(s11487, c11487, in11487_1, in11487_2, c9454);
    wire[0:0] s11488, in11488_1, in11488_2;
    wire c11488;
    assign in11488_1 = {c9458};
    assign in11488_2 = {c9459};
    Full_Adder FA_11488(s11488, c11488, in11488_1, in11488_2, c9457);
    wire[0:0] s11489, in11489_1, in11489_2;
    wire c11489;
    assign in11489_1 = {c9461};
    assign in11489_2 = {c9462};
    Full_Adder FA_11489(s11489, c11489, in11489_1, in11489_2, c9460);
    wire[0:0] s11490, in11490_1, in11490_2;
    wire c11490;
    assign in11490_1 = {c9464};
    assign in11490_2 = {c9465};
    Full_Adder FA_11490(s11490, c11490, in11490_1, in11490_2, c9463);
    wire[0:0] s11491, in11491_1, in11491_2;
    wire c11491;
    assign in11491_1 = {s9467[0]};
    assign in11491_2 = {s9468[0]};
    Full_Adder FA_11491(s11491, c11491, in11491_1, in11491_2, c9466);
    wire[0:0] s11492, in11492_1, in11492_2;
    wire c11492;
    assign in11492_1 = {s9470[0]};
    assign in11492_2 = {s9471[0]};
    Full_Adder FA_11492(s11492, c11492, in11492_1, in11492_2, s9469[0]);
    wire[0:0] s11493, in11493_1, in11493_2;
    wire c11493;
    assign in11493_1 = {s9473[0]};
    assign in11493_2 = {s9474[0]};
    Full_Adder FA_11493(s11493, c11493, in11493_1, in11493_2, s9472[0]);
    wire[0:0] s11494, in11494_1, in11494_2;
    wire c11494;
    assign in11494_1 = {s9476[0]};
    assign in11494_2 = {s9477[0]};
    Full_Adder FA_11494(s11494, c11494, in11494_1, in11494_2, s9475[0]);
    wire[0:0] s11495, in11495_1, in11495_2;
    wire c11495;
    assign in11495_1 = {c9468};
    assign in11495_2 = {c9469};
    Full_Adder FA_11495(s11495, c11495, in11495_1, in11495_2, c9467);
    wire[0:0] s11496, in11496_1, in11496_2;
    wire c11496;
    assign in11496_1 = {c9471};
    assign in11496_2 = {c9472};
    Full_Adder FA_11496(s11496, c11496, in11496_1, in11496_2, c9470);
    wire[0:0] s11497, in11497_1, in11497_2;
    wire c11497;
    assign in11497_1 = {c9474};
    assign in11497_2 = {c9475};
    Full_Adder FA_11497(s11497, c11497, in11497_1, in11497_2, c9473);
    wire[0:0] s11498, in11498_1, in11498_2;
    wire c11498;
    assign in11498_1 = {c9477};
    assign in11498_2 = {c9478};
    Full_Adder FA_11498(s11498, c11498, in11498_1, in11498_2, c9476);
    wire[0:0] s11499, in11499_1, in11499_2;
    wire c11499;
    assign in11499_1 = {s9480[0]};
    assign in11499_2 = {s9481[0]};
    Full_Adder FA_11499(s11499, c11499, in11499_1, in11499_2, c9479);
    wire[0:0] s11500, in11500_1, in11500_2;
    wire c11500;
    assign in11500_1 = {s9483[0]};
    assign in11500_2 = {s9484[0]};
    Full_Adder FA_11500(s11500, c11500, in11500_1, in11500_2, s9482[0]);
    wire[0:0] s11501, in11501_1, in11501_2;
    wire c11501;
    assign in11501_1 = {s9486[0]};
    assign in11501_2 = {s9487[0]};
    Full_Adder FA_11501(s11501, c11501, in11501_1, in11501_2, s9485[0]);
    wire[0:0] s11502, in11502_1, in11502_2;
    wire c11502;
    assign in11502_1 = {s9489[0]};
    assign in11502_2 = {s9490[0]};
    Full_Adder FA_11502(s11502, c11502, in11502_1, in11502_2, s9488[0]);
    wire[0:0] s11503, in11503_1, in11503_2;
    wire c11503;
    assign in11503_1 = {c9481};
    assign in11503_2 = {c9482};
    Full_Adder FA_11503(s11503, c11503, in11503_1, in11503_2, c9480);
    wire[0:0] s11504, in11504_1, in11504_2;
    wire c11504;
    assign in11504_1 = {c9484};
    assign in11504_2 = {c9485};
    Full_Adder FA_11504(s11504, c11504, in11504_1, in11504_2, c9483);
    wire[0:0] s11505, in11505_1, in11505_2;
    wire c11505;
    assign in11505_1 = {c9487};
    assign in11505_2 = {c9488};
    Full_Adder FA_11505(s11505, c11505, in11505_1, in11505_2, c9486);
    wire[0:0] s11506, in11506_1, in11506_2;
    wire c11506;
    assign in11506_1 = {c9490};
    assign in11506_2 = {c9491};
    Full_Adder FA_11506(s11506, c11506, in11506_1, in11506_2, c9489);
    wire[0:0] s11507, in11507_1, in11507_2;
    wire c11507;
    assign in11507_1 = {s9493[0]};
    assign in11507_2 = {s9494[0]};
    Full_Adder FA_11507(s11507, c11507, in11507_1, in11507_2, c9492);
    wire[0:0] s11508, in11508_1, in11508_2;
    wire c11508;
    assign in11508_1 = {s9496[0]};
    assign in11508_2 = {s9497[0]};
    Full_Adder FA_11508(s11508, c11508, in11508_1, in11508_2, s9495[0]);
    wire[0:0] s11509, in11509_1, in11509_2;
    wire c11509;
    assign in11509_1 = {s9499[0]};
    assign in11509_2 = {s9500[0]};
    Full_Adder FA_11509(s11509, c11509, in11509_1, in11509_2, s9498[0]);
    wire[0:0] s11510, in11510_1, in11510_2;
    wire c11510;
    assign in11510_1 = {s9502[0]};
    assign in11510_2 = {s9503[0]};
    Full_Adder FA_11510(s11510, c11510, in11510_1, in11510_2, s9501[0]);
    wire[0:0] s11511, in11511_1, in11511_2;
    wire c11511;
    assign in11511_1 = {c9494};
    assign in11511_2 = {c9495};
    Full_Adder FA_11511(s11511, c11511, in11511_1, in11511_2, c9493);
    wire[0:0] s11512, in11512_1, in11512_2;
    wire c11512;
    assign in11512_1 = {c9497};
    assign in11512_2 = {c9498};
    Full_Adder FA_11512(s11512, c11512, in11512_1, in11512_2, c9496);
    wire[0:0] s11513, in11513_1, in11513_2;
    wire c11513;
    assign in11513_1 = {c9500};
    assign in11513_2 = {c9501};
    Full_Adder FA_11513(s11513, c11513, in11513_1, in11513_2, c9499);
    wire[0:0] s11514, in11514_1, in11514_2;
    wire c11514;
    assign in11514_1 = {c9503};
    assign in11514_2 = {c9504};
    Full_Adder FA_11514(s11514, c11514, in11514_1, in11514_2, c9502);
    wire[0:0] s11515, in11515_1, in11515_2;
    wire c11515;
    assign in11515_1 = {s9506[0]};
    assign in11515_2 = {s9507[0]};
    Full_Adder FA_11515(s11515, c11515, in11515_1, in11515_2, c9505);
    wire[0:0] s11516, in11516_1, in11516_2;
    wire c11516;
    assign in11516_1 = {s9509[0]};
    assign in11516_2 = {s9510[0]};
    Full_Adder FA_11516(s11516, c11516, in11516_1, in11516_2, s9508[0]);
    wire[0:0] s11517, in11517_1, in11517_2;
    wire c11517;
    assign in11517_1 = {s9512[0]};
    assign in11517_2 = {s9513[0]};
    Full_Adder FA_11517(s11517, c11517, in11517_1, in11517_2, s9511[0]);
    wire[0:0] s11518, in11518_1, in11518_2;
    wire c11518;
    assign in11518_1 = {s9515[0]};
    assign in11518_2 = {s9516[0]};
    Full_Adder FA_11518(s11518, c11518, in11518_1, in11518_2, s9514[0]);
    wire[0:0] s11519, in11519_1, in11519_2;
    wire c11519;
    assign in11519_1 = {c9507};
    assign in11519_2 = {c9508};
    Full_Adder FA_11519(s11519, c11519, in11519_1, in11519_2, c9506);
    wire[0:0] s11520, in11520_1, in11520_2;
    wire c11520;
    assign in11520_1 = {c9510};
    assign in11520_2 = {c9511};
    Full_Adder FA_11520(s11520, c11520, in11520_1, in11520_2, c9509);
    wire[0:0] s11521, in11521_1, in11521_2;
    wire c11521;
    assign in11521_1 = {c9513};
    assign in11521_2 = {c9514};
    Full_Adder FA_11521(s11521, c11521, in11521_1, in11521_2, c9512);
    wire[0:0] s11522, in11522_1, in11522_2;
    wire c11522;
    assign in11522_1 = {c9516};
    assign in11522_2 = {c9517};
    Full_Adder FA_11522(s11522, c11522, in11522_1, in11522_2, c9515);
    wire[0:0] s11523, in11523_1, in11523_2;
    wire c11523;
    assign in11523_1 = {s9519[0]};
    assign in11523_2 = {s9520[0]};
    Full_Adder FA_11523(s11523, c11523, in11523_1, in11523_2, c9518);
    wire[0:0] s11524, in11524_1, in11524_2;
    wire c11524;
    assign in11524_1 = {s9522[0]};
    assign in11524_2 = {s9523[0]};
    Full_Adder FA_11524(s11524, c11524, in11524_1, in11524_2, s9521[0]);
    wire[0:0] s11525, in11525_1, in11525_2;
    wire c11525;
    assign in11525_1 = {s9525[0]};
    assign in11525_2 = {s9526[0]};
    Full_Adder FA_11525(s11525, c11525, in11525_1, in11525_2, s9524[0]);
    wire[0:0] s11526, in11526_1, in11526_2;
    wire c11526;
    assign in11526_1 = {s9528[0]};
    assign in11526_2 = {s9529[0]};
    Full_Adder FA_11526(s11526, c11526, in11526_1, in11526_2, s9527[0]);
    wire[0:0] s11527, in11527_1, in11527_2;
    wire c11527;
    assign in11527_1 = {c9520};
    assign in11527_2 = {c9521};
    Full_Adder FA_11527(s11527, c11527, in11527_1, in11527_2, c9519);
    wire[0:0] s11528, in11528_1, in11528_2;
    wire c11528;
    assign in11528_1 = {c9523};
    assign in11528_2 = {c9524};
    Full_Adder FA_11528(s11528, c11528, in11528_1, in11528_2, c9522);
    wire[0:0] s11529, in11529_1, in11529_2;
    wire c11529;
    assign in11529_1 = {c9526};
    assign in11529_2 = {c9527};
    Full_Adder FA_11529(s11529, c11529, in11529_1, in11529_2, c9525);
    wire[0:0] s11530, in11530_1, in11530_2;
    wire c11530;
    assign in11530_1 = {c9529};
    assign in11530_2 = {c9530};
    Full_Adder FA_11530(s11530, c11530, in11530_1, in11530_2, c9528);
    wire[0:0] s11531, in11531_1, in11531_2;
    wire c11531;
    assign in11531_1 = {s9532[0]};
    assign in11531_2 = {s9533[0]};
    Full_Adder FA_11531(s11531, c11531, in11531_1, in11531_2, c9531);
    wire[0:0] s11532, in11532_1, in11532_2;
    wire c11532;
    assign in11532_1 = {s9535[0]};
    assign in11532_2 = {s9536[0]};
    Full_Adder FA_11532(s11532, c11532, in11532_1, in11532_2, s9534[0]);
    wire[0:0] s11533, in11533_1, in11533_2;
    wire c11533;
    assign in11533_1 = {s9538[0]};
    assign in11533_2 = {s9539[0]};
    Full_Adder FA_11533(s11533, c11533, in11533_1, in11533_2, s9537[0]);
    wire[0:0] s11534, in11534_1, in11534_2;
    wire c11534;
    assign in11534_1 = {s9541[0]};
    assign in11534_2 = {s9542[0]};
    Full_Adder FA_11534(s11534, c11534, in11534_1, in11534_2, s9540[0]);
    wire[0:0] s11535, in11535_1, in11535_2;
    wire c11535;
    assign in11535_1 = {c9533};
    assign in11535_2 = {c9534};
    Full_Adder FA_11535(s11535, c11535, in11535_1, in11535_2, c9532);
    wire[0:0] s11536, in11536_1, in11536_2;
    wire c11536;
    assign in11536_1 = {c9536};
    assign in11536_2 = {c9537};
    Full_Adder FA_11536(s11536, c11536, in11536_1, in11536_2, c9535);
    wire[0:0] s11537, in11537_1, in11537_2;
    wire c11537;
    assign in11537_1 = {c9539};
    assign in11537_2 = {c9540};
    Full_Adder FA_11537(s11537, c11537, in11537_1, in11537_2, c9538);
    wire[0:0] s11538, in11538_1, in11538_2;
    wire c11538;
    assign in11538_1 = {c9542};
    assign in11538_2 = {c9543};
    Full_Adder FA_11538(s11538, c11538, in11538_1, in11538_2, c9541);
    wire[0:0] s11539, in11539_1, in11539_2;
    wire c11539;
    assign in11539_1 = {s9545[0]};
    assign in11539_2 = {s9546[0]};
    Full_Adder FA_11539(s11539, c11539, in11539_1, in11539_2, c9544);
    wire[0:0] s11540, in11540_1, in11540_2;
    wire c11540;
    assign in11540_1 = {s9548[0]};
    assign in11540_2 = {s9549[0]};
    Full_Adder FA_11540(s11540, c11540, in11540_1, in11540_2, s9547[0]);
    wire[0:0] s11541, in11541_1, in11541_2;
    wire c11541;
    assign in11541_1 = {s9551[0]};
    assign in11541_2 = {s9552[0]};
    Full_Adder FA_11541(s11541, c11541, in11541_1, in11541_2, s9550[0]);
    wire[0:0] s11542, in11542_1, in11542_2;
    wire c11542;
    assign in11542_1 = {s9554[0]};
    assign in11542_2 = {s9555[0]};
    Full_Adder FA_11542(s11542, c11542, in11542_1, in11542_2, s9553[0]);
    wire[0:0] s11543, in11543_1, in11543_2;
    wire c11543;
    assign in11543_1 = {c9546};
    assign in11543_2 = {c9547};
    Full_Adder FA_11543(s11543, c11543, in11543_1, in11543_2, c9545);
    wire[0:0] s11544, in11544_1, in11544_2;
    wire c11544;
    assign in11544_1 = {c9549};
    assign in11544_2 = {c9550};
    Full_Adder FA_11544(s11544, c11544, in11544_1, in11544_2, c9548);
    wire[0:0] s11545, in11545_1, in11545_2;
    wire c11545;
    assign in11545_1 = {c9552};
    assign in11545_2 = {c9553};
    Full_Adder FA_11545(s11545, c11545, in11545_1, in11545_2, c9551);
    wire[0:0] s11546, in11546_1, in11546_2;
    wire c11546;
    assign in11546_1 = {c9555};
    assign in11546_2 = {c9556};
    Full_Adder FA_11546(s11546, c11546, in11546_1, in11546_2, c9554);
    wire[0:0] s11547, in11547_1, in11547_2;
    wire c11547;
    assign in11547_1 = {s9558[0]};
    assign in11547_2 = {s9559[0]};
    Full_Adder FA_11547(s11547, c11547, in11547_1, in11547_2, c9557);
    wire[0:0] s11548, in11548_1, in11548_2;
    wire c11548;
    assign in11548_1 = {s9561[0]};
    assign in11548_2 = {s9562[0]};
    Full_Adder FA_11548(s11548, c11548, in11548_1, in11548_2, s9560[0]);
    wire[0:0] s11549, in11549_1, in11549_2;
    wire c11549;
    assign in11549_1 = {s9564[0]};
    assign in11549_2 = {s9565[0]};
    Full_Adder FA_11549(s11549, c11549, in11549_1, in11549_2, s9563[0]);
    wire[0:0] s11550, in11550_1, in11550_2;
    wire c11550;
    assign in11550_1 = {s9567[0]};
    assign in11550_2 = {s9568[0]};
    Full_Adder FA_11550(s11550, c11550, in11550_1, in11550_2, s9566[0]);
    wire[0:0] s11551, in11551_1, in11551_2;
    wire c11551;
    assign in11551_1 = {c9559};
    assign in11551_2 = {c9560};
    Full_Adder FA_11551(s11551, c11551, in11551_1, in11551_2, c9558);
    wire[0:0] s11552, in11552_1, in11552_2;
    wire c11552;
    assign in11552_1 = {c9562};
    assign in11552_2 = {c9563};
    Full_Adder FA_11552(s11552, c11552, in11552_1, in11552_2, c9561);
    wire[0:0] s11553, in11553_1, in11553_2;
    wire c11553;
    assign in11553_1 = {c9565};
    assign in11553_2 = {c9566};
    Full_Adder FA_11553(s11553, c11553, in11553_1, in11553_2, c9564);
    wire[0:0] s11554, in11554_1, in11554_2;
    wire c11554;
    assign in11554_1 = {c9568};
    assign in11554_2 = {c9569};
    Full_Adder FA_11554(s11554, c11554, in11554_1, in11554_2, c9567);
    wire[0:0] s11555, in11555_1, in11555_2;
    wire c11555;
    assign in11555_1 = {s9571[0]};
    assign in11555_2 = {s9572[0]};
    Full_Adder FA_11555(s11555, c11555, in11555_1, in11555_2, c9570);
    wire[0:0] s11556, in11556_1, in11556_2;
    wire c11556;
    assign in11556_1 = {s9574[0]};
    assign in11556_2 = {s9575[0]};
    Full_Adder FA_11556(s11556, c11556, in11556_1, in11556_2, s9573[0]);
    wire[0:0] s11557, in11557_1, in11557_2;
    wire c11557;
    assign in11557_1 = {s9577[0]};
    assign in11557_2 = {s9578[0]};
    Full_Adder FA_11557(s11557, c11557, in11557_1, in11557_2, s9576[0]);
    wire[0:0] s11558, in11558_1, in11558_2;
    wire c11558;
    assign in11558_1 = {s9580[0]};
    assign in11558_2 = {s9581[0]};
    Full_Adder FA_11558(s11558, c11558, in11558_1, in11558_2, s9579[0]);
    wire[0:0] s11559, in11559_1, in11559_2;
    wire c11559;
    assign in11559_1 = {c9572};
    assign in11559_2 = {c9573};
    Full_Adder FA_11559(s11559, c11559, in11559_1, in11559_2, c9571);
    wire[0:0] s11560, in11560_1, in11560_2;
    wire c11560;
    assign in11560_1 = {c9575};
    assign in11560_2 = {c9576};
    Full_Adder FA_11560(s11560, c11560, in11560_1, in11560_2, c9574);
    wire[0:0] s11561, in11561_1, in11561_2;
    wire c11561;
    assign in11561_1 = {c9578};
    assign in11561_2 = {c9579};
    Full_Adder FA_11561(s11561, c11561, in11561_1, in11561_2, c9577);
    wire[0:0] s11562, in11562_1, in11562_2;
    wire c11562;
    assign in11562_1 = {c9581};
    assign in11562_2 = {c9582};
    Full_Adder FA_11562(s11562, c11562, in11562_1, in11562_2, c9580);
    wire[0:0] s11563, in11563_1, in11563_2;
    wire c11563;
    assign in11563_1 = {s9584[0]};
    assign in11563_2 = {s9585[0]};
    Full_Adder FA_11563(s11563, c11563, in11563_1, in11563_2, c9583);
    wire[0:0] s11564, in11564_1, in11564_2;
    wire c11564;
    assign in11564_1 = {s9587[0]};
    assign in11564_2 = {s9588[0]};
    Full_Adder FA_11564(s11564, c11564, in11564_1, in11564_2, s9586[0]);
    wire[0:0] s11565, in11565_1, in11565_2;
    wire c11565;
    assign in11565_1 = {s9590[0]};
    assign in11565_2 = {s9591[0]};
    Full_Adder FA_11565(s11565, c11565, in11565_1, in11565_2, s9589[0]);
    wire[0:0] s11566, in11566_1, in11566_2;
    wire c11566;
    assign in11566_1 = {s9593[0]};
    assign in11566_2 = {s9594[0]};
    Full_Adder FA_11566(s11566, c11566, in11566_1, in11566_2, s9592[0]);
    wire[0:0] s11567, in11567_1, in11567_2;
    wire c11567;
    assign in11567_1 = {c9585};
    assign in11567_2 = {c9586};
    Full_Adder FA_11567(s11567, c11567, in11567_1, in11567_2, c9584);
    wire[0:0] s11568, in11568_1, in11568_2;
    wire c11568;
    assign in11568_1 = {c9588};
    assign in11568_2 = {c9589};
    Full_Adder FA_11568(s11568, c11568, in11568_1, in11568_2, c9587);
    wire[0:0] s11569, in11569_1, in11569_2;
    wire c11569;
    assign in11569_1 = {c9591};
    assign in11569_2 = {c9592};
    Full_Adder FA_11569(s11569, c11569, in11569_1, in11569_2, c9590);
    wire[0:0] s11570, in11570_1, in11570_2;
    wire c11570;
    assign in11570_1 = {c9594};
    assign in11570_2 = {c9595};
    Full_Adder FA_11570(s11570, c11570, in11570_1, in11570_2, c9593);
    wire[0:0] s11571, in11571_1, in11571_2;
    wire c11571;
    assign in11571_1 = {s9597[0]};
    assign in11571_2 = {s9598[0]};
    Full_Adder FA_11571(s11571, c11571, in11571_1, in11571_2, c9596);
    wire[0:0] s11572, in11572_1, in11572_2;
    wire c11572;
    assign in11572_1 = {s9600[0]};
    assign in11572_2 = {s9601[0]};
    Full_Adder FA_11572(s11572, c11572, in11572_1, in11572_2, s9599[0]);
    wire[0:0] s11573, in11573_1, in11573_2;
    wire c11573;
    assign in11573_1 = {s9603[0]};
    assign in11573_2 = {s9604[0]};
    Full_Adder FA_11573(s11573, c11573, in11573_1, in11573_2, s9602[0]);
    wire[0:0] s11574, in11574_1, in11574_2;
    wire c11574;
    assign in11574_1 = {s9606[0]};
    assign in11574_2 = {s9607[0]};
    Full_Adder FA_11574(s11574, c11574, in11574_1, in11574_2, s9605[0]);
    wire[0:0] s11575, in11575_1, in11575_2;
    wire c11575;
    assign in11575_1 = {c9598};
    assign in11575_2 = {c9599};
    Full_Adder FA_11575(s11575, c11575, in11575_1, in11575_2, c9597);
    wire[0:0] s11576, in11576_1, in11576_2;
    wire c11576;
    assign in11576_1 = {c9601};
    assign in11576_2 = {c9602};
    Full_Adder FA_11576(s11576, c11576, in11576_1, in11576_2, c9600);
    wire[0:0] s11577, in11577_1, in11577_2;
    wire c11577;
    assign in11577_1 = {c9604};
    assign in11577_2 = {c9605};
    Full_Adder FA_11577(s11577, c11577, in11577_1, in11577_2, c9603);
    wire[0:0] s11578, in11578_1, in11578_2;
    wire c11578;
    assign in11578_1 = {c9607};
    assign in11578_2 = {c9608};
    Full_Adder FA_11578(s11578, c11578, in11578_1, in11578_2, c9606);
    wire[0:0] s11579, in11579_1, in11579_2;
    wire c11579;
    assign in11579_1 = {s9610[0]};
    assign in11579_2 = {s9611[0]};
    Full_Adder FA_11579(s11579, c11579, in11579_1, in11579_2, c9609);
    wire[0:0] s11580, in11580_1, in11580_2;
    wire c11580;
    assign in11580_1 = {s9613[0]};
    assign in11580_2 = {s9614[0]};
    Full_Adder FA_11580(s11580, c11580, in11580_1, in11580_2, s9612[0]);
    wire[0:0] s11581, in11581_1, in11581_2;
    wire c11581;
    assign in11581_1 = {s9616[0]};
    assign in11581_2 = {s9617[0]};
    Full_Adder FA_11581(s11581, c11581, in11581_1, in11581_2, s9615[0]);
    wire[0:0] s11582, in11582_1, in11582_2;
    wire c11582;
    assign in11582_1 = {s9619[0]};
    assign in11582_2 = {s9620[0]};
    Full_Adder FA_11582(s11582, c11582, in11582_1, in11582_2, s9618[0]);
    wire[0:0] s11583, in11583_1, in11583_2;
    wire c11583;
    assign in11583_1 = {c9611};
    assign in11583_2 = {c9612};
    Full_Adder FA_11583(s11583, c11583, in11583_1, in11583_2, c9610);
    wire[0:0] s11584, in11584_1, in11584_2;
    wire c11584;
    assign in11584_1 = {c9614};
    assign in11584_2 = {c9615};
    Full_Adder FA_11584(s11584, c11584, in11584_1, in11584_2, c9613);
    wire[0:0] s11585, in11585_1, in11585_2;
    wire c11585;
    assign in11585_1 = {c9617};
    assign in11585_2 = {c9618};
    Full_Adder FA_11585(s11585, c11585, in11585_1, in11585_2, c9616);
    wire[0:0] s11586, in11586_1, in11586_2;
    wire c11586;
    assign in11586_1 = {c9620};
    assign in11586_2 = {c9621};
    Full_Adder FA_11586(s11586, c11586, in11586_1, in11586_2, c9619);
    wire[0:0] s11587, in11587_1, in11587_2;
    wire c11587;
    assign in11587_1 = {s9623[0]};
    assign in11587_2 = {s9624[0]};
    Full_Adder FA_11587(s11587, c11587, in11587_1, in11587_2, c9622);
    wire[0:0] s11588, in11588_1, in11588_2;
    wire c11588;
    assign in11588_1 = {s9626[0]};
    assign in11588_2 = {s9627[0]};
    Full_Adder FA_11588(s11588, c11588, in11588_1, in11588_2, s9625[0]);
    wire[0:0] s11589, in11589_1, in11589_2;
    wire c11589;
    assign in11589_1 = {s9629[0]};
    assign in11589_2 = {s9630[0]};
    Full_Adder FA_11589(s11589, c11589, in11589_1, in11589_2, s9628[0]);
    wire[0:0] s11590, in11590_1, in11590_2;
    wire c11590;
    assign in11590_1 = {s9632[0]};
    assign in11590_2 = {s9633[0]};
    Full_Adder FA_11590(s11590, c11590, in11590_1, in11590_2, s9631[0]);
    wire[0:0] s11591, in11591_1, in11591_2;
    wire c11591;
    assign in11591_1 = {c9624};
    assign in11591_2 = {c9625};
    Full_Adder FA_11591(s11591, c11591, in11591_1, in11591_2, c9623);
    wire[0:0] s11592, in11592_1, in11592_2;
    wire c11592;
    assign in11592_1 = {c9627};
    assign in11592_2 = {c9628};
    Full_Adder FA_11592(s11592, c11592, in11592_1, in11592_2, c9626);
    wire[0:0] s11593, in11593_1, in11593_2;
    wire c11593;
    assign in11593_1 = {c9630};
    assign in11593_2 = {c9631};
    Full_Adder FA_11593(s11593, c11593, in11593_1, in11593_2, c9629);
    wire[0:0] s11594, in11594_1, in11594_2;
    wire c11594;
    assign in11594_1 = {c9633};
    assign in11594_2 = {c9634};
    Full_Adder FA_11594(s11594, c11594, in11594_1, in11594_2, c9632);
    wire[0:0] s11595, in11595_1, in11595_2;
    wire c11595;
    assign in11595_1 = {s9636[0]};
    assign in11595_2 = {s9637[0]};
    Full_Adder FA_11595(s11595, c11595, in11595_1, in11595_2, c9635);
    wire[0:0] s11596, in11596_1, in11596_2;
    wire c11596;
    assign in11596_1 = {s9639[0]};
    assign in11596_2 = {s9640[0]};
    Full_Adder FA_11596(s11596, c11596, in11596_1, in11596_2, s9638[0]);
    wire[0:0] s11597, in11597_1, in11597_2;
    wire c11597;
    assign in11597_1 = {s9642[0]};
    assign in11597_2 = {s9643[0]};
    Full_Adder FA_11597(s11597, c11597, in11597_1, in11597_2, s9641[0]);
    wire[0:0] s11598, in11598_1, in11598_2;
    wire c11598;
    assign in11598_1 = {s9645[0]};
    assign in11598_2 = {s9646[0]};
    Full_Adder FA_11598(s11598, c11598, in11598_1, in11598_2, s9644[0]);
    wire[0:0] s11599, in11599_1, in11599_2;
    wire c11599;
    assign in11599_1 = {c9637};
    assign in11599_2 = {c9638};
    Full_Adder FA_11599(s11599, c11599, in11599_1, in11599_2, c9636);
    wire[0:0] s11600, in11600_1, in11600_2;
    wire c11600;
    assign in11600_1 = {c9640};
    assign in11600_2 = {c9641};
    Full_Adder FA_11600(s11600, c11600, in11600_1, in11600_2, c9639);
    wire[0:0] s11601, in11601_1, in11601_2;
    wire c11601;
    assign in11601_1 = {c9643};
    assign in11601_2 = {c9644};
    Full_Adder FA_11601(s11601, c11601, in11601_1, in11601_2, c9642);
    wire[0:0] s11602, in11602_1, in11602_2;
    wire c11602;
    assign in11602_1 = {c9646};
    assign in11602_2 = {c9647};
    Full_Adder FA_11602(s11602, c11602, in11602_1, in11602_2, c9645);
    wire[0:0] s11603, in11603_1, in11603_2;
    wire c11603;
    assign in11603_1 = {s9649[0]};
    assign in11603_2 = {s9650[0]};
    Full_Adder FA_11603(s11603, c11603, in11603_1, in11603_2, c9648);
    wire[0:0] s11604, in11604_1, in11604_2;
    wire c11604;
    assign in11604_1 = {s9652[0]};
    assign in11604_2 = {s9653[0]};
    Full_Adder FA_11604(s11604, c11604, in11604_1, in11604_2, s9651[0]);
    wire[0:0] s11605, in11605_1, in11605_2;
    wire c11605;
    assign in11605_1 = {s9655[0]};
    assign in11605_2 = {s9656[0]};
    Full_Adder FA_11605(s11605, c11605, in11605_1, in11605_2, s9654[0]);
    wire[0:0] s11606, in11606_1, in11606_2;
    wire c11606;
    assign in11606_1 = {s9658[0]};
    assign in11606_2 = {s9659[0]};
    Full_Adder FA_11606(s11606, c11606, in11606_1, in11606_2, s9657[0]);
    wire[0:0] s11607, in11607_1, in11607_2;
    wire c11607;
    assign in11607_1 = {c9650};
    assign in11607_2 = {c9651};
    Full_Adder FA_11607(s11607, c11607, in11607_1, in11607_2, c9649);
    wire[0:0] s11608, in11608_1, in11608_2;
    wire c11608;
    assign in11608_1 = {c9653};
    assign in11608_2 = {c9654};
    Full_Adder FA_11608(s11608, c11608, in11608_1, in11608_2, c9652);
    wire[0:0] s11609, in11609_1, in11609_2;
    wire c11609;
    assign in11609_1 = {c9656};
    assign in11609_2 = {c9657};
    Full_Adder FA_11609(s11609, c11609, in11609_1, in11609_2, c9655);
    wire[0:0] s11610, in11610_1, in11610_2;
    wire c11610;
    assign in11610_1 = {c9659};
    assign in11610_2 = {c9660};
    Full_Adder FA_11610(s11610, c11610, in11610_1, in11610_2, c9658);
    wire[0:0] s11611, in11611_1, in11611_2;
    wire c11611;
    assign in11611_1 = {s9662[0]};
    assign in11611_2 = {s9663[0]};
    Full_Adder FA_11611(s11611, c11611, in11611_1, in11611_2, c9661);
    wire[0:0] s11612, in11612_1, in11612_2;
    wire c11612;
    assign in11612_1 = {s9665[0]};
    assign in11612_2 = {s9666[0]};
    Full_Adder FA_11612(s11612, c11612, in11612_1, in11612_2, s9664[0]);
    wire[0:0] s11613, in11613_1, in11613_2;
    wire c11613;
    assign in11613_1 = {s9668[0]};
    assign in11613_2 = {s9669[0]};
    Full_Adder FA_11613(s11613, c11613, in11613_1, in11613_2, s9667[0]);
    wire[0:0] s11614, in11614_1, in11614_2;
    wire c11614;
    assign in11614_1 = {s9671[0]};
    assign in11614_2 = {s9672[0]};
    Full_Adder FA_11614(s11614, c11614, in11614_1, in11614_2, s9670[0]);
    wire[0:0] s11615, in11615_1, in11615_2;
    wire c11615;
    assign in11615_1 = {c9663};
    assign in11615_2 = {c9664};
    Full_Adder FA_11615(s11615, c11615, in11615_1, in11615_2, c9662);
    wire[0:0] s11616, in11616_1, in11616_2;
    wire c11616;
    assign in11616_1 = {c9666};
    assign in11616_2 = {c9667};
    Full_Adder FA_11616(s11616, c11616, in11616_1, in11616_2, c9665);
    wire[0:0] s11617, in11617_1, in11617_2;
    wire c11617;
    assign in11617_1 = {c9669};
    assign in11617_2 = {c9670};
    Full_Adder FA_11617(s11617, c11617, in11617_1, in11617_2, c9668);
    wire[0:0] s11618, in11618_1, in11618_2;
    wire c11618;
    assign in11618_1 = {c9672};
    assign in11618_2 = {c9673};
    Full_Adder FA_11618(s11618, c11618, in11618_1, in11618_2, c9671);
    wire[0:0] s11619, in11619_1, in11619_2;
    wire c11619;
    assign in11619_1 = {s9675[0]};
    assign in11619_2 = {s9676[0]};
    Full_Adder FA_11619(s11619, c11619, in11619_1, in11619_2, c9674);
    wire[0:0] s11620, in11620_1, in11620_2;
    wire c11620;
    assign in11620_1 = {s9678[0]};
    assign in11620_2 = {s9679[0]};
    Full_Adder FA_11620(s11620, c11620, in11620_1, in11620_2, s9677[0]);
    wire[0:0] s11621, in11621_1, in11621_2;
    wire c11621;
    assign in11621_1 = {s9681[0]};
    assign in11621_2 = {s9682[0]};
    Full_Adder FA_11621(s11621, c11621, in11621_1, in11621_2, s9680[0]);
    wire[0:0] s11622, in11622_1, in11622_2;
    wire c11622;
    assign in11622_1 = {s9684[0]};
    assign in11622_2 = {s9685[0]};
    Full_Adder FA_11622(s11622, c11622, in11622_1, in11622_2, s9683[0]);
    wire[0:0] s11623, in11623_1, in11623_2;
    wire c11623;
    assign in11623_1 = {c9676};
    assign in11623_2 = {c9677};
    Full_Adder FA_11623(s11623, c11623, in11623_1, in11623_2, c9675);
    wire[0:0] s11624, in11624_1, in11624_2;
    wire c11624;
    assign in11624_1 = {c9679};
    assign in11624_2 = {c9680};
    Full_Adder FA_11624(s11624, c11624, in11624_1, in11624_2, c9678);
    wire[0:0] s11625, in11625_1, in11625_2;
    wire c11625;
    assign in11625_1 = {c9682};
    assign in11625_2 = {c9683};
    Full_Adder FA_11625(s11625, c11625, in11625_1, in11625_2, c9681);
    wire[0:0] s11626, in11626_1, in11626_2;
    wire c11626;
    assign in11626_1 = {c9685};
    assign in11626_2 = {c9686};
    Full_Adder FA_11626(s11626, c11626, in11626_1, in11626_2, c9684);
    wire[0:0] s11627, in11627_1, in11627_2;
    wire c11627;
    assign in11627_1 = {s9688[0]};
    assign in11627_2 = {s9689[0]};
    Full_Adder FA_11627(s11627, c11627, in11627_1, in11627_2, c9687);
    wire[0:0] s11628, in11628_1, in11628_2;
    wire c11628;
    assign in11628_1 = {s9691[0]};
    assign in11628_2 = {s9692[0]};
    Full_Adder FA_11628(s11628, c11628, in11628_1, in11628_2, s9690[0]);
    wire[0:0] s11629, in11629_1, in11629_2;
    wire c11629;
    assign in11629_1 = {s9694[0]};
    assign in11629_2 = {s9695[0]};
    Full_Adder FA_11629(s11629, c11629, in11629_1, in11629_2, s9693[0]);
    wire[0:0] s11630, in11630_1, in11630_2;
    wire c11630;
    assign in11630_1 = {s9697[0]};
    assign in11630_2 = {s9698[0]};
    Full_Adder FA_11630(s11630, c11630, in11630_1, in11630_2, s9696[0]);
    wire[0:0] s11631, in11631_1, in11631_2;
    wire c11631;
    assign in11631_1 = {c9689};
    assign in11631_2 = {c9690};
    Full_Adder FA_11631(s11631, c11631, in11631_1, in11631_2, c9688);
    wire[0:0] s11632, in11632_1, in11632_2;
    wire c11632;
    assign in11632_1 = {c9692};
    assign in11632_2 = {c9693};
    Full_Adder FA_11632(s11632, c11632, in11632_1, in11632_2, c9691);
    wire[0:0] s11633, in11633_1, in11633_2;
    wire c11633;
    assign in11633_1 = {c9695};
    assign in11633_2 = {c9696};
    Full_Adder FA_11633(s11633, c11633, in11633_1, in11633_2, c9694);
    wire[0:0] s11634, in11634_1, in11634_2;
    wire c11634;
    assign in11634_1 = {c9698};
    assign in11634_2 = {c9699};
    Full_Adder FA_11634(s11634, c11634, in11634_1, in11634_2, c9697);
    wire[0:0] s11635, in11635_1, in11635_2;
    wire c11635;
    assign in11635_1 = {s9701[0]};
    assign in11635_2 = {s9702[0]};
    Full_Adder FA_11635(s11635, c11635, in11635_1, in11635_2, c9700);
    wire[0:0] s11636, in11636_1, in11636_2;
    wire c11636;
    assign in11636_1 = {s9704[0]};
    assign in11636_2 = {s9705[0]};
    Full_Adder FA_11636(s11636, c11636, in11636_1, in11636_2, s9703[0]);
    wire[0:0] s11637, in11637_1, in11637_2;
    wire c11637;
    assign in11637_1 = {s9707[0]};
    assign in11637_2 = {s9708[0]};
    Full_Adder FA_11637(s11637, c11637, in11637_1, in11637_2, s9706[0]);
    wire[0:0] s11638, in11638_1, in11638_2;
    wire c11638;
    assign in11638_1 = {s9710[0]};
    assign in11638_2 = {s9711[0]};
    Full_Adder FA_11638(s11638, c11638, in11638_1, in11638_2, s9709[0]);
    wire[0:0] s11639, in11639_1, in11639_2;
    wire c11639;
    assign in11639_1 = {c9702};
    assign in11639_2 = {c9703};
    Full_Adder FA_11639(s11639, c11639, in11639_1, in11639_2, c9701);
    wire[0:0] s11640, in11640_1, in11640_2;
    wire c11640;
    assign in11640_1 = {c9705};
    assign in11640_2 = {c9706};
    Full_Adder FA_11640(s11640, c11640, in11640_1, in11640_2, c9704);
    wire[0:0] s11641, in11641_1, in11641_2;
    wire c11641;
    assign in11641_1 = {c9708};
    assign in11641_2 = {c9709};
    Full_Adder FA_11641(s11641, c11641, in11641_1, in11641_2, c9707);
    wire[0:0] s11642, in11642_1, in11642_2;
    wire c11642;
    assign in11642_1 = {c9711};
    assign in11642_2 = {c9712};
    Full_Adder FA_11642(s11642, c11642, in11642_1, in11642_2, c9710);
    wire[0:0] s11643, in11643_1, in11643_2;
    wire c11643;
    assign in11643_1 = {s9714[0]};
    assign in11643_2 = {s9715[0]};
    Full_Adder FA_11643(s11643, c11643, in11643_1, in11643_2, c9713);
    wire[0:0] s11644, in11644_1, in11644_2;
    wire c11644;
    assign in11644_1 = {s9717[0]};
    assign in11644_2 = {s9718[0]};
    Full_Adder FA_11644(s11644, c11644, in11644_1, in11644_2, s9716[0]);
    wire[0:0] s11645, in11645_1, in11645_2;
    wire c11645;
    assign in11645_1 = {s9720[0]};
    assign in11645_2 = {s9721[0]};
    Full_Adder FA_11645(s11645, c11645, in11645_1, in11645_2, s9719[0]);
    wire[0:0] s11646, in11646_1, in11646_2;
    wire c11646;
    assign in11646_1 = {s9723[0]};
    assign in11646_2 = {s9724[0]};
    Full_Adder FA_11646(s11646, c11646, in11646_1, in11646_2, s9722[0]);
    wire[0:0] s11647, in11647_1, in11647_2;
    wire c11647;
    assign in11647_1 = {c9715};
    assign in11647_2 = {c9716};
    Full_Adder FA_11647(s11647, c11647, in11647_1, in11647_2, c9714);
    wire[0:0] s11648, in11648_1, in11648_2;
    wire c11648;
    assign in11648_1 = {c9718};
    assign in11648_2 = {c9719};
    Full_Adder FA_11648(s11648, c11648, in11648_1, in11648_2, c9717);
    wire[0:0] s11649, in11649_1, in11649_2;
    wire c11649;
    assign in11649_1 = {c9721};
    assign in11649_2 = {c9722};
    Full_Adder FA_11649(s11649, c11649, in11649_1, in11649_2, c9720);
    wire[0:0] s11650, in11650_1, in11650_2;
    wire c11650;
    assign in11650_1 = {c9724};
    assign in11650_2 = {c9725};
    Full_Adder FA_11650(s11650, c11650, in11650_1, in11650_2, c9723);
    wire[0:0] s11651, in11651_1, in11651_2;
    wire c11651;
    assign in11651_1 = {s9727[0]};
    assign in11651_2 = {s9728[0]};
    Full_Adder FA_11651(s11651, c11651, in11651_1, in11651_2, c9726);
    wire[0:0] s11652, in11652_1, in11652_2;
    wire c11652;
    assign in11652_1 = {s9730[0]};
    assign in11652_2 = {s9731[0]};
    Full_Adder FA_11652(s11652, c11652, in11652_1, in11652_2, s9729[0]);
    wire[0:0] s11653, in11653_1, in11653_2;
    wire c11653;
    assign in11653_1 = {s9733[0]};
    assign in11653_2 = {s9734[0]};
    Full_Adder FA_11653(s11653, c11653, in11653_1, in11653_2, s9732[0]);
    wire[0:0] s11654, in11654_1, in11654_2;
    wire c11654;
    assign in11654_1 = {s9736[0]};
    assign in11654_2 = {s9737[0]};
    Full_Adder FA_11654(s11654, c11654, in11654_1, in11654_2, s9735[0]);
    wire[0:0] s11655, in11655_1, in11655_2;
    wire c11655;
    assign in11655_1 = {c9728};
    assign in11655_2 = {c9729};
    Full_Adder FA_11655(s11655, c11655, in11655_1, in11655_2, c9727);
    wire[0:0] s11656, in11656_1, in11656_2;
    wire c11656;
    assign in11656_1 = {c9731};
    assign in11656_2 = {c9732};
    Full_Adder FA_11656(s11656, c11656, in11656_1, in11656_2, c9730);
    wire[0:0] s11657, in11657_1, in11657_2;
    wire c11657;
    assign in11657_1 = {c9734};
    assign in11657_2 = {c9735};
    Full_Adder FA_11657(s11657, c11657, in11657_1, in11657_2, c9733);
    wire[0:0] s11658, in11658_1, in11658_2;
    wire c11658;
    assign in11658_1 = {c9737};
    assign in11658_2 = {c9738};
    Full_Adder FA_11658(s11658, c11658, in11658_1, in11658_2, c9736);
    wire[0:0] s11659, in11659_1, in11659_2;
    wire c11659;
    assign in11659_1 = {s9740[0]};
    assign in11659_2 = {s9741[0]};
    Full_Adder FA_11659(s11659, c11659, in11659_1, in11659_2, c9739);
    wire[0:0] s11660, in11660_1, in11660_2;
    wire c11660;
    assign in11660_1 = {s9743[0]};
    assign in11660_2 = {s9744[0]};
    Full_Adder FA_11660(s11660, c11660, in11660_1, in11660_2, s9742[0]);
    wire[0:0] s11661, in11661_1, in11661_2;
    wire c11661;
    assign in11661_1 = {s9746[0]};
    assign in11661_2 = {s9747[0]};
    Full_Adder FA_11661(s11661, c11661, in11661_1, in11661_2, s9745[0]);
    wire[0:0] s11662, in11662_1, in11662_2;
    wire c11662;
    assign in11662_1 = {s9749[0]};
    assign in11662_2 = {s9750[0]};
    Full_Adder FA_11662(s11662, c11662, in11662_1, in11662_2, s9748[0]);
    wire[0:0] s11663, in11663_1, in11663_2;
    wire c11663;
    assign in11663_1 = {c9741};
    assign in11663_2 = {c9742};
    Full_Adder FA_11663(s11663, c11663, in11663_1, in11663_2, c9740);
    wire[0:0] s11664, in11664_1, in11664_2;
    wire c11664;
    assign in11664_1 = {c9744};
    assign in11664_2 = {c9745};
    Full_Adder FA_11664(s11664, c11664, in11664_1, in11664_2, c9743);
    wire[0:0] s11665, in11665_1, in11665_2;
    wire c11665;
    assign in11665_1 = {c9747};
    assign in11665_2 = {c9748};
    Full_Adder FA_11665(s11665, c11665, in11665_1, in11665_2, c9746);
    wire[0:0] s11666, in11666_1, in11666_2;
    wire c11666;
    assign in11666_1 = {c9750};
    assign in11666_2 = {c9751};
    Full_Adder FA_11666(s11666, c11666, in11666_1, in11666_2, c9749);
    wire[0:0] s11667, in11667_1, in11667_2;
    wire c11667;
    assign in11667_1 = {s9753[0]};
    assign in11667_2 = {s9754[0]};
    Full_Adder FA_11667(s11667, c11667, in11667_1, in11667_2, c9752);
    wire[0:0] s11668, in11668_1, in11668_2;
    wire c11668;
    assign in11668_1 = {s9756[0]};
    assign in11668_2 = {s9757[0]};
    Full_Adder FA_11668(s11668, c11668, in11668_1, in11668_2, s9755[0]);
    wire[0:0] s11669, in11669_1, in11669_2;
    wire c11669;
    assign in11669_1 = {s9759[0]};
    assign in11669_2 = {s9760[0]};
    Full_Adder FA_11669(s11669, c11669, in11669_1, in11669_2, s9758[0]);
    wire[0:0] s11670, in11670_1, in11670_2;
    wire c11670;
    assign in11670_1 = {s9762[0]};
    assign in11670_2 = {s9763[0]};
    Full_Adder FA_11670(s11670, c11670, in11670_1, in11670_2, s9761[0]);
    wire[0:0] s11671, in11671_1, in11671_2;
    wire c11671;
    assign in11671_1 = {c9754};
    assign in11671_2 = {c9755};
    Full_Adder FA_11671(s11671, c11671, in11671_1, in11671_2, c9753);
    wire[0:0] s11672, in11672_1, in11672_2;
    wire c11672;
    assign in11672_1 = {c9757};
    assign in11672_2 = {c9758};
    Full_Adder FA_11672(s11672, c11672, in11672_1, in11672_2, c9756);
    wire[0:0] s11673, in11673_1, in11673_2;
    wire c11673;
    assign in11673_1 = {c9760};
    assign in11673_2 = {c9761};
    Full_Adder FA_11673(s11673, c11673, in11673_1, in11673_2, c9759);
    wire[0:0] s11674, in11674_1, in11674_2;
    wire c11674;
    assign in11674_1 = {c9763};
    assign in11674_2 = {c9764};
    Full_Adder FA_11674(s11674, c11674, in11674_1, in11674_2, c9762);
    wire[0:0] s11675, in11675_1, in11675_2;
    wire c11675;
    assign in11675_1 = {s9766[0]};
    assign in11675_2 = {s9767[0]};
    Full_Adder FA_11675(s11675, c11675, in11675_1, in11675_2, c9765);
    wire[0:0] s11676, in11676_1, in11676_2;
    wire c11676;
    assign in11676_1 = {s9769[0]};
    assign in11676_2 = {s9770[0]};
    Full_Adder FA_11676(s11676, c11676, in11676_1, in11676_2, s9768[0]);
    wire[0:0] s11677, in11677_1, in11677_2;
    wire c11677;
    assign in11677_1 = {s9772[0]};
    assign in11677_2 = {s9773[0]};
    Full_Adder FA_11677(s11677, c11677, in11677_1, in11677_2, s9771[0]);
    wire[0:0] s11678, in11678_1, in11678_2;
    wire c11678;
    assign in11678_1 = {s9775[0]};
    assign in11678_2 = {s9776[0]};
    Full_Adder FA_11678(s11678, c11678, in11678_1, in11678_2, s9774[0]);
    wire[0:0] s11679, in11679_1, in11679_2;
    wire c11679;
    assign in11679_1 = {c9767};
    assign in11679_2 = {c9768};
    Full_Adder FA_11679(s11679, c11679, in11679_1, in11679_2, c9766);
    wire[0:0] s11680, in11680_1, in11680_2;
    wire c11680;
    assign in11680_1 = {c9770};
    assign in11680_2 = {c9771};
    Full_Adder FA_11680(s11680, c11680, in11680_1, in11680_2, c9769);
    wire[0:0] s11681, in11681_1, in11681_2;
    wire c11681;
    assign in11681_1 = {c9773};
    assign in11681_2 = {c9774};
    Full_Adder FA_11681(s11681, c11681, in11681_1, in11681_2, c9772);
    wire[0:0] s11682, in11682_1, in11682_2;
    wire c11682;
    assign in11682_1 = {c9776};
    assign in11682_2 = {c9777};
    Full_Adder FA_11682(s11682, c11682, in11682_1, in11682_2, c9775);
    wire[0:0] s11683, in11683_1, in11683_2;
    wire c11683;
    assign in11683_1 = {s9779[0]};
    assign in11683_2 = {s9780[0]};
    Full_Adder FA_11683(s11683, c11683, in11683_1, in11683_2, c9778);
    wire[0:0] s11684, in11684_1, in11684_2;
    wire c11684;
    assign in11684_1 = {s9782[0]};
    assign in11684_2 = {s9783[0]};
    Full_Adder FA_11684(s11684, c11684, in11684_1, in11684_2, s9781[0]);
    wire[0:0] s11685, in11685_1, in11685_2;
    wire c11685;
    assign in11685_1 = {s9785[0]};
    assign in11685_2 = {s9786[0]};
    Full_Adder FA_11685(s11685, c11685, in11685_1, in11685_2, s9784[0]);
    wire[0:0] s11686, in11686_1, in11686_2;
    wire c11686;
    assign in11686_1 = {s9788[0]};
    assign in11686_2 = {s9789[0]};
    Full_Adder FA_11686(s11686, c11686, in11686_1, in11686_2, s9787[0]);
    wire[0:0] s11687, in11687_1, in11687_2;
    wire c11687;
    assign in11687_1 = {c9780};
    assign in11687_2 = {c9781};
    Full_Adder FA_11687(s11687, c11687, in11687_1, in11687_2, c9779);
    wire[0:0] s11688, in11688_1, in11688_2;
    wire c11688;
    assign in11688_1 = {c9783};
    assign in11688_2 = {c9784};
    Full_Adder FA_11688(s11688, c11688, in11688_1, in11688_2, c9782);
    wire[0:0] s11689, in11689_1, in11689_2;
    wire c11689;
    assign in11689_1 = {c9786};
    assign in11689_2 = {c9787};
    Full_Adder FA_11689(s11689, c11689, in11689_1, in11689_2, c9785);
    wire[0:0] s11690, in11690_1, in11690_2;
    wire c11690;
    assign in11690_1 = {c9789};
    assign in11690_2 = {c9790};
    Full_Adder FA_11690(s11690, c11690, in11690_1, in11690_2, c9788);
    wire[0:0] s11691, in11691_1, in11691_2;
    wire c11691;
    assign in11691_1 = {s9792[0]};
    assign in11691_2 = {s9793[0]};
    Full_Adder FA_11691(s11691, c11691, in11691_1, in11691_2, c9791);
    wire[0:0] s11692, in11692_1, in11692_2;
    wire c11692;
    assign in11692_1 = {s9795[0]};
    assign in11692_2 = {s9796[0]};
    Full_Adder FA_11692(s11692, c11692, in11692_1, in11692_2, s9794[0]);
    wire[0:0] s11693, in11693_1, in11693_2;
    wire c11693;
    assign in11693_1 = {s9798[0]};
    assign in11693_2 = {s9799[0]};
    Full_Adder FA_11693(s11693, c11693, in11693_1, in11693_2, s9797[0]);
    wire[0:0] s11694, in11694_1, in11694_2;
    wire c11694;
    assign in11694_1 = {s9801[0]};
    assign in11694_2 = {s9802[0]};
    Full_Adder FA_11694(s11694, c11694, in11694_1, in11694_2, s9800[0]);
    wire[0:0] s11695, in11695_1, in11695_2;
    wire c11695;
    assign in11695_1 = {c9793};
    assign in11695_2 = {c9794};
    Full_Adder FA_11695(s11695, c11695, in11695_1, in11695_2, c9792);
    wire[0:0] s11696, in11696_1, in11696_2;
    wire c11696;
    assign in11696_1 = {c9796};
    assign in11696_2 = {c9797};
    Full_Adder FA_11696(s11696, c11696, in11696_1, in11696_2, c9795);
    wire[0:0] s11697, in11697_1, in11697_2;
    wire c11697;
    assign in11697_1 = {c9799};
    assign in11697_2 = {c9800};
    Full_Adder FA_11697(s11697, c11697, in11697_1, in11697_2, c9798);
    wire[0:0] s11698, in11698_1, in11698_2;
    wire c11698;
    assign in11698_1 = {c9802};
    assign in11698_2 = {c9803};
    Full_Adder FA_11698(s11698, c11698, in11698_1, in11698_2, c9801);
    wire[0:0] s11699, in11699_1, in11699_2;
    wire c11699;
    assign in11699_1 = {s9805[0]};
    assign in11699_2 = {s9806[0]};
    Full_Adder FA_11699(s11699, c11699, in11699_1, in11699_2, c9804);
    wire[0:0] s11700, in11700_1, in11700_2;
    wire c11700;
    assign in11700_1 = {s9808[0]};
    assign in11700_2 = {s9809[0]};
    Full_Adder FA_11700(s11700, c11700, in11700_1, in11700_2, s9807[0]);
    wire[0:0] s11701, in11701_1, in11701_2;
    wire c11701;
    assign in11701_1 = {s9811[0]};
    assign in11701_2 = {s9812[0]};
    Full_Adder FA_11701(s11701, c11701, in11701_1, in11701_2, s9810[0]);
    wire[0:0] s11702, in11702_1, in11702_2;
    wire c11702;
    assign in11702_1 = {s9814[0]};
    assign in11702_2 = {s9815[0]};
    Full_Adder FA_11702(s11702, c11702, in11702_1, in11702_2, s9813[0]);
    wire[0:0] s11703, in11703_1, in11703_2;
    wire c11703;
    assign in11703_1 = {c9806};
    assign in11703_2 = {c9807};
    Full_Adder FA_11703(s11703, c11703, in11703_1, in11703_2, c9805);
    wire[0:0] s11704, in11704_1, in11704_2;
    wire c11704;
    assign in11704_1 = {c9809};
    assign in11704_2 = {c9810};
    Full_Adder FA_11704(s11704, c11704, in11704_1, in11704_2, c9808);
    wire[0:0] s11705, in11705_1, in11705_2;
    wire c11705;
    assign in11705_1 = {c9812};
    assign in11705_2 = {c9813};
    Full_Adder FA_11705(s11705, c11705, in11705_1, in11705_2, c9811);
    wire[0:0] s11706, in11706_1, in11706_2;
    wire c11706;
    assign in11706_1 = {c9815};
    assign in11706_2 = {c9816};
    Full_Adder FA_11706(s11706, c11706, in11706_1, in11706_2, c9814);
    wire[0:0] s11707, in11707_1, in11707_2;
    wire c11707;
    assign in11707_1 = {s9818[0]};
    assign in11707_2 = {s9819[0]};
    Full_Adder FA_11707(s11707, c11707, in11707_1, in11707_2, c9817);
    wire[0:0] s11708, in11708_1, in11708_2;
    wire c11708;
    assign in11708_1 = {s9821[0]};
    assign in11708_2 = {s9822[0]};
    Full_Adder FA_11708(s11708, c11708, in11708_1, in11708_2, s9820[0]);
    wire[0:0] s11709, in11709_1, in11709_2;
    wire c11709;
    assign in11709_1 = {s9824[0]};
    assign in11709_2 = {s9825[0]};
    Full_Adder FA_11709(s11709, c11709, in11709_1, in11709_2, s9823[0]);
    wire[0:0] s11710, in11710_1, in11710_2;
    wire c11710;
    assign in11710_1 = {s9827[0]};
    assign in11710_2 = {s9828[0]};
    Full_Adder FA_11710(s11710, c11710, in11710_1, in11710_2, s9826[0]);
    wire[0:0] s11711, in11711_1, in11711_2;
    wire c11711;
    assign in11711_1 = {c9819};
    assign in11711_2 = {c9820};
    Full_Adder FA_11711(s11711, c11711, in11711_1, in11711_2, c9818);
    wire[0:0] s11712, in11712_1, in11712_2;
    wire c11712;
    assign in11712_1 = {c9822};
    assign in11712_2 = {c9823};
    Full_Adder FA_11712(s11712, c11712, in11712_1, in11712_2, c9821);
    wire[0:0] s11713, in11713_1, in11713_2;
    wire c11713;
    assign in11713_1 = {c9825};
    assign in11713_2 = {c9826};
    Full_Adder FA_11713(s11713, c11713, in11713_1, in11713_2, c9824);
    wire[0:0] s11714, in11714_1, in11714_2;
    wire c11714;
    assign in11714_1 = {c9828};
    assign in11714_2 = {c9829};
    Full_Adder FA_11714(s11714, c11714, in11714_1, in11714_2, c9827);
    wire[0:0] s11715, in11715_1, in11715_2;
    wire c11715;
    assign in11715_1 = {s9831[0]};
    assign in11715_2 = {s9832[0]};
    Full_Adder FA_11715(s11715, c11715, in11715_1, in11715_2, c9830);
    wire[0:0] s11716, in11716_1, in11716_2;
    wire c11716;
    assign in11716_1 = {s9834[0]};
    assign in11716_2 = {s9835[0]};
    Full_Adder FA_11716(s11716, c11716, in11716_1, in11716_2, s9833[0]);
    wire[0:0] s11717, in11717_1, in11717_2;
    wire c11717;
    assign in11717_1 = {s9837[0]};
    assign in11717_2 = {s9838[0]};
    Full_Adder FA_11717(s11717, c11717, in11717_1, in11717_2, s9836[0]);
    wire[0:0] s11718, in11718_1, in11718_2;
    wire c11718;
    assign in11718_1 = {s9840[0]};
    assign in11718_2 = {s9841[0]};
    Full_Adder FA_11718(s11718, c11718, in11718_1, in11718_2, s9839[0]);
    wire[0:0] s11719, in11719_1, in11719_2;
    wire c11719;
    assign in11719_1 = {c9832};
    assign in11719_2 = {c9833};
    Full_Adder FA_11719(s11719, c11719, in11719_1, in11719_2, c9831);
    wire[0:0] s11720, in11720_1, in11720_2;
    wire c11720;
    assign in11720_1 = {c9835};
    assign in11720_2 = {c9836};
    Full_Adder FA_11720(s11720, c11720, in11720_1, in11720_2, c9834);
    wire[0:0] s11721, in11721_1, in11721_2;
    wire c11721;
    assign in11721_1 = {c9838};
    assign in11721_2 = {c9839};
    Full_Adder FA_11721(s11721, c11721, in11721_1, in11721_2, c9837);
    wire[0:0] s11722, in11722_1, in11722_2;
    wire c11722;
    assign in11722_1 = {c9841};
    assign in11722_2 = {c9842};
    Full_Adder FA_11722(s11722, c11722, in11722_1, in11722_2, c9840);
    wire[0:0] s11723, in11723_1, in11723_2;
    wire c11723;
    assign in11723_1 = {s9844[0]};
    assign in11723_2 = {s9845[0]};
    Full_Adder FA_11723(s11723, c11723, in11723_1, in11723_2, c9843);
    wire[0:0] s11724, in11724_1, in11724_2;
    wire c11724;
    assign in11724_1 = {s9847[0]};
    assign in11724_2 = {s9848[0]};
    Full_Adder FA_11724(s11724, c11724, in11724_1, in11724_2, s9846[0]);
    wire[0:0] s11725, in11725_1, in11725_2;
    wire c11725;
    assign in11725_1 = {s9850[0]};
    assign in11725_2 = {s9851[0]};
    Full_Adder FA_11725(s11725, c11725, in11725_1, in11725_2, s9849[0]);
    wire[0:0] s11726, in11726_1, in11726_2;
    wire c11726;
    assign in11726_1 = {s9853[0]};
    assign in11726_2 = {s9854[0]};
    Full_Adder FA_11726(s11726, c11726, in11726_1, in11726_2, s9852[0]);
    wire[0:0] s11727, in11727_1, in11727_2;
    wire c11727;
    assign in11727_1 = {c9845};
    assign in11727_2 = {c9846};
    Full_Adder FA_11727(s11727, c11727, in11727_1, in11727_2, c9844);
    wire[0:0] s11728, in11728_1, in11728_2;
    wire c11728;
    assign in11728_1 = {c9848};
    assign in11728_2 = {c9849};
    Full_Adder FA_11728(s11728, c11728, in11728_1, in11728_2, c9847);
    wire[0:0] s11729, in11729_1, in11729_2;
    wire c11729;
    assign in11729_1 = {c9851};
    assign in11729_2 = {c9852};
    Full_Adder FA_11729(s11729, c11729, in11729_1, in11729_2, c9850);
    wire[0:0] s11730, in11730_1, in11730_2;
    wire c11730;
    assign in11730_1 = {c9854};
    assign in11730_2 = {c9855};
    Full_Adder FA_11730(s11730, c11730, in11730_1, in11730_2, c9853);
    wire[0:0] s11731, in11731_1, in11731_2;
    wire c11731;
    assign in11731_1 = {s9857[0]};
    assign in11731_2 = {s9858[0]};
    Full_Adder FA_11731(s11731, c11731, in11731_1, in11731_2, c9856);
    wire[0:0] s11732, in11732_1, in11732_2;
    wire c11732;
    assign in11732_1 = {s9860[0]};
    assign in11732_2 = {s9861[0]};
    Full_Adder FA_11732(s11732, c11732, in11732_1, in11732_2, s9859[0]);
    wire[0:0] s11733, in11733_1, in11733_2;
    wire c11733;
    assign in11733_1 = {s9863[0]};
    assign in11733_2 = {s9864[0]};
    Full_Adder FA_11733(s11733, c11733, in11733_1, in11733_2, s9862[0]);
    wire[0:0] s11734, in11734_1, in11734_2;
    wire c11734;
    assign in11734_1 = {s9866[0]};
    assign in11734_2 = {s9867[0]};
    Full_Adder FA_11734(s11734, c11734, in11734_1, in11734_2, s9865[0]);
    wire[0:0] s11735, in11735_1, in11735_2;
    wire c11735;
    assign in11735_1 = {c9858};
    assign in11735_2 = {c9859};
    Full_Adder FA_11735(s11735, c11735, in11735_1, in11735_2, c9857);
    wire[0:0] s11736, in11736_1, in11736_2;
    wire c11736;
    assign in11736_1 = {c9861};
    assign in11736_2 = {c9862};
    Full_Adder FA_11736(s11736, c11736, in11736_1, in11736_2, c9860);
    wire[0:0] s11737, in11737_1, in11737_2;
    wire c11737;
    assign in11737_1 = {c9864};
    assign in11737_2 = {c9865};
    Full_Adder FA_11737(s11737, c11737, in11737_1, in11737_2, c9863);
    wire[0:0] s11738, in11738_1, in11738_2;
    wire c11738;
    assign in11738_1 = {c9867};
    assign in11738_2 = {c9868};
    Full_Adder FA_11738(s11738, c11738, in11738_1, in11738_2, c9866);
    wire[0:0] s11739, in11739_1, in11739_2;
    wire c11739;
    assign in11739_1 = {s9870[0]};
    assign in11739_2 = {s9871[0]};
    Full_Adder FA_11739(s11739, c11739, in11739_1, in11739_2, c9869);
    wire[0:0] s11740, in11740_1, in11740_2;
    wire c11740;
    assign in11740_1 = {s9873[0]};
    assign in11740_2 = {s9874[0]};
    Full_Adder FA_11740(s11740, c11740, in11740_1, in11740_2, s9872[0]);
    wire[0:0] s11741, in11741_1, in11741_2;
    wire c11741;
    assign in11741_1 = {s9876[0]};
    assign in11741_2 = {s9877[0]};
    Full_Adder FA_11741(s11741, c11741, in11741_1, in11741_2, s9875[0]);
    wire[0:0] s11742, in11742_1, in11742_2;
    wire c11742;
    assign in11742_1 = {s9879[0]};
    assign in11742_2 = {s9880[0]};
    Full_Adder FA_11742(s11742, c11742, in11742_1, in11742_2, s9878[0]);
    wire[0:0] s11743, in11743_1, in11743_2;
    wire c11743;
    assign in11743_1 = {c9871};
    assign in11743_2 = {c9872};
    Full_Adder FA_11743(s11743, c11743, in11743_1, in11743_2, c9870);
    wire[0:0] s11744, in11744_1, in11744_2;
    wire c11744;
    assign in11744_1 = {c9874};
    assign in11744_2 = {c9875};
    Full_Adder FA_11744(s11744, c11744, in11744_1, in11744_2, c9873);
    wire[0:0] s11745, in11745_1, in11745_2;
    wire c11745;
    assign in11745_1 = {c9877};
    assign in11745_2 = {c9878};
    Full_Adder FA_11745(s11745, c11745, in11745_1, in11745_2, c9876);
    wire[0:0] s11746, in11746_1, in11746_2;
    wire c11746;
    assign in11746_1 = {c9880};
    assign in11746_2 = {c9881};
    Full_Adder FA_11746(s11746, c11746, in11746_1, in11746_2, c9879);
    wire[0:0] s11747, in11747_1, in11747_2;
    wire c11747;
    assign in11747_1 = {s9883[0]};
    assign in11747_2 = {s9884[0]};
    Full_Adder FA_11747(s11747, c11747, in11747_1, in11747_2, c9882);
    wire[0:0] s11748, in11748_1, in11748_2;
    wire c11748;
    assign in11748_1 = {s9886[0]};
    assign in11748_2 = {s9887[0]};
    Full_Adder FA_11748(s11748, c11748, in11748_1, in11748_2, s9885[0]);
    wire[0:0] s11749, in11749_1, in11749_2;
    wire c11749;
    assign in11749_1 = {s9889[0]};
    assign in11749_2 = {s9890[0]};
    Full_Adder FA_11749(s11749, c11749, in11749_1, in11749_2, s9888[0]);
    wire[0:0] s11750, in11750_1, in11750_2;
    wire c11750;
    assign in11750_1 = {s9892[0]};
    assign in11750_2 = {s9893[0]};
    Full_Adder FA_11750(s11750, c11750, in11750_1, in11750_2, s9891[0]);
    wire[0:0] s11751, in11751_1, in11751_2;
    wire c11751;
    assign in11751_1 = {c9884};
    assign in11751_2 = {c9885};
    Full_Adder FA_11751(s11751, c11751, in11751_1, in11751_2, c9883);
    wire[0:0] s11752, in11752_1, in11752_2;
    wire c11752;
    assign in11752_1 = {c9887};
    assign in11752_2 = {c9888};
    Full_Adder FA_11752(s11752, c11752, in11752_1, in11752_2, c9886);
    wire[0:0] s11753, in11753_1, in11753_2;
    wire c11753;
    assign in11753_1 = {c9890};
    assign in11753_2 = {c9891};
    Full_Adder FA_11753(s11753, c11753, in11753_1, in11753_2, c9889);
    wire[0:0] s11754, in11754_1, in11754_2;
    wire c11754;
    assign in11754_1 = {c9893};
    assign in11754_2 = {c9894};
    Full_Adder FA_11754(s11754, c11754, in11754_1, in11754_2, c9892);
    wire[0:0] s11755, in11755_1, in11755_2;
    wire c11755;
    assign in11755_1 = {s9896[0]};
    assign in11755_2 = {s9897[0]};
    Full_Adder FA_11755(s11755, c11755, in11755_1, in11755_2, c9895);
    wire[0:0] s11756, in11756_1, in11756_2;
    wire c11756;
    assign in11756_1 = {s9899[0]};
    assign in11756_2 = {s9900[0]};
    Full_Adder FA_11756(s11756, c11756, in11756_1, in11756_2, s9898[0]);
    wire[0:0] s11757, in11757_1, in11757_2;
    wire c11757;
    assign in11757_1 = {s9902[0]};
    assign in11757_2 = {s9903[0]};
    Full_Adder FA_11757(s11757, c11757, in11757_1, in11757_2, s9901[0]);
    wire[0:0] s11758, in11758_1, in11758_2;
    wire c11758;
    assign in11758_1 = {s9905[0]};
    assign in11758_2 = {s9906[0]};
    Full_Adder FA_11758(s11758, c11758, in11758_1, in11758_2, s9904[0]);
    wire[0:0] s11759, in11759_1, in11759_2;
    wire c11759;
    assign in11759_1 = {c9897};
    assign in11759_2 = {c9898};
    Full_Adder FA_11759(s11759, c11759, in11759_1, in11759_2, c9896);
    wire[0:0] s11760, in11760_1, in11760_2;
    wire c11760;
    assign in11760_1 = {c9900};
    assign in11760_2 = {c9901};
    Full_Adder FA_11760(s11760, c11760, in11760_1, in11760_2, c9899);
    wire[0:0] s11761, in11761_1, in11761_2;
    wire c11761;
    assign in11761_1 = {c9903};
    assign in11761_2 = {c9904};
    Full_Adder FA_11761(s11761, c11761, in11761_1, in11761_2, c9902);
    wire[0:0] s11762, in11762_1, in11762_2;
    wire c11762;
    assign in11762_1 = {c9906};
    assign in11762_2 = {c9907};
    Full_Adder FA_11762(s11762, c11762, in11762_1, in11762_2, c9905);
    wire[0:0] s11763, in11763_1, in11763_2;
    wire c11763;
    assign in11763_1 = {s9909[0]};
    assign in11763_2 = {s9910[0]};
    Full_Adder FA_11763(s11763, c11763, in11763_1, in11763_2, c9908);
    wire[0:0] s11764, in11764_1, in11764_2;
    wire c11764;
    assign in11764_1 = {s9912[0]};
    assign in11764_2 = {s9913[0]};
    Full_Adder FA_11764(s11764, c11764, in11764_1, in11764_2, s9911[0]);
    wire[0:0] s11765, in11765_1, in11765_2;
    wire c11765;
    assign in11765_1 = {s9915[0]};
    assign in11765_2 = {s9916[0]};
    Full_Adder FA_11765(s11765, c11765, in11765_1, in11765_2, s9914[0]);
    wire[0:0] s11766, in11766_1, in11766_2;
    wire c11766;
    assign in11766_1 = {s9918[0]};
    assign in11766_2 = {s9919[0]};
    Full_Adder FA_11766(s11766, c11766, in11766_1, in11766_2, s9917[0]);
    wire[0:0] s11767, in11767_1, in11767_2;
    wire c11767;
    assign in11767_1 = {c9910};
    assign in11767_2 = {c9911};
    Full_Adder FA_11767(s11767, c11767, in11767_1, in11767_2, c9909);
    wire[0:0] s11768, in11768_1, in11768_2;
    wire c11768;
    assign in11768_1 = {c9913};
    assign in11768_2 = {c9914};
    Full_Adder FA_11768(s11768, c11768, in11768_1, in11768_2, c9912);
    wire[0:0] s11769, in11769_1, in11769_2;
    wire c11769;
    assign in11769_1 = {c9916};
    assign in11769_2 = {c9917};
    Full_Adder FA_11769(s11769, c11769, in11769_1, in11769_2, c9915);
    wire[0:0] s11770, in11770_1, in11770_2;
    wire c11770;
    assign in11770_1 = {c9919};
    assign in11770_2 = {c9920};
    Full_Adder FA_11770(s11770, c11770, in11770_1, in11770_2, c9918);
    wire[0:0] s11771, in11771_1, in11771_2;
    wire c11771;
    assign in11771_1 = {s9922[0]};
    assign in11771_2 = {s9923[0]};
    Full_Adder FA_11771(s11771, c11771, in11771_1, in11771_2, c9921);
    wire[0:0] s11772, in11772_1, in11772_2;
    wire c11772;
    assign in11772_1 = {s9925[0]};
    assign in11772_2 = {s9926[0]};
    Full_Adder FA_11772(s11772, c11772, in11772_1, in11772_2, s9924[0]);
    wire[0:0] s11773, in11773_1, in11773_2;
    wire c11773;
    assign in11773_1 = {s9928[0]};
    assign in11773_2 = {s9929[0]};
    Full_Adder FA_11773(s11773, c11773, in11773_1, in11773_2, s9927[0]);
    wire[0:0] s11774, in11774_1, in11774_2;
    wire c11774;
    assign in11774_1 = {s9931[0]};
    assign in11774_2 = {s9932[0]};
    Full_Adder FA_11774(s11774, c11774, in11774_1, in11774_2, s9930[0]);
    wire[0:0] s11775, in11775_1, in11775_2;
    wire c11775;
    assign in11775_1 = {c9923};
    assign in11775_2 = {c9924};
    Full_Adder FA_11775(s11775, c11775, in11775_1, in11775_2, c9922);
    wire[0:0] s11776, in11776_1, in11776_2;
    wire c11776;
    assign in11776_1 = {c9926};
    assign in11776_2 = {c9927};
    Full_Adder FA_11776(s11776, c11776, in11776_1, in11776_2, c9925);
    wire[0:0] s11777, in11777_1, in11777_2;
    wire c11777;
    assign in11777_1 = {c9929};
    assign in11777_2 = {c9930};
    Full_Adder FA_11777(s11777, c11777, in11777_1, in11777_2, c9928);
    wire[0:0] s11778, in11778_1, in11778_2;
    wire c11778;
    assign in11778_1 = {c9932};
    assign in11778_2 = {c9933};
    Full_Adder FA_11778(s11778, c11778, in11778_1, in11778_2, c9931);
    wire[0:0] s11779, in11779_1, in11779_2;
    wire c11779;
    assign in11779_1 = {s9935[0]};
    assign in11779_2 = {s9936[0]};
    Full_Adder FA_11779(s11779, c11779, in11779_1, in11779_2, c9934);
    wire[0:0] s11780, in11780_1, in11780_2;
    wire c11780;
    assign in11780_1 = {s9938[0]};
    assign in11780_2 = {s9939[0]};
    Full_Adder FA_11780(s11780, c11780, in11780_1, in11780_2, s9937[0]);
    wire[0:0] s11781, in11781_1, in11781_2;
    wire c11781;
    assign in11781_1 = {s9941[0]};
    assign in11781_2 = {s9942[0]};
    Full_Adder FA_11781(s11781, c11781, in11781_1, in11781_2, s9940[0]);
    wire[0:0] s11782, in11782_1, in11782_2;
    wire c11782;
    assign in11782_1 = {s9944[0]};
    assign in11782_2 = {s9945[0]};
    Full_Adder FA_11782(s11782, c11782, in11782_1, in11782_2, s9943[0]);
    wire[0:0] s11783, in11783_1, in11783_2;
    wire c11783;
    assign in11783_1 = {c9936};
    assign in11783_2 = {c9937};
    Full_Adder FA_11783(s11783, c11783, in11783_1, in11783_2, c9935);
    wire[0:0] s11784, in11784_1, in11784_2;
    wire c11784;
    assign in11784_1 = {c9939};
    assign in11784_2 = {c9940};
    Full_Adder FA_11784(s11784, c11784, in11784_1, in11784_2, c9938);
    wire[0:0] s11785, in11785_1, in11785_2;
    wire c11785;
    assign in11785_1 = {c9942};
    assign in11785_2 = {c9943};
    Full_Adder FA_11785(s11785, c11785, in11785_1, in11785_2, c9941);
    wire[0:0] s11786, in11786_1, in11786_2;
    wire c11786;
    assign in11786_1 = {c9945};
    assign in11786_2 = {c9946};
    Full_Adder FA_11786(s11786, c11786, in11786_1, in11786_2, c9944);
    wire[0:0] s11787, in11787_1, in11787_2;
    wire c11787;
    assign in11787_1 = {s9948[0]};
    assign in11787_2 = {s9949[0]};
    Full_Adder FA_11787(s11787, c11787, in11787_1, in11787_2, c9947);
    wire[0:0] s11788, in11788_1, in11788_2;
    wire c11788;
    assign in11788_1 = {s9951[0]};
    assign in11788_2 = {s9952[0]};
    Full_Adder FA_11788(s11788, c11788, in11788_1, in11788_2, s9950[0]);
    wire[0:0] s11789, in11789_1, in11789_2;
    wire c11789;
    assign in11789_1 = {s9954[0]};
    assign in11789_2 = {s9955[0]};
    Full_Adder FA_11789(s11789, c11789, in11789_1, in11789_2, s9953[0]);
    wire[0:0] s11790, in11790_1, in11790_2;
    wire c11790;
    assign in11790_1 = {s9957[0]};
    assign in11790_2 = {s9958[0]};
    Full_Adder FA_11790(s11790, c11790, in11790_1, in11790_2, s9956[0]);
    wire[0:0] s11791, in11791_1, in11791_2;
    wire c11791;
    assign in11791_1 = {c9949};
    assign in11791_2 = {c9950};
    Full_Adder FA_11791(s11791, c11791, in11791_1, in11791_2, c9948);
    wire[0:0] s11792, in11792_1, in11792_2;
    wire c11792;
    assign in11792_1 = {c9952};
    assign in11792_2 = {c9953};
    Full_Adder FA_11792(s11792, c11792, in11792_1, in11792_2, c9951);
    wire[0:0] s11793, in11793_1, in11793_2;
    wire c11793;
    assign in11793_1 = {c9955};
    assign in11793_2 = {c9956};
    Full_Adder FA_11793(s11793, c11793, in11793_1, in11793_2, c9954);
    wire[0:0] s11794, in11794_1, in11794_2;
    wire c11794;
    assign in11794_1 = {c9958};
    assign in11794_2 = {c9959};
    Full_Adder FA_11794(s11794, c11794, in11794_1, in11794_2, c9957);
    wire[0:0] s11795, in11795_1, in11795_2;
    wire c11795;
    assign in11795_1 = {s9961[0]};
    assign in11795_2 = {s9962[0]};
    Full_Adder FA_11795(s11795, c11795, in11795_1, in11795_2, c9960);
    wire[0:0] s11796, in11796_1, in11796_2;
    wire c11796;
    assign in11796_1 = {s9964[0]};
    assign in11796_2 = {s9965[0]};
    Full_Adder FA_11796(s11796, c11796, in11796_1, in11796_2, s9963[0]);
    wire[0:0] s11797, in11797_1, in11797_2;
    wire c11797;
    assign in11797_1 = {s9967[0]};
    assign in11797_2 = {s9968[0]};
    Full_Adder FA_11797(s11797, c11797, in11797_1, in11797_2, s9966[0]);
    wire[0:0] s11798, in11798_1, in11798_2;
    wire c11798;
    assign in11798_1 = {s9970[0]};
    assign in11798_2 = {s9971[0]};
    Full_Adder FA_11798(s11798, c11798, in11798_1, in11798_2, s9969[0]);
    wire[0:0] s11799, in11799_1, in11799_2;
    wire c11799;
    assign in11799_1 = {c9962};
    assign in11799_2 = {c9963};
    Full_Adder FA_11799(s11799, c11799, in11799_1, in11799_2, c9961);
    wire[0:0] s11800, in11800_1, in11800_2;
    wire c11800;
    assign in11800_1 = {c9965};
    assign in11800_2 = {c9966};
    Full_Adder FA_11800(s11800, c11800, in11800_1, in11800_2, c9964);
    wire[0:0] s11801, in11801_1, in11801_2;
    wire c11801;
    assign in11801_1 = {c9968};
    assign in11801_2 = {c9969};
    Full_Adder FA_11801(s11801, c11801, in11801_1, in11801_2, c9967);
    wire[0:0] s11802, in11802_1, in11802_2;
    wire c11802;
    assign in11802_1 = {c9971};
    assign in11802_2 = {c9972};
    Full_Adder FA_11802(s11802, c11802, in11802_1, in11802_2, c9970);
    wire[0:0] s11803, in11803_1, in11803_2;
    wire c11803;
    assign in11803_1 = {s9974[0]};
    assign in11803_2 = {s9975[0]};
    Full_Adder FA_11803(s11803, c11803, in11803_1, in11803_2, c9973);
    wire[0:0] s11804, in11804_1, in11804_2;
    wire c11804;
    assign in11804_1 = {s9977[0]};
    assign in11804_2 = {s9978[0]};
    Full_Adder FA_11804(s11804, c11804, in11804_1, in11804_2, s9976[0]);
    wire[0:0] s11805, in11805_1, in11805_2;
    wire c11805;
    assign in11805_1 = {s9980[0]};
    assign in11805_2 = {s9981[0]};
    Full_Adder FA_11805(s11805, c11805, in11805_1, in11805_2, s9979[0]);
    wire[0:0] s11806, in11806_1, in11806_2;
    wire c11806;
    assign in11806_1 = {s9983[0]};
    assign in11806_2 = {s9984[0]};
    Full_Adder FA_11806(s11806, c11806, in11806_1, in11806_2, s9982[0]);
    wire[0:0] s11807, in11807_1, in11807_2;
    wire c11807;
    assign in11807_1 = {c9975};
    assign in11807_2 = {c9976};
    Full_Adder FA_11807(s11807, c11807, in11807_1, in11807_2, c9974);
    wire[0:0] s11808, in11808_1, in11808_2;
    wire c11808;
    assign in11808_1 = {c9978};
    assign in11808_2 = {c9979};
    Full_Adder FA_11808(s11808, c11808, in11808_1, in11808_2, c9977);
    wire[0:0] s11809, in11809_1, in11809_2;
    wire c11809;
    assign in11809_1 = {c9981};
    assign in11809_2 = {c9982};
    Full_Adder FA_11809(s11809, c11809, in11809_1, in11809_2, c9980);
    wire[0:0] s11810, in11810_1, in11810_2;
    wire c11810;
    assign in11810_1 = {c9984};
    assign in11810_2 = {c9985};
    Full_Adder FA_11810(s11810, c11810, in11810_1, in11810_2, c9983);
    wire[0:0] s11811, in11811_1, in11811_2;
    wire c11811;
    assign in11811_1 = {s9987[0]};
    assign in11811_2 = {s9988[0]};
    Full_Adder FA_11811(s11811, c11811, in11811_1, in11811_2, c9986);
    wire[0:0] s11812, in11812_1, in11812_2;
    wire c11812;
    assign in11812_1 = {s9990[0]};
    assign in11812_2 = {s9991[0]};
    Full_Adder FA_11812(s11812, c11812, in11812_1, in11812_2, s9989[0]);
    wire[0:0] s11813, in11813_1, in11813_2;
    wire c11813;
    assign in11813_1 = {s9993[0]};
    assign in11813_2 = {s9994[0]};
    Full_Adder FA_11813(s11813, c11813, in11813_1, in11813_2, s9992[0]);
    wire[0:0] s11814, in11814_1, in11814_2;
    wire c11814;
    assign in11814_1 = {s9996[0]};
    assign in11814_2 = {s9997[0]};
    Full_Adder FA_11814(s11814, c11814, in11814_1, in11814_2, s9995[0]);
    wire[0:0] s11815, in11815_1, in11815_2;
    wire c11815;
    assign in11815_1 = {c9988};
    assign in11815_2 = {c9989};
    Full_Adder FA_11815(s11815, c11815, in11815_1, in11815_2, c9987);
    wire[0:0] s11816, in11816_1, in11816_2;
    wire c11816;
    assign in11816_1 = {c9991};
    assign in11816_2 = {c9992};
    Full_Adder FA_11816(s11816, c11816, in11816_1, in11816_2, c9990);
    wire[0:0] s11817, in11817_1, in11817_2;
    wire c11817;
    assign in11817_1 = {c9994};
    assign in11817_2 = {c9995};
    Full_Adder FA_11817(s11817, c11817, in11817_1, in11817_2, c9993);
    wire[0:0] s11818, in11818_1, in11818_2;
    wire c11818;
    assign in11818_1 = {c9997};
    assign in11818_2 = {c9998};
    Full_Adder FA_11818(s11818, c11818, in11818_1, in11818_2, c9996);
    wire[0:0] s11819, in11819_1, in11819_2;
    wire c11819;
    assign in11819_1 = {s10000[0]};
    assign in11819_2 = {s10001[0]};
    Full_Adder FA_11819(s11819, c11819, in11819_1, in11819_2, c9999);
    wire[0:0] s11820, in11820_1, in11820_2;
    wire c11820;
    assign in11820_1 = {s10003[0]};
    assign in11820_2 = {s10004[0]};
    Full_Adder FA_11820(s11820, c11820, in11820_1, in11820_2, s10002[0]);
    wire[0:0] s11821, in11821_1, in11821_2;
    wire c11821;
    assign in11821_1 = {s10006[0]};
    assign in11821_2 = {s10007[0]};
    Full_Adder FA_11821(s11821, c11821, in11821_1, in11821_2, s10005[0]);
    wire[0:0] s11822, in11822_1, in11822_2;
    wire c11822;
    assign in11822_1 = {s10009[0]};
    assign in11822_2 = {s10010[0]};
    Full_Adder FA_11822(s11822, c11822, in11822_1, in11822_2, s10008[0]);
    wire[0:0] s11823, in11823_1, in11823_2;
    wire c11823;
    assign in11823_1 = {c10001};
    assign in11823_2 = {c10002};
    Full_Adder FA_11823(s11823, c11823, in11823_1, in11823_2, c10000);
    wire[0:0] s11824, in11824_1, in11824_2;
    wire c11824;
    assign in11824_1 = {c10004};
    assign in11824_2 = {c10005};
    Full_Adder FA_11824(s11824, c11824, in11824_1, in11824_2, c10003);
    wire[0:0] s11825, in11825_1, in11825_2;
    wire c11825;
    assign in11825_1 = {c10007};
    assign in11825_2 = {c10008};
    Full_Adder FA_11825(s11825, c11825, in11825_1, in11825_2, c10006);
    wire[0:0] s11826, in11826_1, in11826_2;
    wire c11826;
    assign in11826_1 = {c10010};
    assign in11826_2 = {c10011};
    Full_Adder FA_11826(s11826, c11826, in11826_1, in11826_2, c10009);
    wire[0:0] s11827, in11827_1, in11827_2;
    wire c11827;
    assign in11827_1 = {s10013[0]};
    assign in11827_2 = {s10014[0]};
    Full_Adder FA_11827(s11827, c11827, in11827_1, in11827_2, c10012);
    wire[0:0] s11828, in11828_1, in11828_2;
    wire c11828;
    assign in11828_1 = {s10016[0]};
    assign in11828_2 = {s10017[0]};
    Full_Adder FA_11828(s11828, c11828, in11828_1, in11828_2, s10015[0]);
    wire[0:0] s11829, in11829_1, in11829_2;
    wire c11829;
    assign in11829_1 = {s10019[0]};
    assign in11829_2 = {s10020[0]};
    Full_Adder FA_11829(s11829, c11829, in11829_1, in11829_2, s10018[0]);
    wire[0:0] s11830, in11830_1, in11830_2;
    wire c11830;
    assign in11830_1 = {s10022[0]};
    assign in11830_2 = {s10023[0]};
    Full_Adder FA_11830(s11830, c11830, in11830_1, in11830_2, s10021[0]);
    wire[0:0] s11831, in11831_1, in11831_2;
    wire c11831;
    assign in11831_1 = {c10014};
    assign in11831_2 = {c10015};
    Full_Adder FA_11831(s11831, c11831, in11831_1, in11831_2, c10013);
    wire[0:0] s11832, in11832_1, in11832_2;
    wire c11832;
    assign in11832_1 = {c10017};
    assign in11832_2 = {c10018};
    Full_Adder FA_11832(s11832, c11832, in11832_1, in11832_2, c10016);
    wire[0:0] s11833, in11833_1, in11833_2;
    wire c11833;
    assign in11833_1 = {c10020};
    assign in11833_2 = {c10021};
    Full_Adder FA_11833(s11833, c11833, in11833_1, in11833_2, c10019);
    wire[0:0] s11834, in11834_1, in11834_2;
    wire c11834;
    assign in11834_1 = {c10023};
    assign in11834_2 = {c10024};
    Full_Adder FA_11834(s11834, c11834, in11834_1, in11834_2, c10022);
    wire[0:0] s11835, in11835_1, in11835_2;
    wire c11835;
    assign in11835_1 = {s10026[0]};
    assign in11835_2 = {s10027[0]};
    Full_Adder FA_11835(s11835, c11835, in11835_1, in11835_2, c10025);
    wire[0:0] s11836, in11836_1, in11836_2;
    wire c11836;
    assign in11836_1 = {s10029[0]};
    assign in11836_2 = {s10030[0]};
    Full_Adder FA_11836(s11836, c11836, in11836_1, in11836_2, s10028[0]);
    wire[0:0] s11837, in11837_1, in11837_2;
    wire c11837;
    assign in11837_1 = {s10032[0]};
    assign in11837_2 = {s10033[0]};
    Full_Adder FA_11837(s11837, c11837, in11837_1, in11837_2, s10031[0]);
    wire[0:0] s11838, in11838_1, in11838_2;
    wire c11838;
    assign in11838_1 = {s10035[0]};
    assign in11838_2 = {s10036[0]};
    Full_Adder FA_11838(s11838, c11838, in11838_1, in11838_2, s10034[0]);
    wire[0:0] s11839, in11839_1, in11839_2;
    wire c11839;
    assign in11839_1 = {c10027};
    assign in11839_2 = {c10028};
    Full_Adder FA_11839(s11839, c11839, in11839_1, in11839_2, c10026);
    wire[0:0] s11840, in11840_1, in11840_2;
    wire c11840;
    assign in11840_1 = {c10030};
    assign in11840_2 = {c10031};
    Full_Adder FA_11840(s11840, c11840, in11840_1, in11840_2, c10029);
    wire[0:0] s11841, in11841_1, in11841_2;
    wire c11841;
    assign in11841_1 = {c10033};
    assign in11841_2 = {c10034};
    Full_Adder FA_11841(s11841, c11841, in11841_1, in11841_2, c10032);
    wire[0:0] s11842, in11842_1, in11842_2;
    wire c11842;
    assign in11842_1 = {c10036};
    assign in11842_2 = {c10037};
    Full_Adder FA_11842(s11842, c11842, in11842_1, in11842_2, c10035);
    wire[0:0] s11843, in11843_1, in11843_2;
    wire c11843;
    assign in11843_1 = {s10039[0]};
    assign in11843_2 = {s10040[0]};
    Full_Adder FA_11843(s11843, c11843, in11843_1, in11843_2, c10038);
    wire[0:0] s11844, in11844_1, in11844_2;
    wire c11844;
    assign in11844_1 = {s10042[0]};
    assign in11844_2 = {s10043[0]};
    Full_Adder FA_11844(s11844, c11844, in11844_1, in11844_2, s10041[0]);
    wire[0:0] s11845, in11845_1, in11845_2;
    wire c11845;
    assign in11845_1 = {s10045[0]};
    assign in11845_2 = {s10046[0]};
    Full_Adder FA_11845(s11845, c11845, in11845_1, in11845_2, s10044[0]);
    wire[0:0] s11846, in11846_1, in11846_2;
    wire c11846;
    assign in11846_1 = {s10048[0]};
    assign in11846_2 = {s10049[0]};
    Full_Adder FA_11846(s11846, c11846, in11846_1, in11846_2, s10047[0]);
    wire[0:0] s11847, in11847_1, in11847_2;
    wire c11847;
    assign in11847_1 = {c10040};
    assign in11847_2 = {c10041};
    Full_Adder FA_11847(s11847, c11847, in11847_1, in11847_2, c10039);
    wire[0:0] s11848, in11848_1, in11848_2;
    wire c11848;
    assign in11848_1 = {c10043};
    assign in11848_2 = {c10044};
    Full_Adder FA_11848(s11848, c11848, in11848_1, in11848_2, c10042);
    wire[0:0] s11849, in11849_1, in11849_2;
    wire c11849;
    assign in11849_1 = {c10046};
    assign in11849_2 = {c10047};
    Full_Adder FA_11849(s11849, c11849, in11849_1, in11849_2, c10045);
    wire[0:0] s11850, in11850_1, in11850_2;
    wire c11850;
    assign in11850_1 = {c10049};
    assign in11850_2 = {c10050};
    Full_Adder FA_11850(s11850, c11850, in11850_1, in11850_2, c10048);
    wire[0:0] s11851, in11851_1, in11851_2;
    wire c11851;
    assign in11851_1 = {s10052[0]};
    assign in11851_2 = {s10053[0]};
    Full_Adder FA_11851(s11851, c11851, in11851_1, in11851_2, c10051);
    wire[0:0] s11852, in11852_1, in11852_2;
    wire c11852;
    assign in11852_1 = {s10055[0]};
    assign in11852_2 = {s10056[0]};
    Full_Adder FA_11852(s11852, c11852, in11852_1, in11852_2, s10054[0]);
    wire[0:0] s11853, in11853_1, in11853_2;
    wire c11853;
    assign in11853_1 = {s10058[0]};
    assign in11853_2 = {s10059[0]};
    Full_Adder FA_11853(s11853, c11853, in11853_1, in11853_2, s10057[0]);
    wire[0:0] s11854, in11854_1, in11854_2;
    wire c11854;
    assign in11854_1 = {s10061[0]};
    assign in11854_2 = {s10062[0]};
    Full_Adder FA_11854(s11854, c11854, in11854_1, in11854_2, s10060[0]);
    wire[0:0] s11855, in11855_1, in11855_2;
    wire c11855;
    assign in11855_1 = {c10053};
    assign in11855_2 = {c10054};
    Full_Adder FA_11855(s11855, c11855, in11855_1, in11855_2, c10052);
    wire[0:0] s11856, in11856_1, in11856_2;
    wire c11856;
    assign in11856_1 = {c10056};
    assign in11856_2 = {c10057};
    Full_Adder FA_11856(s11856, c11856, in11856_1, in11856_2, c10055);
    wire[0:0] s11857, in11857_1, in11857_2;
    wire c11857;
    assign in11857_1 = {c10059};
    assign in11857_2 = {c10060};
    Full_Adder FA_11857(s11857, c11857, in11857_1, in11857_2, c10058);
    wire[0:0] s11858, in11858_1, in11858_2;
    wire c11858;
    assign in11858_1 = {c10062};
    assign in11858_2 = {c10063};
    Full_Adder FA_11858(s11858, c11858, in11858_1, in11858_2, c10061);
    wire[0:0] s11859, in11859_1, in11859_2;
    wire c11859;
    assign in11859_1 = {s10065[0]};
    assign in11859_2 = {s10066[0]};
    Full_Adder FA_11859(s11859, c11859, in11859_1, in11859_2, c10064);
    wire[0:0] s11860, in11860_1, in11860_2;
    wire c11860;
    assign in11860_1 = {s10068[0]};
    assign in11860_2 = {s10069[0]};
    Full_Adder FA_11860(s11860, c11860, in11860_1, in11860_2, s10067[0]);
    wire[0:0] s11861, in11861_1, in11861_2;
    wire c11861;
    assign in11861_1 = {s10071[0]};
    assign in11861_2 = {s10072[0]};
    Full_Adder FA_11861(s11861, c11861, in11861_1, in11861_2, s10070[0]);
    wire[0:0] s11862, in11862_1, in11862_2;
    wire c11862;
    assign in11862_1 = {s10074[0]};
    assign in11862_2 = {s10075[0]};
    Full_Adder FA_11862(s11862, c11862, in11862_1, in11862_2, s10073[0]);
    wire[0:0] s11863, in11863_1, in11863_2;
    wire c11863;
    assign in11863_1 = {c10066};
    assign in11863_2 = {c10067};
    Full_Adder FA_11863(s11863, c11863, in11863_1, in11863_2, c10065);
    wire[0:0] s11864, in11864_1, in11864_2;
    wire c11864;
    assign in11864_1 = {c10069};
    assign in11864_2 = {c10070};
    Full_Adder FA_11864(s11864, c11864, in11864_1, in11864_2, c10068);
    wire[0:0] s11865, in11865_1, in11865_2;
    wire c11865;
    assign in11865_1 = {c10072};
    assign in11865_2 = {c10073};
    Full_Adder FA_11865(s11865, c11865, in11865_1, in11865_2, c10071);
    wire[0:0] s11866, in11866_1, in11866_2;
    wire c11866;
    assign in11866_1 = {c10075};
    assign in11866_2 = {c10076};
    Full_Adder FA_11866(s11866, c11866, in11866_1, in11866_2, c10074);
    wire[0:0] s11867, in11867_1, in11867_2;
    wire c11867;
    assign in11867_1 = {s10078[0]};
    assign in11867_2 = {s10079[0]};
    Full_Adder FA_11867(s11867, c11867, in11867_1, in11867_2, c10077);
    wire[0:0] s11868, in11868_1, in11868_2;
    wire c11868;
    assign in11868_1 = {s10081[0]};
    assign in11868_2 = {s10082[0]};
    Full_Adder FA_11868(s11868, c11868, in11868_1, in11868_2, s10080[0]);
    wire[0:0] s11869, in11869_1, in11869_2;
    wire c11869;
    assign in11869_1 = {s10084[0]};
    assign in11869_2 = {s10085[0]};
    Full_Adder FA_11869(s11869, c11869, in11869_1, in11869_2, s10083[0]);
    wire[0:0] s11870, in11870_1, in11870_2;
    wire c11870;
    assign in11870_1 = {s10087[0]};
    assign in11870_2 = {s10088[0]};
    Full_Adder FA_11870(s11870, c11870, in11870_1, in11870_2, s10086[0]);
    wire[0:0] s11871, in11871_1, in11871_2;
    wire c11871;
    assign in11871_1 = {c10079};
    assign in11871_2 = {c10080};
    Full_Adder FA_11871(s11871, c11871, in11871_1, in11871_2, c10078);
    wire[0:0] s11872, in11872_1, in11872_2;
    wire c11872;
    assign in11872_1 = {c10082};
    assign in11872_2 = {c10083};
    Full_Adder FA_11872(s11872, c11872, in11872_1, in11872_2, c10081);
    wire[0:0] s11873, in11873_1, in11873_2;
    wire c11873;
    assign in11873_1 = {c10085};
    assign in11873_2 = {c10086};
    Full_Adder FA_11873(s11873, c11873, in11873_1, in11873_2, c10084);
    wire[0:0] s11874, in11874_1, in11874_2;
    wire c11874;
    assign in11874_1 = {c10088};
    assign in11874_2 = {c10089};
    Full_Adder FA_11874(s11874, c11874, in11874_1, in11874_2, c10087);
    wire[0:0] s11875, in11875_1, in11875_2;
    wire c11875;
    assign in11875_1 = {s10091[0]};
    assign in11875_2 = {s10092[0]};
    Full_Adder FA_11875(s11875, c11875, in11875_1, in11875_2, c10090);
    wire[0:0] s11876, in11876_1, in11876_2;
    wire c11876;
    assign in11876_1 = {s10094[0]};
    assign in11876_2 = {s10095[0]};
    Full_Adder FA_11876(s11876, c11876, in11876_1, in11876_2, s10093[0]);
    wire[0:0] s11877, in11877_1, in11877_2;
    wire c11877;
    assign in11877_1 = {s10097[0]};
    assign in11877_2 = {s10098[0]};
    Full_Adder FA_11877(s11877, c11877, in11877_1, in11877_2, s10096[0]);
    wire[0:0] s11878, in11878_1, in11878_2;
    wire c11878;
    assign in11878_1 = {s10100[0]};
    assign in11878_2 = {s10101[0]};
    Full_Adder FA_11878(s11878, c11878, in11878_1, in11878_2, s10099[0]);
    wire[0:0] s11879, in11879_1, in11879_2;
    wire c11879;
    assign in11879_1 = {c10092};
    assign in11879_2 = {c10093};
    Full_Adder FA_11879(s11879, c11879, in11879_1, in11879_2, c10091);
    wire[0:0] s11880, in11880_1, in11880_2;
    wire c11880;
    assign in11880_1 = {c10095};
    assign in11880_2 = {c10096};
    Full_Adder FA_11880(s11880, c11880, in11880_1, in11880_2, c10094);
    wire[0:0] s11881, in11881_1, in11881_2;
    wire c11881;
    assign in11881_1 = {c10098};
    assign in11881_2 = {c10099};
    Full_Adder FA_11881(s11881, c11881, in11881_1, in11881_2, c10097);
    wire[0:0] s11882, in11882_1, in11882_2;
    wire c11882;
    assign in11882_1 = {c10101};
    assign in11882_2 = {c10102};
    Full_Adder FA_11882(s11882, c11882, in11882_1, in11882_2, c10100);
    wire[0:0] s11883, in11883_1, in11883_2;
    wire c11883;
    assign in11883_1 = {s10104[0]};
    assign in11883_2 = {s10105[0]};
    Full_Adder FA_11883(s11883, c11883, in11883_1, in11883_2, c10103);
    wire[0:0] s11884, in11884_1, in11884_2;
    wire c11884;
    assign in11884_1 = {s10107[0]};
    assign in11884_2 = {s10108[0]};
    Full_Adder FA_11884(s11884, c11884, in11884_1, in11884_2, s10106[0]);
    wire[0:0] s11885, in11885_1, in11885_2;
    wire c11885;
    assign in11885_1 = {s10110[0]};
    assign in11885_2 = {s10111[0]};
    Full_Adder FA_11885(s11885, c11885, in11885_1, in11885_2, s10109[0]);
    wire[0:0] s11886, in11886_1, in11886_2;
    wire c11886;
    assign in11886_1 = {s10113[0]};
    assign in11886_2 = {s10114[0]};
    Full_Adder FA_11886(s11886, c11886, in11886_1, in11886_2, s10112[0]);
    wire[0:0] s11887, in11887_1, in11887_2;
    wire c11887;
    assign in11887_1 = {c10105};
    assign in11887_2 = {c10106};
    Full_Adder FA_11887(s11887, c11887, in11887_1, in11887_2, c10104);
    wire[0:0] s11888, in11888_1, in11888_2;
    wire c11888;
    assign in11888_1 = {c10108};
    assign in11888_2 = {c10109};
    Full_Adder FA_11888(s11888, c11888, in11888_1, in11888_2, c10107);
    wire[0:0] s11889, in11889_1, in11889_2;
    wire c11889;
    assign in11889_1 = {c10111};
    assign in11889_2 = {c10112};
    Full_Adder FA_11889(s11889, c11889, in11889_1, in11889_2, c10110);
    wire[0:0] s11890, in11890_1, in11890_2;
    wire c11890;
    assign in11890_1 = {c10114};
    assign in11890_2 = {c10115};
    Full_Adder FA_11890(s11890, c11890, in11890_1, in11890_2, c10113);
    wire[0:0] s11891, in11891_1, in11891_2;
    wire c11891;
    assign in11891_1 = {s10117[0]};
    assign in11891_2 = {s10118[0]};
    Full_Adder FA_11891(s11891, c11891, in11891_1, in11891_2, c10116);
    wire[0:0] s11892, in11892_1, in11892_2;
    wire c11892;
    assign in11892_1 = {s10120[0]};
    assign in11892_2 = {s10121[0]};
    Full_Adder FA_11892(s11892, c11892, in11892_1, in11892_2, s10119[0]);
    wire[0:0] s11893, in11893_1, in11893_2;
    wire c11893;
    assign in11893_1 = {s10123[0]};
    assign in11893_2 = {s10124[0]};
    Full_Adder FA_11893(s11893, c11893, in11893_1, in11893_2, s10122[0]);
    wire[0:0] s11894, in11894_1, in11894_2;
    wire c11894;
    assign in11894_1 = {s10126[0]};
    assign in11894_2 = {s10127[0]};
    Full_Adder FA_11894(s11894, c11894, in11894_1, in11894_2, s10125[0]);
    wire[0:0] s11895, in11895_1, in11895_2;
    wire c11895;
    assign in11895_1 = {c10118};
    assign in11895_2 = {c10119};
    Full_Adder FA_11895(s11895, c11895, in11895_1, in11895_2, c10117);
    wire[0:0] s11896, in11896_1, in11896_2;
    wire c11896;
    assign in11896_1 = {c10121};
    assign in11896_2 = {c10122};
    Full_Adder FA_11896(s11896, c11896, in11896_1, in11896_2, c10120);
    wire[0:0] s11897, in11897_1, in11897_2;
    wire c11897;
    assign in11897_1 = {c10124};
    assign in11897_2 = {c10125};
    Full_Adder FA_11897(s11897, c11897, in11897_1, in11897_2, c10123);
    wire[0:0] s11898, in11898_1, in11898_2;
    wire c11898;
    assign in11898_1 = {c10127};
    assign in11898_2 = {c10128};
    Full_Adder FA_11898(s11898, c11898, in11898_1, in11898_2, c10126);
    wire[0:0] s11899, in11899_1, in11899_2;
    wire c11899;
    assign in11899_1 = {s10130[0]};
    assign in11899_2 = {s10131[0]};
    Full_Adder FA_11899(s11899, c11899, in11899_1, in11899_2, c10129);
    wire[0:0] s11900, in11900_1, in11900_2;
    wire c11900;
    assign in11900_1 = {s10133[0]};
    assign in11900_2 = {s10134[0]};
    Full_Adder FA_11900(s11900, c11900, in11900_1, in11900_2, s10132[0]);
    wire[0:0] s11901, in11901_1, in11901_2;
    wire c11901;
    assign in11901_1 = {s10136[0]};
    assign in11901_2 = {s10137[0]};
    Full_Adder FA_11901(s11901, c11901, in11901_1, in11901_2, s10135[0]);
    wire[0:0] s11902, in11902_1, in11902_2;
    wire c11902;
    assign in11902_1 = {s10139[0]};
    assign in11902_2 = {s10140[0]};
    Full_Adder FA_11902(s11902, c11902, in11902_1, in11902_2, s10138[0]);
    wire[0:0] s11903, in11903_1, in11903_2;
    wire c11903;
    assign in11903_1 = {c10131};
    assign in11903_2 = {c10132};
    Full_Adder FA_11903(s11903, c11903, in11903_1, in11903_2, c10130);
    wire[0:0] s11904, in11904_1, in11904_2;
    wire c11904;
    assign in11904_1 = {c10134};
    assign in11904_2 = {c10135};
    Full_Adder FA_11904(s11904, c11904, in11904_1, in11904_2, c10133);
    wire[0:0] s11905, in11905_1, in11905_2;
    wire c11905;
    assign in11905_1 = {c10137};
    assign in11905_2 = {c10138};
    Full_Adder FA_11905(s11905, c11905, in11905_1, in11905_2, c10136);
    wire[0:0] s11906, in11906_1, in11906_2;
    wire c11906;
    assign in11906_1 = {c10140};
    assign in11906_2 = {c10141};
    Full_Adder FA_11906(s11906, c11906, in11906_1, in11906_2, c10139);
    wire[0:0] s11907, in11907_1, in11907_2;
    wire c11907;
    assign in11907_1 = {s10143[0]};
    assign in11907_2 = {s10144[0]};
    Full_Adder FA_11907(s11907, c11907, in11907_1, in11907_2, c10142);
    wire[0:0] s11908, in11908_1, in11908_2;
    wire c11908;
    assign in11908_1 = {s10146[0]};
    assign in11908_2 = {s10147[0]};
    Full_Adder FA_11908(s11908, c11908, in11908_1, in11908_2, s10145[0]);
    wire[0:0] s11909, in11909_1, in11909_2;
    wire c11909;
    assign in11909_1 = {s10149[0]};
    assign in11909_2 = {s10150[0]};
    Full_Adder FA_11909(s11909, c11909, in11909_1, in11909_2, s10148[0]);
    wire[0:0] s11910, in11910_1, in11910_2;
    wire c11910;
    assign in11910_1 = {s10152[0]};
    assign in11910_2 = {s10153[0]};
    Full_Adder FA_11910(s11910, c11910, in11910_1, in11910_2, s10151[0]);
    wire[0:0] s11911, in11911_1, in11911_2;
    wire c11911;
    assign in11911_1 = {c10144};
    assign in11911_2 = {c10145};
    Full_Adder FA_11911(s11911, c11911, in11911_1, in11911_2, c10143);
    wire[0:0] s11912, in11912_1, in11912_2;
    wire c11912;
    assign in11912_1 = {c10147};
    assign in11912_2 = {c10148};
    Full_Adder FA_11912(s11912, c11912, in11912_1, in11912_2, c10146);
    wire[0:0] s11913, in11913_1, in11913_2;
    wire c11913;
    assign in11913_1 = {c10150};
    assign in11913_2 = {c10151};
    Full_Adder FA_11913(s11913, c11913, in11913_1, in11913_2, c10149);
    wire[0:0] s11914, in11914_1, in11914_2;
    wire c11914;
    assign in11914_1 = {c10153};
    assign in11914_2 = {c10154};
    Full_Adder FA_11914(s11914, c11914, in11914_1, in11914_2, c10152);
    wire[0:0] s11915, in11915_1, in11915_2;
    wire c11915;
    assign in11915_1 = {s10156[0]};
    assign in11915_2 = {s10157[0]};
    Full_Adder FA_11915(s11915, c11915, in11915_1, in11915_2, c10155);
    wire[0:0] s11916, in11916_1, in11916_2;
    wire c11916;
    assign in11916_1 = {s10159[0]};
    assign in11916_2 = {s10160[0]};
    Full_Adder FA_11916(s11916, c11916, in11916_1, in11916_2, s10158[0]);
    wire[0:0] s11917, in11917_1, in11917_2;
    wire c11917;
    assign in11917_1 = {s10162[0]};
    assign in11917_2 = {s10163[0]};
    Full_Adder FA_11917(s11917, c11917, in11917_1, in11917_2, s10161[0]);
    wire[0:0] s11918, in11918_1, in11918_2;
    wire c11918;
    assign in11918_1 = {s10165[0]};
    assign in11918_2 = {s10166[0]};
    Full_Adder FA_11918(s11918, c11918, in11918_1, in11918_2, s10164[0]);
    wire[0:0] s11919, in11919_1, in11919_2;
    wire c11919;
    assign in11919_1 = {c10157};
    assign in11919_2 = {c10158};
    Full_Adder FA_11919(s11919, c11919, in11919_1, in11919_2, c10156);
    wire[0:0] s11920, in11920_1, in11920_2;
    wire c11920;
    assign in11920_1 = {c10160};
    assign in11920_2 = {c10161};
    Full_Adder FA_11920(s11920, c11920, in11920_1, in11920_2, c10159);
    wire[0:0] s11921, in11921_1, in11921_2;
    wire c11921;
    assign in11921_1 = {c10163};
    assign in11921_2 = {c10164};
    Full_Adder FA_11921(s11921, c11921, in11921_1, in11921_2, c10162);
    wire[0:0] s11922, in11922_1, in11922_2;
    wire c11922;
    assign in11922_1 = {c10166};
    assign in11922_2 = {c10167};
    Full_Adder FA_11922(s11922, c11922, in11922_1, in11922_2, c10165);
    wire[0:0] s11923, in11923_1, in11923_2;
    wire c11923;
    assign in11923_1 = {s10169[0]};
    assign in11923_2 = {s10170[0]};
    Full_Adder FA_11923(s11923, c11923, in11923_1, in11923_2, c10168);
    wire[0:0] s11924, in11924_1, in11924_2;
    wire c11924;
    assign in11924_1 = {s10172[0]};
    assign in11924_2 = {s10173[0]};
    Full_Adder FA_11924(s11924, c11924, in11924_1, in11924_2, s10171[0]);
    wire[0:0] s11925, in11925_1, in11925_2;
    wire c11925;
    assign in11925_1 = {s10175[0]};
    assign in11925_2 = {s10176[0]};
    Full_Adder FA_11925(s11925, c11925, in11925_1, in11925_2, s10174[0]);
    wire[0:0] s11926, in11926_1, in11926_2;
    wire c11926;
    assign in11926_1 = {s10178[0]};
    assign in11926_2 = {s10179[0]};
    Full_Adder FA_11926(s11926, c11926, in11926_1, in11926_2, s10177[0]);
    wire[0:0] s11927, in11927_1, in11927_2;
    wire c11927;
    assign in11927_1 = {c10170};
    assign in11927_2 = {c10171};
    Full_Adder FA_11927(s11927, c11927, in11927_1, in11927_2, c10169);
    wire[0:0] s11928, in11928_1, in11928_2;
    wire c11928;
    assign in11928_1 = {c10173};
    assign in11928_2 = {c10174};
    Full_Adder FA_11928(s11928, c11928, in11928_1, in11928_2, c10172);
    wire[0:0] s11929, in11929_1, in11929_2;
    wire c11929;
    assign in11929_1 = {c10176};
    assign in11929_2 = {c10177};
    Full_Adder FA_11929(s11929, c11929, in11929_1, in11929_2, c10175);
    wire[0:0] s11930, in11930_1, in11930_2;
    wire c11930;
    assign in11930_1 = {c10179};
    assign in11930_2 = {c10180};
    Full_Adder FA_11930(s11930, c11930, in11930_1, in11930_2, c10178);
    wire[0:0] s11931, in11931_1, in11931_2;
    wire c11931;
    assign in11931_1 = {s10182[0]};
    assign in11931_2 = {s10183[0]};
    Full_Adder FA_11931(s11931, c11931, in11931_1, in11931_2, c10181);
    wire[0:0] s11932, in11932_1, in11932_2;
    wire c11932;
    assign in11932_1 = {s10185[0]};
    assign in11932_2 = {s10186[0]};
    Full_Adder FA_11932(s11932, c11932, in11932_1, in11932_2, s10184[0]);
    wire[0:0] s11933, in11933_1, in11933_2;
    wire c11933;
    assign in11933_1 = {s10188[0]};
    assign in11933_2 = {s10189[0]};
    Full_Adder FA_11933(s11933, c11933, in11933_1, in11933_2, s10187[0]);
    wire[0:0] s11934, in11934_1, in11934_2;
    wire c11934;
    assign in11934_1 = {s10191[0]};
    assign in11934_2 = {s10192[0]};
    Full_Adder FA_11934(s11934, c11934, in11934_1, in11934_2, s10190[0]);
    wire[0:0] s11935, in11935_1, in11935_2;
    wire c11935;
    assign in11935_1 = {c10183};
    assign in11935_2 = {c10184};
    Full_Adder FA_11935(s11935, c11935, in11935_1, in11935_2, c10182);
    wire[0:0] s11936, in11936_1, in11936_2;
    wire c11936;
    assign in11936_1 = {c10186};
    assign in11936_2 = {c10187};
    Full_Adder FA_11936(s11936, c11936, in11936_1, in11936_2, c10185);
    wire[0:0] s11937, in11937_1, in11937_2;
    wire c11937;
    assign in11937_1 = {c10189};
    assign in11937_2 = {c10190};
    Full_Adder FA_11937(s11937, c11937, in11937_1, in11937_2, c10188);
    wire[0:0] s11938, in11938_1, in11938_2;
    wire c11938;
    assign in11938_1 = {c10192};
    assign in11938_2 = {c10193};
    Full_Adder FA_11938(s11938, c11938, in11938_1, in11938_2, c10191);
    wire[0:0] s11939, in11939_1, in11939_2;
    wire c11939;
    assign in11939_1 = {s10195[0]};
    assign in11939_2 = {s10196[0]};
    Full_Adder FA_11939(s11939, c11939, in11939_1, in11939_2, c10194);
    wire[0:0] s11940, in11940_1, in11940_2;
    wire c11940;
    assign in11940_1 = {s10198[0]};
    assign in11940_2 = {s10199[0]};
    Full_Adder FA_11940(s11940, c11940, in11940_1, in11940_2, s10197[0]);
    wire[0:0] s11941, in11941_1, in11941_2;
    wire c11941;
    assign in11941_1 = {s10201[0]};
    assign in11941_2 = {s10202[0]};
    Full_Adder FA_11941(s11941, c11941, in11941_1, in11941_2, s10200[0]);
    wire[0:0] s11942, in11942_1, in11942_2;
    wire c11942;
    assign in11942_1 = {s10204[0]};
    assign in11942_2 = {s10205[0]};
    Full_Adder FA_11942(s11942, c11942, in11942_1, in11942_2, s10203[0]);
    wire[0:0] s11943, in11943_1, in11943_2;
    wire c11943;
    assign in11943_1 = {c10196};
    assign in11943_2 = {c10197};
    Full_Adder FA_11943(s11943, c11943, in11943_1, in11943_2, c10195);
    wire[0:0] s11944, in11944_1, in11944_2;
    wire c11944;
    assign in11944_1 = {c10199};
    assign in11944_2 = {c10200};
    Full_Adder FA_11944(s11944, c11944, in11944_1, in11944_2, c10198);
    wire[0:0] s11945, in11945_1, in11945_2;
    wire c11945;
    assign in11945_1 = {c10202};
    assign in11945_2 = {c10203};
    Full_Adder FA_11945(s11945, c11945, in11945_1, in11945_2, c10201);
    wire[0:0] s11946, in11946_1, in11946_2;
    wire c11946;
    assign in11946_1 = {c10205};
    assign in11946_2 = {c10206};
    Full_Adder FA_11946(s11946, c11946, in11946_1, in11946_2, c10204);
    wire[0:0] s11947, in11947_1, in11947_2;
    wire c11947;
    assign in11947_1 = {s10208[0]};
    assign in11947_2 = {s10209[0]};
    Full_Adder FA_11947(s11947, c11947, in11947_1, in11947_2, c10207);
    wire[0:0] s11948, in11948_1, in11948_2;
    wire c11948;
    assign in11948_1 = {s10211[0]};
    assign in11948_2 = {s10212[0]};
    Full_Adder FA_11948(s11948, c11948, in11948_1, in11948_2, s10210[0]);
    wire[0:0] s11949, in11949_1, in11949_2;
    wire c11949;
    assign in11949_1 = {s10214[0]};
    assign in11949_2 = {s10215[0]};
    Full_Adder FA_11949(s11949, c11949, in11949_1, in11949_2, s10213[0]);
    wire[0:0] s11950, in11950_1, in11950_2;
    wire c11950;
    assign in11950_1 = {s10217[0]};
    assign in11950_2 = {s10218[0]};
    Full_Adder FA_11950(s11950, c11950, in11950_1, in11950_2, s10216[0]);
    wire[0:0] s11951, in11951_1, in11951_2;
    wire c11951;
    assign in11951_1 = {c10209};
    assign in11951_2 = {c10210};
    Full_Adder FA_11951(s11951, c11951, in11951_1, in11951_2, c10208);
    wire[0:0] s11952, in11952_1, in11952_2;
    wire c11952;
    assign in11952_1 = {c10212};
    assign in11952_2 = {c10213};
    Full_Adder FA_11952(s11952, c11952, in11952_1, in11952_2, c10211);
    wire[0:0] s11953, in11953_1, in11953_2;
    wire c11953;
    assign in11953_1 = {c10215};
    assign in11953_2 = {c10216};
    Full_Adder FA_11953(s11953, c11953, in11953_1, in11953_2, c10214);
    wire[0:0] s11954, in11954_1, in11954_2;
    wire c11954;
    assign in11954_1 = {c10218};
    assign in11954_2 = {c10219};
    Full_Adder FA_11954(s11954, c11954, in11954_1, in11954_2, c10217);
    wire[0:0] s11955, in11955_1, in11955_2;
    wire c11955;
    assign in11955_1 = {s10221[0]};
    assign in11955_2 = {s10222[0]};
    Full_Adder FA_11955(s11955, c11955, in11955_1, in11955_2, c10220);
    wire[0:0] s11956, in11956_1, in11956_2;
    wire c11956;
    assign in11956_1 = {s10224[0]};
    assign in11956_2 = {s10225[0]};
    Full_Adder FA_11956(s11956, c11956, in11956_1, in11956_2, s10223[0]);
    wire[0:0] s11957, in11957_1, in11957_2;
    wire c11957;
    assign in11957_1 = {s10227[0]};
    assign in11957_2 = {s10228[0]};
    Full_Adder FA_11957(s11957, c11957, in11957_1, in11957_2, s10226[0]);
    wire[0:0] s11958, in11958_1, in11958_2;
    wire c11958;
    assign in11958_1 = {s10230[0]};
    assign in11958_2 = {s10231[0]};
    Full_Adder FA_11958(s11958, c11958, in11958_1, in11958_2, s10229[0]);
    wire[0:0] s11959, in11959_1, in11959_2;
    wire c11959;
    assign in11959_1 = {c10222};
    assign in11959_2 = {c10223};
    Full_Adder FA_11959(s11959, c11959, in11959_1, in11959_2, c10221);
    wire[0:0] s11960, in11960_1, in11960_2;
    wire c11960;
    assign in11960_1 = {c10225};
    assign in11960_2 = {c10226};
    Full_Adder FA_11960(s11960, c11960, in11960_1, in11960_2, c10224);
    wire[0:0] s11961, in11961_1, in11961_2;
    wire c11961;
    assign in11961_1 = {c10228};
    assign in11961_2 = {c10229};
    Full_Adder FA_11961(s11961, c11961, in11961_1, in11961_2, c10227);
    wire[0:0] s11962, in11962_1, in11962_2;
    wire c11962;
    assign in11962_1 = {c10231};
    assign in11962_2 = {c10232};
    Full_Adder FA_11962(s11962, c11962, in11962_1, in11962_2, c10230);
    wire[0:0] s11963, in11963_1, in11963_2;
    wire c11963;
    assign in11963_1 = {s10234[0]};
    assign in11963_2 = {s10235[0]};
    Full_Adder FA_11963(s11963, c11963, in11963_1, in11963_2, c10233);
    wire[0:0] s11964, in11964_1, in11964_2;
    wire c11964;
    assign in11964_1 = {s10237[0]};
    assign in11964_2 = {s10238[0]};
    Full_Adder FA_11964(s11964, c11964, in11964_1, in11964_2, s10236[0]);
    wire[0:0] s11965, in11965_1, in11965_2;
    wire c11965;
    assign in11965_1 = {s10240[0]};
    assign in11965_2 = {s10241[0]};
    Full_Adder FA_11965(s11965, c11965, in11965_1, in11965_2, s10239[0]);
    wire[0:0] s11966, in11966_1, in11966_2;
    wire c11966;
    assign in11966_1 = {s10243[0]};
    assign in11966_2 = {s10244[0]};
    Full_Adder FA_11966(s11966, c11966, in11966_1, in11966_2, s10242[0]);
    wire[0:0] s11967, in11967_1, in11967_2;
    wire c11967;
    assign in11967_1 = {c10235};
    assign in11967_2 = {c10236};
    Full_Adder FA_11967(s11967, c11967, in11967_1, in11967_2, c10234);
    wire[0:0] s11968, in11968_1, in11968_2;
    wire c11968;
    assign in11968_1 = {c10238};
    assign in11968_2 = {c10239};
    Full_Adder FA_11968(s11968, c11968, in11968_1, in11968_2, c10237);
    wire[0:0] s11969, in11969_1, in11969_2;
    wire c11969;
    assign in11969_1 = {c10241};
    assign in11969_2 = {c10242};
    Full_Adder FA_11969(s11969, c11969, in11969_1, in11969_2, c10240);
    wire[0:0] s11970, in11970_1, in11970_2;
    wire c11970;
    assign in11970_1 = {c10244};
    assign in11970_2 = {c10245};
    Full_Adder FA_11970(s11970, c11970, in11970_1, in11970_2, c10243);
    wire[0:0] s11971, in11971_1, in11971_2;
    wire c11971;
    assign in11971_1 = {s10247[0]};
    assign in11971_2 = {s10248[0]};
    Full_Adder FA_11971(s11971, c11971, in11971_1, in11971_2, c10246);
    wire[0:0] s11972, in11972_1, in11972_2;
    wire c11972;
    assign in11972_1 = {s10250[0]};
    assign in11972_2 = {s10251[0]};
    Full_Adder FA_11972(s11972, c11972, in11972_1, in11972_2, s10249[0]);
    wire[0:0] s11973, in11973_1, in11973_2;
    wire c11973;
    assign in11973_1 = {s10253[0]};
    assign in11973_2 = {s10254[0]};
    Full_Adder FA_11973(s11973, c11973, in11973_1, in11973_2, s10252[0]);
    wire[0:0] s11974, in11974_1, in11974_2;
    wire c11974;
    assign in11974_1 = {s10256[0]};
    assign in11974_2 = {s10257[0]};
    Full_Adder FA_11974(s11974, c11974, in11974_1, in11974_2, s10255[0]);
    wire[0:0] s11975, in11975_1, in11975_2;
    wire c11975;
    assign in11975_1 = {c10248};
    assign in11975_2 = {c10249};
    Full_Adder FA_11975(s11975, c11975, in11975_1, in11975_2, c10247);
    wire[0:0] s11976, in11976_1, in11976_2;
    wire c11976;
    assign in11976_1 = {c10251};
    assign in11976_2 = {c10252};
    Full_Adder FA_11976(s11976, c11976, in11976_1, in11976_2, c10250);
    wire[0:0] s11977, in11977_1, in11977_2;
    wire c11977;
    assign in11977_1 = {c10254};
    assign in11977_2 = {c10255};
    Full_Adder FA_11977(s11977, c11977, in11977_1, in11977_2, c10253);
    wire[0:0] s11978, in11978_1, in11978_2;
    wire c11978;
    assign in11978_1 = {c10257};
    assign in11978_2 = {c10258};
    Full_Adder FA_11978(s11978, c11978, in11978_1, in11978_2, c10256);
    wire[0:0] s11979, in11979_1, in11979_2;
    wire c11979;
    assign in11979_1 = {s10260[0]};
    assign in11979_2 = {s10261[0]};
    Full_Adder FA_11979(s11979, c11979, in11979_1, in11979_2, c10259);
    wire[0:0] s11980, in11980_1, in11980_2;
    wire c11980;
    assign in11980_1 = {s10263[0]};
    assign in11980_2 = {s10264[0]};
    Full_Adder FA_11980(s11980, c11980, in11980_1, in11980_2, s10262[0]);
    wire[0:0] s11981, in11981_1, in11981_2;
    wire c11981;
    assign in11981_1 = {s10266[0]};
    assign in11981_2 = {s10267[0]};
    Full_Adder FA_11981(s11981, c11981, in11981_1, in11981_2, s10265[0]);
    wire[0:0] s11982, in11982_1, in11982_2;
    wire c11982;
    assign in11982_1 = {s10269[0]};
    assign in11982_2 = {s10270[0]};
    Full_Adder FA_11982(s11982, c11982, in11982_1, in11982_2, s10268[0]);
    wire[0:0] s11983, in11983_1, in11983_2;
    wire c11983;
    assign in11983_1 = {c10261};
    assign in11983_2 = {c10262};
    Full_Adder FA_11983(s11983, c11983, in11983_1, in11983_2, c10260);
    wire[0:0] s11984, in11984_1, in11984_2;
    wire c11984;
    assign in11984_1 = {c10264};
    assign in11984_2 = {c10265};
    Full_Adder FA_11984(s11984, c11984, in11984_1, in11984_2, c10263);
    wire[0:0] s11985, in11985_1, in11985_2;
    wire c11985;
    assign in11985_1 = {c10267};
    assign in11985_2 = {c10268};
    Full_Adder FA_11985(s11985, c11985, in11985_1, in11985_2, c10266);
    wire[0:0] s11986, in11986_1, in11986_2;
    wire c11986;
    assign in11986_1 = {c10270};
    assign in11986_2 = {c10271};
    Full_Adder FA_11986(s11986, c11986, in11986_1, in11986_2, c10269);
    wire[0:0] s11987, in11987_1, in11987_2;
    wire c11987;
    assign in11987_1 = {s10273[0]};
    assign in11987_2 = {s10274[0]};
    Full_Adder FA_11987(s11987, c11987, in11987_1, in11987_2, c10272);
    wire[0:0] s11988, in11988_1, in11988_2;
    wire c11988;
    assign in11988_1 = {s10276[0]};
    assign in11988_2 = {s10277[0]};
    Full_Adder FA_11988(s11988, c11988, in11988_1, in11988_2, s10275[0]);
    wire[0:0] s11989, in11989_1, in11989_2;
    wire c11989;
    assign in11989_1 = {s10279[0]};
    assign in11989_2 = {s10280[0]};
    Full_Adder FA_11989(s11989, c11989, in11989_1, in11989_2, s10278[0]);
    wire[0:0] s11990, in11990_1, in11990_2;
    wire c11990;
    assign in11990_1 = {s10282[0]};
    assign in11990_2 = {s10283[0]};
    Full_Adder FA_11990(s11990, c11990, in11990_1, in11990_2, s10281[0]);
    wire[0:0] s11991, in11991_1, in11991_2;
    wire c11991;
    assign in11991_1 = {c10274};
    assign in11991_2 = {c10275};
    Full_Adder FA_11991(s11991, c11991, in11991_1, in11991_2, c10273);
    wire[0:0] s11992, in11992_1, in11992_2;
    wire c11992;
    assign in11992_1 = {c10277};
    assign in11992_2 = {c10278};
    Full_Adder FA_11992(s11992, c11992, in11992_1, in11992_2, c10276);
    wire[0:0] s11993, in11993_1, in11993_2;
    wire c11993;
    assign in11993_1 = {c10280};
    assign in11993_2 = {c10281};
    Full_Adder FA_11993(s11993, c11993, in11993_1, in11993_2, c10279);
    wire[0:0] s11994, in11994_1, in11994_2;
    wire c11994;
    assign in11994_1 = {c10283};
    assign in11994_2 = {c10284};
    Full_Adder FA_11994(s11994, c11994, in11994_1, in11994_2, c10282);
    wire[0:0] s11995, in11995_1, in11995_2;
    wire c11995;
    assign in11995_1 = {s10286[0]};
    assign in11995_2 = {s10287[0]};
    Full_Adder FA_11995(s11995, c11995, in11995_1, in11995_2, c10285);
    wire[0:0] s11996, in11996_1, in11996_2;
    wire c11996;
    assign in11996_1 = {s10289[0]};
    assign in11996_2 = {s10290[0]};
    Full_Adder FA_11996(s11996, c11996, in11996_1, in11996_2, s10288[0]);
    wire[0:0] s11997, in11997_1, in11997_2;
    wire c11997;
    assign in11997_1 = {s10292[0]};
    assign in11997_2 = {s10293[0]};
    Full_Adder FA_11997(s11997, c11997, in11997_1, in11997_2, s10291[0]);
    wire[0:0] s11998, in11998_1, in11998_2;
    wire c11998;
    assign in11998_1 = {s10295[0]};
    assign in11998_2 = {s10296[0]};
    Full_Adder FA_11998(s11998, c11998, in11998_1, in11998_2, s10294[0]);
    wire[0:0] s11999, in11999_1, in11999_2;
    wire c11999;
    assign in11999_1 = {c10287};
    assign in11999_2 = {c10288};
    Full_Adder FA_11999(s11999, c11999, in11999_1, in11999_2, c10286);
    wire[0:0] s12000, in12000_1, in12000_2;
    wire c12000;
    assign in12000_1 = {c10290};
    assign in12000_2 = {c10291};
    Full_Adder FA_12000(s12000, c12000, in12000_1, in12000_2, c10289);
    wire[0:0] s12001, in12001_1, in12001_2;
    wire c12001;
    assign in12001_1 = {c10293};
    assign in12001_2 = {c10294};
    Full_Adder FA_12001(s12001, c12001, in12001_1, in12001_2, c10292);
    wire[0:0] s12002, in12002_1, in12002_2;
    wire c12002;
    assign in12002_1 = {c10296};
    assign in12002_2 = {c10297};
    Full_Adder FA_12002(s12002, c12002, in12002_1, in12002_2, c10295);
    wire[0:0] s12003, in12003_1, in12003_2;
    wire c12003;
    assign in12003_1 = {s10299[0]};
    assign in12003_2 = {s10300[0]};
    Full_Adder FA_12003(s12003, c12003, in12003_1, in12003_2, c10298);
    wire[0:0] s12004, in12004_1, in12004_2;
    wire c12004;
    assign in12004_1 = {s10302[0]};
    assign in12004_2 = {s10303[0]};
    Full_Adder FA_12004(s12004, c12004, in12004_1, in12004_2, s10301[0]);
    wire[0:0] s12005, in12005_1, in12005_2;
    wire c12005;
    assign in12005_1 = {s10305[0]};
    assign in12005_2 = {s10306[0]};
    Full_Adder FA_12005(s12005, c12005, in12005_1, in12005_2, s10304[0]);
    wire[0:0] s12006, in12006_1, in12006_2;
    wire c12006;
    assign in12006_1 = {s10308[0]};
    assign in12006_2 = {s10309[0]};
    Full_Adder FA_12006(s12006, c12006, in12006_1, in12006_2, s10307[0]);
    wire[0:0] s12007, in12007_1, in12007_2;
    wire c12007;
    assign in12007_1 = {c10300};
    assign in12007_2 = {c10301};
    Full_Adder FA_12007(s12007, c12007, in12007_1, in12007_2, c10299);
    wire[0:0] s12008, in12008_1, in12008_2;
    wire c12008;
    assign in12008_1 = {c10303};
    assign in12008_2 = {c10304};
    Full_Adder FA_12008(s12008, c12008, in12008_1, in12008_2, c10302);
    wire[0:0] s12009, in12009_1, in12009_2;
    wire c12009;
    assign in12009_1 = {c10306};
    assign in12009_2 = {c10307};
    Full_Adder FA_12009(s12009, c12009, in12009_1, in12009_2, c10305);
    wire[0:0] s12010, in12010_1, in12010_2;
    wire c12010;
    assign in12010_1 = {c10309};
    assign in12010_2 = {c10310};
    Full_Adder FA_12010(s12010, c12010, in12010_1, in12010_2, c10308);
    wire[0:0] s12011, in12011_1, in12011_2;
    wire c12011;
    assign in12011_1 = {s10312[0]};
    assign in12011_2 = {s10313[0]};
    Full_Adder FA_12011(s12011, c12011, in12011_1, in12011_2, c10311);
    wire[0:0] s12012, in12012_1, in12012_2;
    wire c12012;
    assign in12012_1 = {s10315[0]};
    assign in12012_2 = {s10316[0]};
    Full_Adder FA_12012(s12012, c12012, in12012_1, in12012_2, s10314[0]);
    wire[0:0] s12013, in12013_1, in12013_2;
    wire c12013;
    assign in12013_1 = {s10318[0]};
    assign in12013_2 = {s10319[0]};
    Full_Adder FA_12013(s12013, c12013, in12013_1, in12013_2, s10317[0]);
    wire[0:0] s12014, in12014_1, in12014_2;
    wire c12014;
    assign in12014_1 = {s10321[0]};
    assign in12014_2 = {s10322[0]};
    Full_Adder FA_12014(s12014, c12014, in12014_1, in12014_2, s10320[0]);
    wire[0:0] s12015, in12015_1, in12015_2;
    wire c12015;
    assign in12015_1 = {c10313};
    assign in12015_2 = {c10314};
    Full_Adder FA_12015(s12015, c12015, in12015_1, in12015_2, c10312);
    wire[0:0] s12016, in12016_1, in12016_2;
    wire c12016;
    assign in12016_1 = {c10316};
    assign in12016_2 = {c10317};
    Full_Adder FA_12016(s12016, c12016, in12016_1, in12016_2, c10315);
    wire[0:0] s12017, in12017_1, in12017_2;
    wire c12017;
    assign in12017_1 = {c10319};
    assign in12017_2 = {c10320};
    Full_Adder FA_12017(s12017, c12017, in12017_1, in12017_2, c10318);
    wire[0:0] s12018, in12018_1, in12018_2;
    wire c12018;
    assign in12018_1 = {c10322};
    assign in12018_2 = {c10323};
    Full_Adder FA_12018(s12018, c12018, in12018_1, in12018_2, c10321);
    wire[0:0] s12019, in12019_1, in12019_2;
    wire c12019;
    assign in12019_1 = {s10325[0]};
    assign in12019_2 = {s10326[0]};
    Full_Adder FA_12019(s12019, c12019, in12019_1, in12019_2, c10324);
    wire[0:0] s12020, in12020_1, in12020_2;
    wire c12020;
    assign in12020_1 = {s10328[0]};
    assign in12020_2 = {s10329[0]};
    Full_Adder FA_12020(s12020, c12020, in12020_1, in12020_2, s10327[0]);
    wire[0:0] s12021, in12021_1, in12021_2;
    wire c12021;
    assign in12021_1 = {s10331[0]};
    assign in12021_2 = {s10332[0]};
    Full_Adder FA_12021(s12021, c12021, in12021_1, in12021_2, s10330[0]);
    wire[0:0] s12022, in12022_1, in12022_2;
    wire c12022;
    assign in12022_1 = {s10334[0]};
    assign in12022_2 = {s10335[0]};
    Full_Adder FA_12022(s12022, c12022, in12022_1, in12022_2, s10333[0]);
    wire[0:0] s12023, in12023_1, in12023_2;
    wire c12023;
    assign in12023_1 = {c10326};
    assign in12023_2 = {c10327};
    Full_Adder FA_12023(s12023, c12023, in12023_1, in12023_2, c10325);
    wire[0:0] s12024, in12024_1, in12024_2;
    wire c12024;
    assign in12024_1 = {c10329};
    assign in12024_2 = {c10330};
    Full_Adder FA_12024(s12024, c12024, in12024_1, in12024_2, c10328);
    wire[0:0] s12025, in12025_1, in12025_2;
    wire c12025;
    assign in12025_1 = {c10332};
    assign in12025_2 = {c10333};
    Full_Adder FA_12025(s12025, c12025, in12025_1, in12025_2, c10331);
    wire[0:0] s12026, in12026_1, in12026_2;
    wire c12026;
    assign in12026_1 = {c10335};
    assign in12026_2 = {c10336};
    Full_Adder FA_12026(s12026, c12026, in12026_1, in12026_2, c10334);
    wire[0:0] s12027, in12027_1, in12027_2;
    wire c12027;
    assign in12027_1 = {s10338[0]};
    assign in12027_2 = {s10339[0]};
    Full_Adder FA_12027(s12027, c12027, in12027_1, in12027_2, c10337);
    wire[0:0] s12028, in12028_1, in12028_2;
    wire c12028;
    assign in12028_1 = {s10341[0]};
    assign in12028_2 = {s10342[0]};
    Full_Adder FA_12028(s12028, c12028, in12028_1, in12028_2, s10340[0]);
    wire[0:0] s12029, in12029_1, in12029_2;
    wire c12029;
    assign in12029_1 = {s10344[0]};
    assign in12029_2 = {s10345[0]};
    Full_Adder FA_12029(s12029, c12029, in12029_1, in12029_2, s10343[0]);
    wire[0:0] s12030, in12030_1, in12030_2;
    wire c12030;
    assign in12030_1 = {s10347[0]};
    assign in12030_2 = {s10348[0]};
    Full_Adder FA_12030(s12030, c12030, in12030_1, in12030_2, s10346[0]);
    wire[0:0] s12031, in12031_1, in12031_2;
    wire c12031;
    assign in12031_1 = {c10339};
    assign in12031_2 = {c10340};
    Full_Adder FA_12031(s12031, c12031, in12031_1, in12031_2, c10338);
    wire[0:0] s12032, in12032_1, in12032_2;
    wire c12032;
    assign in12032_1 = {c10342};
    assign in12032_2 = {c10343};
    Full_Adder FA_12032(s12032, c12032, in12032_1, in12032_2, c10341);
    wire[0:0] s12033, in12033_1, in12033_2;
    wire c12033;
    assign in12033_1 = {c10345};
    assign in12033_2 = {c10346};
    Full_Adder FA_12033(s12033, c12033, in12033_1, in12033_2, c10344);
    wire[0:0] s12034, in12034_1, in12034_2;
    wire c12034;
    assign in12034_1 = {c10348};
    assign in12034_2 = {c10349};
    Full_Adder FA_12034(s12034, c12034, in12034_1, in12034_2, c10347);
    wire[0:0] s12035, in12035_1, in12035_2;
    wire c12035;
    assign in12035_1 = {s10351[0]};
    assign in12035_2 = {s10352[0]};
    Full_Adder FA_12035(s12035, c12035, in12035_1, in12035_2, c10350);
    wire[0:0] s12036, in12036_1, in12036_2;
    wire c12036;
    assign in12036_1 = {s10354[0]};
    assign in12036_2 = {s10355[0]};
    Full_Adder FA_12036(s12036, c12036, in12036_1, in12036_2, s10353[0]);
    wire[0:0] s12037, in12037_1, in12037_2;
    wire c12037;
    assign in12037_1 = {s10357[0]};
    assign in12037_2 = {s10358[0]};
    Full_Adder FA_12037(s12037, c12037, in12037_1, in12037_2, s10356[0]);
    wire[0:0] s12038, in12038_1, in12038_2;
    wire c12038;
    assign in12038_1 = {s10360[0]};
    assign in12038_2 = {s10361[0]};
    Full_Adder FA_12038(s12038, c12038, in12038_1, in12038_2, s10359[0]);
    wire[0:0] s12039, in12039_1, in12039_2;
    wire c12039;
    assign in12039_1 = {c10352};
    assign in12039_2 = {c10353};
    Full_Adder FA_12039(s12039, c12039, in12039_1, in12039_2, c10351);
    wire[0:0] s12040, in12040_1, in12040_2;
    wire c12040;
    assign in12040_1 = {c10355};
    assign in12040_2 = {c10356};
    Full_Adder FA_12040(s12040, c12040, in12040_1, in12040_2, c10354);
    wire[0:0] s12041, in12041_1, in12041_2;
    wire c12041;
    assign in12041_1 = {c10358};
    assign in12041_2 = {c10359};
    Full_Adder FA_12041(s12041, c12041, in12041_1, in12041_2, c10357);
    wire[0:0] s12042, in12042_1, in12042_2;
    wire c12042;
    assign in12042_1 = {c10361};
    assign in12042_2 = {c10362};
    Full_Adder FA_12042(s12042, c12042, in12042_1, in12042_2, c10360);
    wire[0:0] s12043, in12043_1, in12043_2;
    wire c12043;
    assign in12043_1 = {s10364[0]};
    assign in12043_2 = {s10365[0]};
    Full_Adder FA_12043(s12043, c12043, in12043_1, in12043_2, c10363);
    wire[0:0] s12044, in12044_1, in12044_2;
    wire c12044;
    assign in12044_1 = {s10367[0]};
    assign in12044_2 = {s10368[0]};
    Full_Adder FA_12044(s12044, c12044, in12044_1, in12044_2, s10366[0]);
    wire[0:0] s12045, in12045_1, in12045_2;
    wire c12045;
    assign in12045_1 = {s10370[0]};
    assign in12045_2 = {s10371[0]};
    Full_Adder FA_12045(s12045, c12045, in12045_1, in12045_2, s10369[0]);
    wire[0:0] s12046, in12046_1, in12046_2;
    wire c12046;
    assign in12046_1 = {s10373[0]};
    assign in12046_2 = {s10374[0]};
    Full_Adder FA_12046(s12046, c12046, in12046_1, in12046_2, s10372[0]);
    wire[0:0] s12047, in12047_1, in12047_2;
    wire c12047;
    assign in12047_1 = {c10365};
    assign in12047_2 = {c10366};
    Full_Adder FA_12047(s12047, c12047, in12047_1, in12047_2, c10364);
    wire[0:0] s12048, in12048_1, in12048_2;
    wire c12048;
    assign in12048_1 = {c10368};
    assign in12048_2 = {c10369};
    Full_Adder FA_12048(s12048, c12048, in12048_1, in12048_2, c10367);
    wire[0:0] s12049, in12049_1, in12049_2;
    wire c12049;
    assign in12049_1 = {c10371};
    assign in12049_2 = {c10372};
    Full_Adder FA_12049(s12049, c12049, in12049_1, in12049_2, c10370);
    wire[0:0] s12050, in12050_1, in12050_2;
    wire c12050;
    assign in12050_1 = {c10374};
    assign in12050_2 = {c10375};
    Full_Adder FA_12050(s12050, c12050, in12050_1, in12050_2, c10373);
    wire[0:0] s12051, in12051_1, in12051_2;
    wire c12051;
    assign in12051_1 = {s10377[0]};
    assign in12051_2 = {s10378[0]};
    Full_Adder FA_12051(s12051, c12051, in12051_1, in12051_2, c10376);
    wire[0:0] s12052, in12052_1, in12052_2;
    wire c12052;
    assign in12052_1 = {s10380[0]};
    assign in12052_2 = {s10381[0]};
    Full_Adder FA_12052(s12052, c12052, in12052_1, in12052_2, s10379[0]);
    wire[0:0] s12053, in12053_1, in12053_2;
    wire c12053;
    assign in12053_1 = {s10383[0]};
    assign in12053_2 = {s10384[0]};
    Full_Adder FA_12053(s12053, c12053, in12053_1, in12053_2, s10382[0]);
    wire[0:0] s12054, in12054_1, in12054_2;
    wire c12054;
    assign in12054_1 = {s10386[0]};
    assign in12054_2 = {s10387[0]};
    Full_Adder FA_12054(s12054, c12054, in12054_1, in12054_2, s10385[0]);
    wire[0:0] s12055, in12055_1, in12055_2;
    wire c12055;
    assign in12055_1 = {c10378};
    assign in12055_2 = {c10379};
    Full_Adder FA_12055(s12055, c12055, in12055_1, in12055_2, c10377);
    wire[0:0] s12056, in12056_1, in12056_2;
    wire c12056;
    assign in12056_1 = {c10381};
    assign in12056_2 = {c10382};
    Full_Adder FA_12056(s12056, c12056, in12056_1, in12056_2, c10380);
    wire[0:0] s12057, in12057_1, in12057_2;
    wire c12057;
    assign in12057_1 = {c10384};
    assign in12057_2 = {c10385};
    Full_Adder FA_12057(s12057, c12057, in12057_1, in12057_2, c10383);
    wire[0:0] s12058, in12058_1, in12058_2;
    wire c12058;
    assign in12058_1 = {c10387};
    assign in12058_2 = {c10388};
    Full_Adder FA_12058(s12058, c12058, in12058_1, in12058_2, c10386);
    wire[0:0] s12059, in12059_1, in12059_2;
    wire c12059;
    assign in12059_1 = {s10390[0]};
    assign in12059_2 = {s10391[0]};
    Full_Adder FA_12059(s12059, c12059, in12059_1, in12059_2, c10389);
    wire[0:0] s12060, in12060_1, in12060_2;
    wire c12060;
    assign in12060_1 = {s10393[0]};
    assign in12060_2 = {s10394[0]};
    Full_Adder FA_12060(s12060, c12060, in12060_1, in12060_2, s10392[0]);
    wire[0:0] s12061, in12061_1, in12061_2;
    wire c12061;
    assign in12061_1 = {s10396[0]};
    assign in12061_2 = {s10397[0]};
    Full_Adder FA_12061(s12061, c12061, in12061_1, in12061_2, s10395[0]);
    wire[0:0] s12062, in12062_1, in12062_2;
    wire c12062;
    assign in12062_1 = {s10399[0]};
    assign in12062_2 = {s10400[0]};
    Full_Adder FA_12062(s12062, c12062, in12062_1, in12062_2, s10398[0]);
    wire[0:0] s12063, in12063_1, in12063_2;
    wire c12063;
    assign in12063_1 = {c10391};
    assign in12063_2 = {c10392};
    Full_Adder FA_12063(s12063, c12063, in12063_1, in12063_2, c10390);
    wire[0:0] s12064, in12064_1, in12064_2;
    wire c12064;
    assign in12064_1 = {c10394};
    assign in12064_2 = {c10395};
    Full_Adder FA_12064(s12064, c12064, in12064_1, in12064_2, c10393);
    wire[0:0] s12065, in12065_1, in12065_2;
    wire c12065;
    assign in12065_1 = {c10397};
    assign in12065_2 = {c10398};
    Full_Adder FA_12065(s12065, c12065, in12065_1, in12065_2, c10396);
    wire[0:0] s12066, in12066_1, in12066_2;
    wire c12066;
    assign in12066_1 = {c10400};
    assign in12066_2 = {c10401};
    Full_Adder FA_12066(s12066, c12066, in12066_1, in12066_2, c10399);
    wire[0:0] s12067, in12067_1, in12067_2;
    wire c12067;
    assign in12067_1 = {s10403[0]};
    assign in12067_2 = {s10404[0]};
    Full_Adder FA_12067(s12067, c12067, in12067_1, in12067_2, c10402);
    wire[0:0] s12068, in12068_1, in12068_2;
    wire c12068;
    assign in12068_1 = {s10406[0]};
    assign in12068_2 = {s10407[0]};
    Full_Adder FA_12068(s12068, c12068, in12068_1, in12068_2, s10405[0]);
    wire[0:0] s12069, in12069_1, in12069_2;
    wire c12069;
    assign in12069_1 = {s10409[0]};
    assign in12069_2 = {s10410[0]};
    Full_Adder FA_12069(s12069, c12069, in12069_1, in12069_2, s10408[0]);
    wire[0:0] s12070, in12070_1, in12070_2;
    wire c12070;
    assign in12070_1 = {s10412[0]};
    assign in12070_2 = {s10413[0]};
    Full_Adder FA_12070(s12070, c12070, in12070_1, in12070_2, s10411[0]);
    wire[0:0] s12071, in12071_1, in12071_2;
    wire c12071;
    assign in12071_1 = {c10404};
    assign in12071_2 = {c10405};
    Full_Adder FA_12071(s12071, c12071, in12071_1, in12071_2, c10403);
    wire[0:0] s12072, in12072_1, in12072_2;
    wire c12072;
    assign in12072_1 = {c10407};
    assign in12072_2 = {c10408};
    Full_Adder FA_12072(s12072, c12072, in12072_1, in12072_2, c10406);
    wire[0:0] s12073, in12073_1, in12073_2;
    wire c12073;
    assign in12073_1 = {c10410};
    assign in12073_2 = {c10411};
    Full_Adder FA_12073(s12073, c12073, in12073_1, in12073_2, c10409);
    wire[0:0] s12074, in12074_1, in12074_2;
    wire c12074;
    assign in12074_1 = {c10413};
    assign in12074_2 = {c10414};
    Full_Adder FA_12074(s12074, c12074, in12074_1, in12074_2, c10412);
    wire[0:0] s12075, in12075_1, in12075_2;
    wire c12075;
    assign in12075_1 = {s10416[0]};
    assign in12075_2 = {s10417[0]};
    Full_Adder FA_12075(s12075, c12075, in12075_1, in12075_2, c10415);
    wire[0:0] s12076, in12076_1, in12076_2;
    wire c12076;
    assign in12076_1 = {s10419[0]};
    assign in12076_2 = {s10420[0]};
    Full_Adder FA_12076(s12076, c12076, in12076_1, in12076_2, s10418[0]);
    wire[0:0] s12077, in12077_1, in12077_2;
    wire c12077;
    assign in12077_1 = {s10422[0]};
    assign in12077_2 = {s10423[0]};
    Full_Adder FA_12077(s12077, c12077, in12077_1, in12077_2, s10421[0]);
    wire[0:0] s12078, in12078_1, in12078_2;
    wire c12078;
    assign in12078_1 = {s10425[0]};
    assign in12078_2 = {s10426[0]};
    Full_Adder FA_12078(s12078, c12078, in12078_1, in12078_2, s10424[0]);
    wire[0:0] s12079, in12079_1, in12079_2;
    wire c12079;
    assign in12079_1 = {c10416};
    assign in12079_2 = {c10417};
    Full_Adder FA_12079(s12079, c12079, in12079_1, in12079_2, pp127[91]);
    wire[0:0] s12080, in12080_1, in12080_2;
    wire c12080;
    assign in12080_1 = {c10419};
    assign in12080_2 = {c10420};
    Full_Adder FA_12080(s12080, c12080, in12080_1, in12080_2, c10418);
    wire[0:0] s12081, in12081_1, in12081_2;
    wire c12081;
    assign in12081_1 = {c10422};
    assign in12081_2 = {c10423};
    Full_Adder FA_12081(s12081, c12081, in12081_1, in12081_2, c10421);
    wire[0:0] s12082, in12082_1, in12082_2;
    wire c12082;
    assign in12082_1 = {c10425};
    assign in12082_2 = {c10426};
    Full_Adder FA_12082(s12082, c12082, in12082_1, in12082_2, c10424);
    wire[0:0] s12083, in12083_1, in12083_2;
    wire c12083;
    assign in12083_1 = {c10428};
    assign in12083_2 = {s10429[0]};
    Full_Adder FA_12083(s12083, c12083, in12083_1, in12083_2, c10427);
    wire[0:0] s12084, in12084_1, in12084_2;
    wire c12084;
    assign in12084_1 = {s10431[0]};
    assign in12084_2 = {s10432[0]};
    Full_Adder FA_12084(s12084, c12084, in12084_1, in12084_2, s10430[0]);
    wire[0:0] s12085, in12085_1, in12085_2;
    wire c12085;
    assign in12085_1 = {s10434[0]};
    assign in12085_2 = {s10435[0]};
    Full_Adder FA_12085(s12085, c12085, in12085_1, in12085_2, s10433[0]);
    wire[0:0] s12086, in12086_1, in12086_2;
    wire c12086;
    assign in12086_1 = {s10437[0]};
    assign in12086_2 = {s10438[0]};
    Full_Adder FA_12086(s12086, c12086, in12086_1, in12086_2, s10436[0]);
    wire[0:0] s12087, in12087_1, in12087_2;
    wire c12087;
    assign in12087_1 = {pp126[93]};
    assign in12087_2 = {pp127[92]};
    Full_Adder FA_12087(s12087, c12087, in12087_1, in12087_2, pp125[94]);
    wire[0:0] s12088, in12088_1, in12088_2;
    wire c12088;
    assign in12088_1 = {c10430};
    assign in12088_2 = {c10431};
    Full_Adder FA_12088(s12088, c12088, in12088_1, in12088_2, c10429);
    wire[0:0] s12089, in12089_1, in12089_2;
    wire c12089;
    assign in12089_1 = {c10433};
    assign in12089_2 = {c10434};
    Full_Adder FA_12089(s12089, c12089, in12089_1, in12089_2, c10432);
    wire[0:0] s12090, in12090_1, in12090_2;
    wire c12090;
    assign in12090_1 = {c10436};
    assign in12090_2 = {c10437};
    Full_Adder FA_12090(s12090, c12090, in12090_1, in12090_2, c10435);
    wire[0:0] s12091, in12091_1, in12091_2;
    wire c12091;
    assign in12091_1 = {c10439};
    assign in12091_2 = {c10440};
    Full_Adder FA_12091(s12091, c12091, in12091_1, in12091_2, c10438);
    wire[0:0] s12092, in12092_1, in12092_2;
    wire c12092;
    assign in12092_1 = {s10442[0]};
    assign in12092_2 = {s10443[0]};
    Full_Adder FA_12092(s12092, c12092, in12092_1, in12092_2, s10441[0]);
    wire[0:0] s12093, in12093_1, in12093_2;
    wire c12093;
    assign in12093_1 = {s10445[0]};
    assign in12093_2 = {s10446[0]};
    Full_Adder FA_12093(s12093, c12093, in12093_1, in12093_2, s10444[0]);
    wire[0:0] s12094, in12094_1, in12094_2;
    wire c12094;
    assign in12094_1 = {s10448[0]};
    assign in12094_2 = {s10449[0]};
    Full_Adder FA_12094(s12094, c12094, in12094_1, in12094_2, s10447[0]);
    wire[0:0] s12095, in12095_1, in12095_2;
    wire c12095;
    assign in12095_1 = {pp124[96]};
    assign in12095_2 = {pp125[95]};
    Full_Adder FA_12095(s12095, c12095, in12095_1, in12095_2, pp123[97]);
    wire[0:0] s12096, in12096_1, in12096_2;
    wire c12096;
    assign in12096_1 = {pp127[93]};
    assign in12096_2 = {c10441};
    Full_Adder FA_12096(s12096, c12096, in12096_1, in12096_2, pp126[94]);
    wire[0:0] s12097, in12097_1, in12097_2;
    wire c12097;
    assign in12097_1 = {c10443};
    assign in12097_2 = {c10444};
    Full_Adder FA_12097(s12097, c12097, in12097_1, in12097_2, c10442);
    wire[0:0] s12098, in12098_1, in12098_2;
    wire c12098;
    assign in12098_1 = {c10446};
    assign in12098_2 = {c10447};
    Full_Adder FA_12098(s12098, c12098, in12098_1, in12098_2, c10445);
    wire[0:0] s12099, in12099_1, in12099_2;
    wire c12099;
    assign in12099_1 = {c10449};
    assign in12099_2 = {c10450};
    Full_Adder FA_12099(s12099, c12099, in12099_1, in12099_2, c10448);
    wire[0:0] s12100, in12100_1, in12100_2;
    wire c12100;
    assign in12100_1 = {s10452[0]};
    assign in12100_2 = {s10453[0]};
    Full_Adder FA_12100(s12100, c12100, in12100_1, in12100_2, c10451);
    wire[0:0] s12101, in12101_1, in12101_2;
    wire c12101;
    assign in12101_1 = {s10455[0]};
    assign in12101_2 = {s10456[0]};
    Full_Adder FA_12101(s12101, c12101, in12101_1, in12101_2, s10454[0]);
    wire[0:0] s12102, in12102_1, in12102_2;
    wire c12102;
    assign in12102_1 = {s10458[0]};
    assign in12102_2 = {s10459[0]};
    Full_Adder FA_12102(s12102, c12102, in12102_1, in12102_2, s10457[0]);
    wire[0:0] s12103, in12103_1, in12103_2;
    wire c12103;
    assign in12103_1 = {pp122[99]};
    assign in12103_2 = {pp123[98]};
    Full_Adder FA_12103(s12103, c12103, in12103_1, in12103_2, pp121[100]);
    wire[0:0] s12104, in12104_1, in12104_2;
    wire c12104;
    assign in12104_1 = {pp125[96]};
    assign in12104_2 = {pp126[95]};
    Full_Adder FA_12104(s12104, c12104, in12104_1, in12104_2, pp124[97]);
    wire[0:0] s12105, in12105_1, in12105_2;
    wire c12105;
    assign in12105_1 = {c10452};
    assign in12105_2 = {c10453};
    Full_Adder FA_12105(s12105, c12105, in12105_1, in12105_2, pp127[94]);
    wire[0:0] s12106, in12106_1, in12106_2;
    wire c12106;
    assign in12106_1 = {c10455};
    assign in12106_2 = {c10456};
    Full_Adder FA_12106(s12106, c12106, in12106_1, in12106_2, c10454);
    wire[0:0] s12107, in12107_1, in12107_2;
    wire c12107;
    assign in12107_1 = {c10458};
    assign in12107_2 = {c10459};
    Full_Adder FA_12107(s12107, c12107, in12107_1, in12107_2, c10457);
    wire[0:0] s12108, in12108_1, in12108_2;
    wire c12108;
    assign in12108_1 = {c10461};
    assign in12108_2 = {s10462[0]};
    Full_Adder FA_12108(s12108, c12108, in12108_1, in12108_2, c10460);
    wire[0:0] s12109, in12109_1, in12109_2;
    wire c12109;
    assign in12109_1 = {s10464[0]};
    assign in12109_2 = {s10465[0]};
    Full_Adder FA_12109(s12109, c12109, in12109_1, in12109_2, s10463[0]);
    wire[0:0] s12110, in12110_1, in12110_2;
    wire c12110;
    assign in12110_1 = {s10467[0]};
    assign in12110_2 = {s10468[0]};
    Full_Adder FA_12110(s12110, c12110, in12110_1, in12110_2, s10466[0]);
    wire[0:0] s12111, in12111_1, in12111_2;
    wire c12111;
    assign in12111_1 = {pp120[102]};
    assign in12111_2 = {pp121[101]};
    Full_Adder FA_12111(s12111, c12111, in12111_1, in12111_2, pp119[103]);
    wire[0:0] s12112, in12112_1, in12112_2;
    wire c12112;
    assign in12112_1 = {pp123[99]};
    assign in12112_2 = {pp124[98]};
    Full_Adder FA_12112(s12112, c12112, in12112_1, in12112_2, pp122[100]);
    wire[0:0] s12113, in12113_1, in12113_2;
    wire c12113;
    assign in12113_1 = {pp126[96]};
    assign in12113_2 = {pp127[95]};
    Full_Adder FA_12113(s12113, c12113, in12113_1, in12113_2, pp125[97]);
    wire[0:0] s12114, in12114_1, in12114_2;
    wire c12114;
    assign in12114_1 = {c10463};
    assign in12114_2 = {c10464};
    Full_Adder FA_12114(s12114, c12114, in12114_1, in12114_2, c10462);
    wire[0:0] s12115, in12115_1, in12115_2;
    wire c12115;
    assign in12115_1 = {c10466};
    assign in12115_2 = {c10467};
    Full_Adder FA_12115(s12115, c12115, in12115_1, in12115_2, c10465);
    wire[0:0] s12116, in12116_1, in12116_2;
    wire c12116;
    assign in12116_1 = {c10469};
    assign in12116_2 = {c10470};
    Full_Adder FA_12116(s12116, c12116, in12116_1, in12116_2, c10468);
    wire[0:0] s12117, in12117_1, in12117_2;
    wire c12117;
    assign in12117_1 = {s10472[0]};
    assign in12117_2 = {s10473[0]};
    Full_Adder FA_12117(s12117, c12117, in12117_1, in12117_2, s10471[0]);
    wire[0:0] s12118, in12118_1, in12118_2;
    wire c12118;
    assign in12118_1 = {s10475[0]};
    assign in12118_2 = {s10476[0]};
    Full_Adder FA_12118(s12118, c12118, in12118_1, in12118_2, s10474[0]);
    wire[0:0] s12119, in12119_1, in12119_2;
    wire c12119;
    assign in12119_1 = {pp118[105]};
    assign in12119_2 = {pp119[104]};
    Full_Adder FA_12119(s12119, c12119, in12119_1, in12119_2, pp117[106]);
    wire[0:0] s12120, in12120_1, in12120_2;
    wire c12120;
    assign in12120_1 = {pp121[102]};
    assign in12120_2 = {pp122[101]};
    Full_Adder FA_12120(s12120, c12120, in12120_1, in12120_2, pp120[103]);
    wire[0:0] s12121, in12121_1, in12121_2;
    wire c12121;
    assign in12121_1 = {pp124[99]};
    assign in12121_2 = {pp125[98]};
    Full_Adder FA_12121(s12121, c12121, in12121_1, in12121_2, pp123[100]);
    wire[0:0] s12122, in12122_1, in12122_2;
    wire c12122;
    assign in12122_1 = {pp127[96]};
    assign in12122_2 = {c10471};
    Full_Adder FA_12122(s12122, c12122, in12122_1, in12122_2, pp126[97]);
    wire[0:0] s12123, in12123_1, in12123_2;
    wire c12123;
    assign in12123_1 = {c10473};
    assign in12123_2 = {c10474};
    Full_Adder FA_12123(s12123, c12123, in12123_1, in12123_2, c10472);
    wire[0:0] s12124, in12124_1, in12124_2;
    wire c12124;
    assign in12124_1 = {c10476};
    assign in12124_2 = {c10477};
    Full_Adder FA_12124(s12124, c12124, in12124_1, in12124_2, c10475);
    wire[0:0] s12125, in12125_1, in12125_2;
    wire c12125;
    assign in12125_1 = {s10479[0]};
    assign in12125_2 = {s10480[0]};
    Full_Adder FA_12125(s12125, c12125, in12125_1, in12125_2, c10478);
    wire[0:0] s12126, in12126_1, in12126_2;
    wire c12126;
    assign in12126_1 = {s10482[0]};
    assign in12126_2 = {s10483[0]};
    Full_Adder FA_12126(s12126, c12126, in12126_1, in12126_2, s10481[0]);
    wire[0:0] s12127, in12127_1, in12127_2;
    wire c12127;
    assign in12127_1 = {pp116[108]};
    assign in12127_2 = {pp117[107]};
    Full_Adder FA_12127(s12127, c12127, in12127_1, in12127_2, pp115[109]);
    wire[0:0] s12128, in12128_1, in12128_2;
    wire c12128;
    assign in12128_1 = {pp119[105]};
    assign in12128_2 = {pp120[104]};
    Full_Adder FA_12128(s12128, c12128, in12128_1, in12128_2, pp118[106]);
    wire[0:0] s12129, in12129_1, in12129_2;
    wire c12129;
    assign in12129_1 = {pp122[102]};
    assign in12129_2 = {pp123[101]};
    Full_Adder FA_12129(s12129, c12129, in12129_1, in12129_2, pp121[103]);
    wire[0:0] s12130, in12130_1, in12130_2;
    wire c12130;
    assign in12130_1 = {pp125[99]};
    assign in12130_2 = {pp126[98]};
    Full_Adder FA_12130(s12130, c12130, in12130_1, in12130_2, pp124[100]);
    wire[0:0] s12131, in12131_1, in12131_2;
    wire c12131;
    assign in12131_1 = {c10479};
    assign in12131_2 = {c10480};
    Full_Adder FA_12131(s12131, c12131, in12131_1, in12131_2, pp127[97]);
    wire[0:0] s12132, in12132_1, in12132_2;
    wire c12132;
    assign in12132_1 = {c10482};
    assign in12132_2 = {c10483};
    Full_Adder FA_12132(s12132, c12132, in12132_1, in12132_2, c10481);
    wire[0:0] s12133, in12133_1, in12133_2;
    wire c12133;
    assign in12133_1 = {c10485};
    assign in12133_2 = {s10486[0]};
    Full_Adder FA_12133(s12133, c12133, in12133_1, in12133_2, c10484);
    wire[0:0] s12134, in12134_1, in12134_2;
    wire c12134;
    assign in12134_1 = {s10488[0]};
    assign in12134_2 = {s10489[0]};
    Full_Adder FA_12134(s12134, c12134, in12134_1, in12134_2, s10487[0]);
    wire[0:0] s12135, in12135_1, in12135_2;
    wire c12135;
    assign in12135_1 = {pp114[111]};
    assign in12135_2 = {pp115[110]};
    Full_Adder FA_12135(s12135, c12135, in12135_1, in12135_2, pp113[112]);
    wire[0:0] s12136, in12136_1, in12136_2;
    wire c12136;
    assign in12136_1 = {pp117[108]};
    assign in12136_2 = {pp118[107]};
    Full_Adder FA_12136(s12136, c12136, in12136_1, in12136_2, pp116[109]);
    wire[0:0] s12137, in12137_1, in12137_2;
    wire c12137;
    assign in12137_1 = {pp120[105]};
    assign in12137_2 = {pp121[104]};
    Full_Adder FA_12137(s12137, c12137, in12137_1, in12137_2, pp119[106]);
    wire[0:0] s12138, in12138_1, in12138_2;
    wire c12138;
    assign in12138_1 = {pp123[102]};
    assign in12138_2 = {pp124[101]};
    Full_Adder FA_12138(s12138, c12138, in12138_1, in12138_2, pp122[103]);
    wire[0:0] s12139, in12139_1, in12139_2;
    wire c12139;
    assign in12139_1 = {pp126[99]};
    assign in12139_2 = {pp127[98]};
    Full_Adder FA_12139(s12139, c12139, in12139_1, in12139_2, pp125[100]);
    wire[0:0] s12140, in12140_1, in12140_2;
    wire c12140;
    assign in12140_1 = {c10487};
    assign in12140_2 = {c10488};
    Full_Adder FA_12140(s12140, c12140, in12140_1, in12140_2, c10486);
    wire[0:0] s12141, in12141_1, in12141_2;
    wire c12141;
    assign in12141_1 = {c10490};
    assign in12141_2 = {c10491};
    Full_Adder FA_12141(s12141, c12141, in12141_1, in12141_2, c10489);
    wire[0:0] s12142, in12142_1, in12142_2;
    wire c12142;
    assign in12142_1 = {s10493[0]};
    assign in12142_2 = {s10494[0]};
    Full_Adder FA_12142(s12142, c12142, in12142_1, in12142_2, s10492[0]);
    wire[0:0] s12143, in12143_1, in12143_2;
    wire c12143;
    assign in12143_1 = {pp112[114]};
    assign in12143_2 = {pp113[113]};
    Full_Adder FA_12143(s12143, c12143, in12143_1, in12143_2, pp111[115]);
    wire[0:0] s12144, in12144_1, in12144_2;
    wire c12144;
    assign in12144_1 = {pp115[111]};
    assign in12144_2 = {pp116[110]};
    Full_Adder FA_12144(s12144, c12144, in12144_1, in12144_2, pp114[112]);
    wire[0:0] s12145, in12145_1, in12145_2;
    wire c12145;
    assign in12145_1 = {pp118[108]};
    assign in12145_2 = {pp119[107]};
    Full_Adder FA_12145(s12145, c12145, in12145_1, in12145_2, pp117[109]);
    wire[0:0] s12146, in12146_1, in12146_2;
    wire c12146;
    assign in12146_1 = {pp121[105]};
    assign in12146_2 = {pp122[104]};
    Full_Adder FA_12146(s12146, c12146, in12146_1, in12146_2, pp120[106]);
    wire[0:0] s12147, in12147_1, in12147_2;
    wire c12147;
    assign in12147_1 = {pp124[102]};
    assign in12147_2 = {pp125[101]};
    Full_Adder FA_12147(s12147, c12147, in12147_1, in12147_2, pp123[103]);
    wire[0:0] s12148, in12148_1, in12148_2;
    wire c12148;
    assign in12148_1 = {pp127[99]};
    assign in12148_2 = {c10492};
    Full_Adder FA_12148(s12148, c12148, in12148_1, in12148_2, pp126[100]);
    wire[0:0] s12149, in12149_1, in12149_2;
    wire c12149;
    assign in12149_1 = {c10494};
    assign in12149_2 = {c10495};
    Full_Adder FA_12149(s12149, c12149, in12149_1, in12149_2, c10493);
    wire[0:0] s12150, in12150_1, in12150_2;
    wire c12150;
    assign in12150_1 = {s10497[0]};
    assign in12150_2 = {s10498[0]};
    Full_Adder FA_12150(s12150, c12150, in12150_1, in12150_2, c10496);
    wire[0:0] s12151, in12151_1, in12151_2;
    wire c12151;
    assign in12151_1 = {pp110[117]};
    assign in12151_2 = {pp111[116]};
    Full_Adder FA_12151(s12151, c12151, in12151_1, in12151_2, pp109[118]);
    wire[0:0] s12152, in12152_1, in12152_2;
    wire c12152;
    assign in12152_1 = {pp113[114]};
    assign in12152_2 = {pp114[113]};
    Full_Adder FA_12152(s12152, c12152, in12152_1, in12152_2, pp112[115]);
    wire[0:0] s12153, in12153_1, in12153_2;
    wire c12153;
    assign in12153_1 = {pp116[111]};
    assign in12153_2 = {pp117[110]};
    Full_Adder FA_12153(s12153, c12153, in12153_1, in12153_2, pp115[112]);
    wire[0:0] s12154, in12154_1, in12154_2;
    wire c12154;
    assign in12154_1 = {pp119[108]};
    assign in12154_2 = {pp120[107]};
    Full_Adder FA_12154(s12154, c12154, in12154_1, in12154_2, pp118[109]);
    wire[0:0] s12155, in12155_1, in12155_2;
    wire c12155;
    assign in12155_1 = {pp122[105]};
    assign in12155_2 = {pp123[104]};
    Full_Adder FA_12155(s12155, c12155, in12155_1, in12155_2, pp121[106]);
    wire[0:0] s12156, in12156_1, in12156_2;
    wire c12156;
    assign in12156_1 = {pp125[102]};
    assign in12156_2 = {pp126[101]};
    Full_Adder FA_12156(s12156, c12156, in12156_1, in12156_2, pp124[103]);
    wire[0:0] s12157, in12157_1, in12157_2;
    wire c12157;
    assign in12157_1 = {c10497};
    assign in12157_2 = {c10498};
    Full_Adder FA_12157(s12157, c12157, in12157_1, in12157_2, pp127[100]);
    wire[0:0] s12158, in12158_1, in12158_2;
    wire c12158;
    assign in12158_1 = {c10500};
    assign in12158_2 = {s10501[0]};
    Full_Adder FA_12158(s12158, c12158, in12158_1, in12158_2, c10499);
    wire[0:0] s12159, in12159_1, in12159_2;
    wire c12159;
    assign in12159_1 = {pp108[120]};
    assign in12159_2 = {pp109[119]};
    Full_Adder FA_12159(s12159, c12159, in12159_1, in12159_2, pp107[121]);
    wire[0:0] s12160, in12160_1, in12160_2;
    wire c12160;
    assign in12160_1 = {pp111[117]};
    assign in12160_2 = {pp112[116]};
    Full_Adder FA_12160(s12160, c12160, in12160_1, in12160_2, pp110[118]);
    wire[0:0] s12161, in12161_1, in12161_2;
    wire c12161;
    assign in12161_1 = {pp114[114]};
    assign in12161_2 = {pp115[113]};
    Full_Adder FA_12161(s12161, c12161, in12161_1, in12161_2, pp113[115]);
    wire[0:0] s12162, in12162_1, in12162_2;
    wire c12162;
    assign in12162_1 = {pp117[111]};
    assign in12162_2 = {pp118[110]};
    Full_Adder FA_12162(s12162, c12162, in12162_1, in12162_2, pp116[112]);
    wire[0:0] s12163, in12163_1, in12163_2;
    wire c12163;
    assign in12163_1 = {pp120[108]};
    assign in12163_2 = {pp121[107]};
    Full_Adder FA_12163(s12163, c12163, in12163_1, in12163_2, pp119[109]);
    wire[0:0] s12164, in12164_1, in12164_2;
    wire c12164;
    assign in12164_1 = {pp123[105]};
    assign in12164_2 = {pp124[104]};
    Full_Adder FA_12164(s12164, c12164, in12164_1, in12164_2, pp122[106]);
    wire[0:0] s12165, in12165_1, in12165_2;
    wire c12165;
    assign in12165_1 = {pp126[102]};
    assign in12165_2 = {pp127[101]};
    Full_Adder FA_12165(s12165, c12165, in12165_1, in12165_2, pp125[103]);
    wire[0:0] s12166, in12166_1, in12166_2;
    wire c12166;
    assign in12166_1 = {c10502};
    assign in12166_2 = {c10503};
    Full_Adder FA_12166(s12166, c12166, in12166_1, in12166_2, c10501);
    wire[0:0] s12167, in12167_1, in12167_2;
    wire c12167;
    assign in12167_1 = {pp106[123]};
    assign in12167_2 = {pp107[122]};
    Full_Adder FA_12167(s12167, c12167, in12167_1, in12167_2, pp105[124]);
    wire[0:0] s12168, in12168_1, in12168_2;
    wire c12168;
    assign in12168_1 = {pp109[120]};
    assign in12168_2 = {pp110[119]};
    Full_Adder FA_12168(s12168, c12168, in12168_1, in12168_2, pp108[121]);
    wire[0:0] s12169, in12169_1, in12169_2;
    wire c12169;
    assign in12169_1 = {pp112[117]};
    assign in12169_2 = {pp113[116]};
    Full_Adder FA_12169(s12169, c12169, in12169_1, in12169_2, pp111[118]);
    wire[0:0] s12170, in12170_1, in12170_2;
    wire c12170;
    assign in12170_1 = {pp115[114]};
    assign in12170_2 = {pp116[113]};
    Full_Adder FA_12170(s12170, c12170, in12170_1, in12170_2, pp114[115]);
    wire[0:0] s12171, in12171_1, in12171_2;
    wire c12171;
    assign in12171_1 = {pp118[111]};
    assign in12171_2 = {pp119[110]};
    Full_Adder FA_12171(s12171, c12171, in12171_1, in12171_2, pp117[112]);
    wire[0:0] s12172, in12172_1, in12172_2;
    wire c12172;
    assign in12172_1 = {pp121[108]};
    assign in12172_2 = {pp122[107]};
    Full_Adder FA_12172(s12172, c12172, in12172_1, in12172_2, pp120[109]);
    wire[0:0] s12173, in12173_1, in12173_2;
    wire c12173;
    assign in12173_1 = {pp124[105]};
    assign in12173_2 = {pp125[104]};
    Full_Adder FA_12173(s12173, c12173, in12173_1, in12173_2, pp123[106]);
    wire[0:0] s12174, in12174_1, in12174_2;
    wire c12174;
    assign in12174_1 = {pp127[102]};
    assign in12174_2 = {c10504};
    Full_Adder FA_12174(s12174, c12174, in12174_1, in12174_2, pp126[103]);
    wire[0:0] s12175, in12175_1, in12175_2;
    wire c12175;
    assign in12175_1 = {pp104[126]};
    assign in12175_2 = {pp105[125]};
    Full_Adder FA_12175(s12175, c12175, in12175_1, in12175_2, pp103[127]);
    wire[0:0] s12176, in12176_1, in12176_2;
    wire c12176;
    assign in12176_1 = {pp107[123]};
    assign in12176_2 = {pp108[122]};
    Full_Adder FA_12176(s12176, c12176, in12176_1, in12176_2, pp106[124]);
    wire[0:0] s12177, in12177_1, in12177_2;
    wire c12177;
    assign in12177_1 = {pp110[120]};
    assign in12177_2 = {pp111[119]};
    Full_Adder FA_12177(s12177, c12177, in12177_1, in12177_2, pp109[121]);
    wire[0:0] s12178, in12178_1, in12178_2;
    wire c12178;
    assign in12178_1 = {pp113[117]};
    assign in12178_2 = {pp114[116]};
    Full_Adder FA_12178(s12178, c12178, in12178_1, in12178_2, pp112[118]);
    wire[0:0] s12179, in12179_1, in12179_2;
    wire c12179;
    assign in12179_1 = {pp116[114]};
    assign in12179_2 = {pp117[113]};
    Full_Adder FA_12179(s12179, c12179, in12179_1, in12179_2, pp115[115]);
    wire[0:0] s12180, in12180_1, in12180_2;
    wire c12180;
    assign in12180_1 = {pp119[111]};
    assign in12180_2 = {pp120[110]};
    Full_Adder FA_12180(s12180, c12180, in12180_1, in12180_2, pp118[112]);
    wire[0:0] s12181, in12181_1, in12181_2;
    wire c12181;
    assign in12181_1 = {pp122[108]};
    assign in12181_2 = {pp123[107]};
    Full_Adder FA_12181(s12181, c12181, in12181_1, in12181_2, pp121[109]);
    wire[0:0] s12182, in12182_1, in12182_2;
    wire c12182;
    assign in12182_1 = {pp125[105]};
    assign in12182_2 = {pp126[104]};
    Full_Adder FA_12182(s12182, c12182, in12182_1, in12182_2, pp124[106]);
    wire[0:0] s12183, in12183_1, in12183_2;
    wire c12183;
    assign in12183_1 = {pp105[126]};
    assign in12183_2 = {pp106[125]};
    Full_Adder FA_12183(s12183, c12183, in12183_1, in12183_2, pp104[127]);
    wire[0:0] s12184, in12184_1, in12184_2;
    wire c12184;
    assign in12184_1 = {pp108[123]};
    assign in12184_2 = {pp109[122]};
    Full_Adder FA_12184(s12184, c12184, in12184_1, in12184_2, pp107[124]);
    wire[0:0] s12185, in12185_1, in12185_2;
    wire c12185;
    assign in12185_1 = {pp111[120]};
    assign in12185_2 = {pp112[119]};
    Full_Adder FA_12185(s12185, c12185, in12185_1, in12185_2, pp110[121]);
    wire[0:0] s12186, in12186_1, in12186_2;
    wire c12186;
    assign in12186_1 = {pp114[117]};
    assign in12186_2 = {pp115[116]};
    Full_Adder FA_12186(s12186, c12186, in12186_1, in12186_2, pp113[118]);
    wire[0:0] s12187, in12187_1, in12187_2;
    wire c12187;
    assign in12187_1 = {pp117[114]};
    assign in12187_2 = {pp118[113]};
    Full_Adder FA_12187(s12187, c12187, in12187_1, in12187_2, pp116[115]);
    wire[0:0] s12188, in12188_1, in12188_2;
    wire c12188;
    assign in12188_1 = {pp120[111]};
    assign in12188_2 = {pp121[110]};
    Full_Adder FA_12188(s12188, c12188, in12188_1, in12188_2, pp119[112]);
    wire[0:0] s12189, in12189_1, in12189_2;
    wire c12189;
    assign in12189_1 = {pp123[108]};
    assign in12189_2 = {pp124[107]};
    Full_Adder FA_12189(s12189, c12189, in12189_1, in12189_2, pp122[109]);
    wire[0:0] s12190, in12190_1, in12190_2;
    wire c12190;
    assign in12190_1 = {pp106[126]};
    assign in12190_2 = {pp107[125]};
    Full_Adder FA_12190(s12190, c12190, in12190_1, in12190_2, pp105[127]);
    wire[0:0] s12191, in12191_1, in12191_2;
    wire c12191;
    assign in12191_1 = {pp109[123]};
    assign in12191_2 = {pp110[122]};
    Full_Adder FA_12191(s12191, c12191, in12191_1, in12191_2, pp108[124]);
    wire[0:0] s12192, in12192_1, in12192_2;
    wire c12192;
    assign in12192_1 = {pp112[120]};
    assign in12192_2 = {pp113[119]};
    Full_Adder FA_12192(s12192, c12192, in12192_1, in12192_2, pp111[121]);
    wire[0:0] s12193, in12193_1, in12193_2;
    wire c12193;
    assign in12193_1 = {pp115[117]};
    assign in12193_2 = {pp116[116]};
    Full_Adder FA_12193(s12193, c12193, in12193_1, in12193_2, pp114[118]);
    wire[0:0] s12194, in12194_1, in12194_2;
    wire c12194;
    assign in12194_1 = {pp118[114]};
    assign in12194_2 = {pp119[113]};
    Full_Adder FA_12194(s12194, c12194, in12194_1, in12194_2, pp117[115]);
    wire[0:0] s12195, in12195_1, in12195_2;
    wire c12195;
    assign in12195_1 = {pp121[111]};
    assign in12195_2 = {pp122[110]};
    Full_Adder FA_12195(s12195, c12195, in12195_1, in12195_2, pp120[112]);
    wire[0:0] s12196, in12196_1, in12196_2;
    wire c12196;
    assign in12196_1 = {pp107[126]};
    assign in12196_2 = {pp108[125]};
    Full_Adder FA_12196(s12196, c12196, in12196_1, in12196_2, pp106[127]);
    wire[0:0] s12197, in12197_1, in12197_2;
    wire c12197;
    assign in12197_1 = {pp110[123]};
    assign in12197_2 = {pp111[122]};
    Full_Adder FA_12197(s12197, c12197, in12197_1, in12197_2, pp109[124]);
    wire[0:0] s12198, in12198_1, in12198_2;
    wire c12198;
    assign in12198_1 = {pp113[120]};
    assign in12198_2 = {pp114[119]};
    Full_Adder FA_12198(s12198, c12198, in12198_1, in12198_2, pp112[121]);
    wire[0:0] s12199, in12199_1, in12199_2;
    wire c12199;
    assign in12199_1 = {pp116[117]};
    assign in12199_2 = {pp117[116]};
    Full_Adder FA_12199(s12199, c12199, in12199_1, in12199_2, pp115[118]);
    wire[0:0] s12200, in12200_1, in12200_2;
    wire c12200;
    assign in12200_1 = {pp119[114]};
    assign in12200_2 = {pp120[113]};
    Full_Adder FA_12200(s12200, c12200, in12200_1, in12200_2, pp118[115]);
    wire[0:0] s12201, in12201_1, in12201_2;
    wire c12201;
    assign in12201_1 = {pp108[126]};
    assign in12201_2 = {pp109[125]};
    Full_Adder FA_12201(s12201, c12201, in12201_1, in12201_2, pp107[127]);
    wire[0:0] s12202, in12202_1, in12202_2;
    wire c12202;
    assign in12202_1 = {pp111[123]};
    assign in12202_2 = {pp112[122]};
    Full_Adder FA_12202(s12202, c12202, in12202_1, in12202_2, pp110[124]);
    wire[0:0] s12203, in12203_1, in12203_2;
    wire c12203;
    assign in12203_1 = {pp114[120]};
    assign in12203_2 = {pp115[119]};
    Full_Adder FA_12203(s12203, c12203, in12203_1, in12203_2, pp113[121]);
    wire[0:0] s12204, in12204_1, in12204_2;
    wire c12204;
    assign in12204_1 = {pp117[117]};
    assign in12204_2 = {pp118[116]};
    Full_Adder FA_12204(s12204, c12204, in12204_1, in12204_2, pp116[118]);
    wire[0:0] s12205, in12205_1, in12205_2;
    wire c12205;
    assign in12205_1 = {pp109[126]};
    assign in12205_2 = {pp110[125]};
    Full_Adder FA_12205(s12205, c12205, in12205_1, in12205_2, pp108[127]);
    wire[0:0] s12206, in12206_1, in12206_2;
    wire c12206;
    assign in12206_1 = {pp112[123]};
    assign in12206_2 = {pp113[122]};
    Full_Adder FA_12206(s12206, c12206, in12206_1, in12206_2, pp111[124]);
    wire[0:0] s12207, in12207_1, in12207_2;
    wire c12207;
    assign in12207_1 = {pp115[120]};
    assign in12207_2 = {pp116[119]};
    Full_Adder FA_12207(s12207, c12207, in12207_1, in12207_2, pp114[121]);
    wire[0:0] s12208, in12208_1, in12208_2;
    wire c12208;
    assign in12208_1 = {pp110[126]};
    assign in12208_2 = {pp111[125]};
    Full_Adder FA_12208(s12208, c12208, in12208_1, in12208_2, pp109[127]);
    wire[0:0] s12209, in12209_1, in12209_2;
    wire c12209;
    assign in12209_1 = {pp113[123]};
    assign in12209_2 = {pp114[122]};
    Full_Adder FA_12209(s12209, c12209, in12209_1, in12209_2, pp112[124]);
    wire[0:0] s12210, in12210_1, in12210_2;
    wire c12210;
    assign in12210_1 = {pp111[126]};
    assign in12210_2 = {pp112[125]};
    Full_Adder FA_12210(s12210, c12210, in12210_1, in12210_2, pp110[127]);

    /*Stage 6*/
    wire[0:0] s12211, in12211_1, in12211_2;
    wire c12211;
    assign in12211_1 = {pp0[12]};
    assign in12211_2 = {pp1[11]};
    Half_Adder HA_12211(s12211, c12211, in12211_1, in12211_2);
    wire[0:0] s12212, in12212_1, in12212_2;
    wire c12212;
    assign in12212_1 = {pp1[12]};
    assign in12212_2 = {pp2[11]};
    Full_Adder FA_12212(s12212, c12212, in12212_1, in12212_2, pp0[13]);
    wire[0:0] s12213, in12213_1, in12213_2;
    wire c12213;
    assign in12213_1 = {pp3[10]};
    assign in12213_2 = {pp4[9]};
    Half_Adder HA_12213(s12213, c12213, in12213_1, in12213_2);
    wire[0:0] s12214, in12214_1, in12214_2;
    wire c12214;
    assign in12214_1 = {pp1[13]};
    assign in12214_2 = {pp2[12]};
    Full_Adder FA_12214(s12214, c12214, in12214_1, in12214_2, pp0[14]);
    wire[0:0] s12215, in12215_1, in12215_2;
    wire c12215;
    assign in12215_1 = {pp4[10]};
    assign in12215_2 = {pp5[9]};
    Full_Adder FA_12215(s12215, c12215, in12215_1, in12215_2, pp3[11]);
    wire[0:0] s12216, in12216_1, in12216_2;
    wire c12216;
    assign in12216_1 = {pp6[8]};
    assign in12216_2 = {pp7[7]};
    Half_Adder HA_12216(s12216, c12216, in12216_1, in12216_2);
    wire[0:0] s12217, in12217_1, in12217_2;
    wire c12217;
    assign in12217_1 = {pp1[14]};
    assign in12217_2 = {pp2[13]};
    Full_Adder FA_12217(s12217, c12217, in12217_1, in12217_2, pp0[15]);
    wire[0:0] s12218, in12218_1, in12218_2;
    wire c12218;
    assign in12218_1 = {pp4[11]};
    assign in12218_2 = {pp5[10]};
    Full_Adder FA_12218(s12218, c12218, in12218_1, in12218_2, pp3[12]);
    wire[0:0] s12219, in12219_1, in12219_2;
    wire c12219;
    assign in12219_1 = {pp7[8]};
    assign in12219_2 = {pp8[7]};
    Full_Adder FA_12219(s12219, c12219, in12219_1, in12219_2, pp6[9]);
    wire[0:0] s12220, in12220_1, in12220_2;
    wire c12220;
    assign in12220_1 = {pp9[6]};
    assign in12220_2 = {pp10[5]};
    Half_Adder HA_12220(s12220, c12220, in12220_1, in12220_2);
    wire[0:0] s12221, in12221_1, in12221_2;
    wire c12221;
    assign in12221_1 = {pp1[15]};
    assign in12221_2 = {pp2[14]};
    Full_Adder FA_12221(s12221, c12221, in12221_1, in12221_2, pp0[16]);
    wire[0:0] s12222, in12222_1, in12222_2;
    wire c12222;
    assign in12222_1 = {pp4[12]};
    assign in12222_2 = {pp5[11]};
    Full_Adder FA_12222(s12222, c12222, in12222_1, in12222_2, pp3[13]);
    wire[0:0] s12223, in12223_1, in12223_2;
    wire c12223;
    assign in12223_1 = {pp7[9]};
    assign in12223_2 = {pp8[8]};
    Full_Adder FA_12223(s12223, c12223, in12223_1, in12223_2, pp6[10]);
    wire[0:0] s12224, in12224_1, in12224_2;
    wire c12224;
    assign in12224_1 = {pp10[6]};
    assign in12224_2 = {pp11[5]};
    Full_Adder FA_12224(s12224, c12224, in12224_1, in12224_2, pp9[7]);
    wire[0:0] s12225, in12225_1, in12225_2;
    wire c12225;
    assign in12225_1 = {pp12[4]};
    assign in12225_2 = {pp13[3]};
    Half_Adder HA_12225(s12225, c12225, in12225_1, in12225_2);
    wire[0:0] s12226, in12226_1, in12226_2;
    wire c12226;
    assign in12226_1 = {pp1[16]};
    assign in12226_2 = {pp2[15]};
    Full_Adder FA_12226(s12226, c12226, in12226_1, in12226_2, pp0[17]);
    wire[0:0] s12227, in12227_1, in12227_2;
    wire c12227;
    assign in12227_1 = {pp4[13]};
    assign in12227_2 = {pp5[12]};
    Full_Adder FA_12227(s12227, c12227, in12227_1, in12227_2, pp3[14]);
    wire[0:0] s12228, in12228_1, in12228_2;
    wire c12228;
    assign in12228_1 = {pp7[10]};
    assign in12228_2 = {pp8[9]};
    Full_Adder FA_12228(s12228, c12228, in12228_1, in12228_2, pp6[11]);
    wire[0:0] s12229, in12229_1, in12229_2;
    wire c12229;
    assign in12229_1 = {pp10[7]};
    assign in12229_2 = {pp11[6]};
    Full_Adder FA_12229(s12229, c12229, in12229_1, in12229_2, pp9[8]);
    wire[0:0] s12230, in12230_1, in12230_2;
    wire c12230;
    assign in12230_1 = {pp13[4]};
    assign in12230_2 = {pp14[3]};
    Full_Adder FA_12230(s12230, c12230, in12230_1, in12230_2, pp12[5]);
    wire[0:0] s12231, in12231_1, in12231_2;
    wire c12231;
    assign in12231_1 = {pp15[2]};
    assign in12231_2 = {pp16[1]};
    Half_Adder HA_12231(s12231, c12231, in12231_1, in12231_2);
    wire[0:0] s12232, in12232_1, in12232_2;
    wire c12232;
    assign in12232_1 = {pp3[15]};
    assign in12232_2 = {pp4[14]};
    Full_Adder FA_12232(s12232, c12232, in12232_1, in12232_2, pp2[16]);
    wire[0:0] s12233, in12233_1, in12233_2;
    wire c12233;
    assign in12233_1 = {pp6[12]};
    assign in12233_2 = {pp7[11]};
    Full_Adder FA_12233(s12233, c12233, in12233_1, in12233_2, pp5[13]);
    wire[0:0] s12234, in12234_1, in12234_2;
    wire c12234;
    assign in12234_1 = {pp9[9]};
    assign in12234_2 = {pp10[8]};
    Full_Adder FA_12234(s12234, c12234, in12234_1, in12234_2, pp8[10]);
    wire[0:0] s12235, in12235_1, in12235_2;
    wire c12235;
    assign in12235_1 = {pp12[6]};
    assign in12235_2 = {pp13[5]};
    Full_Adder FA_12235(s12235, c12235, in12235_1, in12235_2, pp11[7]);
    wire[0:0] s12236, in12236_1, in12236_2;
    wire c12236;
    assign in12236_1 = {pp15[3]};
    assign in12236_2 = {pp16[2]};
    Full_Adder FA_12236(s12236, c12236, in12236_1, in12236_2, pp14[4]);
    wire[0:0] s12237, in12237_1, in12237_2;
    wire c12237;
    assign in12237_1 = {pp18[0]};
    assign in12237_2 = {s10507[0]};
    Full_Adder FA_12237(s12237, c12237, in12237_1, in12237_2, pp17[1]);
    wire[0:0] s12238, in12238_1, in12238_2;
    wire c12238;
    assign in12238_1 = {pp6[13]};
    assign in12238_2 = {pp7[12]};
    Full_Adder FA_12238(s12238, c12238, in12238_1, in12238_2, pp5[14]);
    wire[0:0] s12239, in12239_1, in12239_2;
    wire c12239;
    assign in12239_1 = {pp9[10]};
    assign in12239_2 = {pp10[9]};
    Full_Adder FA_12239(s12239, c12239, in12239_1, in12239_2, pp8[11]);
    wire[0:0] s12240, in12240_1, in12240_2;
    wire c12240;
    assign in12240_1 = {pp12[7]};
    assign in12240_2 = {pp13[6]};
    Full_Adder FA_12240(s12240, c12240, in12240_1, in12240_2, pp11[8]);
    wire[0:0] s12241, in12241_1, in12241_2;
    wire c12241;
    assign in12241_1 = {pp15[4]};
    assign in12241_2 = {pp16[3]};
    Full_Adder FA_12241(s12241, c12241, in12241_1, in12241_2, pp14[5]);
    wire[0:0] s12242, in12242_1, in12242_2;
    wire c12242;
    assign in12242_1 = {pp18[1]};
    assign in12242_2 = {pp19[0]};
    Full_Adder FA_12242(s12242, c12242, in12242_1, in12242_2, pp17[2]);
    wire[0:0] s12243, in12243_1, in12243_2;
    wire c12243;
    assign in12243_1 = {s10508[0]};
    assign in12243_2 = {s10509[0]};
    Full_Adder FA_12243(s12243, c12243, in12243_1, in12243_2, c10507);
    wire[0:0] s12244, in12244_1, in12244_2;
    wire c12244;
    assign in12244_1 = {pp9[11]};
    assign in12244_2 = {pp10[10]};
    Full_Adder FA_12244(s12244, c12244, in12244_1, in12244_2, pp8[12]);
    wire[0:0] s12245, in12245_1, in12245_2;
    wire c12245;
    assign in12245_1 = {pp12[8]};
    assign in12245_2 = {pp13[7]};
    Full_Adder FA_12245(s12245, c12245, in12245_1, in12245_2, pp11[9]);
    wire[0:0] s12246, in12246_1, in12246_2;
    wire c12246;
    assign in12246_1 = {pp15[5]};
    assign in12246_2 = {pp16[4]};
    Full_Adder FA_12246(s12246, c12246, in12246_1, in12246_2, pp14[6]);
    wire[0:0] s12247, in12247_1, in12247_2;
    wire c12247;
    assign in12247_1 = {pp18[2]};
    assign in12247_2 = {pp19[1]};
    Full_Adder FA_12247(s12247, c12247, in12247_1, in12247_2, pp17[3]);
    wire[0:0] s12248, in12248_1, in12248_2;
    wire c12248;
    assign in12248_1 = {c10508};
    assign in12248_2 = {c10509};
    Full_Adder FA_12248(s12248, c12248, in12248_1, in12248_2, pp20[0]);
    wire[0:0] s12249, in12249_1, in12249_2;
    wire c12249;
    assign in12249_1 = {s10511[0]};
    assign in12249_2 = {s10512[0]};
    Full_Adder FA_12249(s12249, c12249, in12249_1, in12249_2, s10510[0]);
    wire[0:0] s12250, in12250_1, in12250_2;
    wire c12250;
    assign in12250_1 = {pp12[9]};
    assign in12250_2 = {pp13[8]};
    Full_Adder FA_12250(s12250, c12250, in12250_1, in12250_2, pp11[10]);
    wire[0:0] s12251, in12251_1, in12251_2;
    wire c12251;
    assign in12251_1 = {pp15[6]};
    assign in12251_2 = {pp16[5]};
    Full_Adder FA_12251(s12251, c12251, in12251_1, in12251_2, pp14[7]);
    wire[0:0] s12252, in12252_1, in12252_2;
    wire c12252;
    assign in12252_1 = {pp18[3]};
    assign in12252_2 = {pp19[2]};
    Full_Adder FA_12252(s12252, c12252, in12252_1, in12252_2, pp17[4]);
    wire[0:0] s12253, in12253_1, in12253_2;
    wire c12253;
    assign in12253_1 = {pp21[0]};
    assign in12253_2 = {c10510};
    Full_Adder FA_12253(s12253, c12253, in12253_1, in12253_2, pp20[1]);
    wire[0:0] s12254, in12254_1, in12254_2;
    wire c12254;
    assign in12254_1 = {c10512};
    assign in12254_2 = {s10513[0]};
    Full_Adder FA_12254(s12254, c12254, in12254_1, in12254_2, c10511);
    wire[0:0] s12255, in12255_1, in12255_2;
    wire c12255;
    assign in12255_1 = {s10515[0]};
    assign in12255_2 = {s10516[0]};
    Full_Adder FA_12255(s12255, c12255, in12255_1, in12255_2, s10514[0]);
    wire[0:0] s12256, in12256_1, in12256_2;
    wire c12256;
    assign in12256_1 = {pp15[7]};
    assign in12256_2 = {pp16[6]};
    Full_Adder FA_12256(s12256, c12256, in12256_1, in12256_2, pp14[8]);
    wire[0:0] s12257, in12257_1, in12257_2;
    wire c12257;
    assign in12257_1 = {pp18[4]};
    assign in12257_2 = {pp19[3]};
    Full_Adder FA_12257(s12257, c12257, in12257_1, in12257_2, pp17[5]);
    wire[0:0] s12258, in12258_1, in12258_2;
    wire c12258;
    assign in12258_1 = {pp21[1]};
    assign in12258_2 = {pp22[0]};
    Full_Adder FA_12258(s12258, c12258, in12258_1, in12258_2, pp20[2]);
    wire[0:0] s12259, in12259_1, in12259_2;
    wire c12259;
    assign in12259_1 = {c10514};
    assign in12259_2 = {c10515};
    Full_Adder FA_12259(s12259, c12259, in12259_1, in12259_2, c10513);
    wire[0:0] s12260, in12260_1, in12260_2;
    wire c12260;
    assign in12260_1 = {s10517[0]};
    assign in12260_2 = {s10518[0]};
    Full_Adder FA_12260(s12260, c12260, in12260_1, in12260_2, c10516);
    wire[0:0] s12261, in12261_1, in12261_2;
    wire c12261;
    assign in12261_1 = {s10520[0]};
    assign in12261_2 = {s10521[0]};
    Full_Adder FA_12261(s12261, c12261, in12261_1, in12261_2, s10519[0]);
    wire[0:0] s12262, in12262_1, in12262_2;
    wire c12262;
    assign in12262_1 = {pp18[5]};
    assign in12262_2 = {pp19[4]};
    Full_Adder FA_12262(s12262, c12262, in12262_1, in12262_2, pp17[6]);
    wire[0:0] s12263, in12263_1, in12263_2;
    wire c12263;
    assign in12263_1 = {pp21[2]};
    assign in12263_2 = {pp22[1]};
    Full_Adder FA_12263(s12263, c12263, in12263_1, in12263_2, pp20[3]);
    wire[0:0] s12264, in12264_1, in12264_2;
    wire c12264;
    assign in12264_1 = {c10517};
    assign in12264_2 = {c10518};
    Full_Adder FA_12264(s12264, c12264, in12264_1, in12264_2, pp23[0]);
    wire[0:0] s12265, in12265_1, in12265_2;
    wire c12265;
    assign in12265_1 = {c10520};
    assign in12265_2 = {c10521};
    Full_Adder FA_12265(s12265, c12265, in12265_1, in12265_2, c10519);
    wire[0:0] s12266, in12266_1, in12266_2;
    wire c12266;
    assign in12266_1 = {s10523[0]};
    assign in12266_2 = {s10524[0]};
    Full_Adder FA_12266(s12266, c12266, in12266_1, in12266_2, s10522[0]);
    wire[0:0] s12267, in12267_1, in12267_2;
    wire c12267;
    assign in12267_1 = {s10526[0]};
    assign in12267_2 = {s10527[0]};
    Full_Adder FA_12267(s12267, c12267, in12267_1, in12267_2, s10525[0]);
    wire[0:0] s12268, in12268_1, in12268_2;
    wire c12268;
    assign in12268_1 = {pp21[3]};
    assign in12268_2 = {pp22[2]};
    Full_Adder FA_12268(s12268, c12268, in12268_1, in12268_2, pp20[4]);
    wire[0:0] s12269, in12269_1, in12269_2;
    wire c12269;
    assign in12269_1 = {pp24[0]};
    assign in12269_2 = {c10522};
    Full_Adder FA_12269(s12269, c12269, in12269_1, in12269_2, pp23[1]);
    wire[0:0] s12270, in12270_1, in12270_2;
    wire c12270;
    assign in12270_1 = {c10524};
    assign in12270_2 = {c10525};
    Full_Adder FA_12270(s12270, c12270, in12270_1, in12270_2, c10523);
    wire[0:0] s12271, in12271_1, in12271_2;
    wire c12271;
    assign in12271_1 = {c10527};
    assign in12271_2 = {s10528[0]};
    Full_Adder FA_12271(s12271, c12271, in12271_1, in12271_2, c10526);
    wire[0:0] s12272, in12272_1, in12272_2;
    wire c12272;
    assign in12272_1 = {s10530[0]};
    assign in12272_2 = {s10531[0]};
    Full_Adder FA_12272(s12272, c12272, in12272_1, in12272_2, s10529[0]);
    wire[0:0] s12273, in12273_1, in12273_2;
    wire c12273;
    assign in12273_1 = {s10533[0]};
    assign in12273_2 = {s10534[0]};
    Full_Adder FA_12273(s12273, c12273, in12273_1, in12273_2, s10532[0]);
    wire[0:0] s12274, in12274_1, in12274_2;
    wire c12274;
    assign in12274_1 = {pp24[1]};
    assign in12274_2 = {pp25[0]};
    Full_Adder FA_12274(s12274, c12274, in12274_1, in12274_2, pp23[2]);
    wire[0:0] s12275, in12275_1, in12275_2;
    wire c12275;
    assign in12275_1 = {c10529};
    assign in12275_2 = {c10530};
    Full_Adder FA_12275(s12275, c12275, in12275_1, in12275_2, c10528);
    wire[0:0] s12276, in12276_1, in12276_2;
    wire c12276;
    assign in12276_1 = {c10532};
    assign in12276_2 = {c10533};
    Full_Adder FA_12276(s12276, c12276, in12276_1, in12276_2, c10531);
    wire[0:0] s12277, in12277_1, in12277_2;
    wire c12277;
    assign in12277_1 = {s10535[0]};
    assign in12277_2 = {s10536[0]};
    Full_Adder FA_12277(s12277, c12277, in12277_1, in12277_2, c10534);
    wire[0:0] s12278, in12278_1, in12278_2;
    wire c12278;
    assign in12278_1 = {s10538[0]};
    assign in12278_2 = {s10539[0]};
    Full_Adder FA_12278(s12278, c12278, in12278_1, in12278_2, s10537[0]);
    wire[0:0] s12279, in12279_1, in12279_2;
    wire c12279;
    assign in12279_1 = {s10541[0]};
    assign in12279_2 = {s10542[0]};
    Full_Adder FA_12279(s12279, c12279, in12279_1, in12279_2, s10540[0]);
    wire[0:0] s12280, in12280_1, in12280_2;
    wire c12280;
    assign in12280_1 = {s8011[0]};
    assign in12280_2 = {c10535};
    Full_Adder FA_12280(s12280, c12280, in12280_1, in12280_2, pp26[0]);
    wire[0:0] s12281, in12281_1, in12281_2;
    wire c12281;
    assign in12281_1 = {c10537};
    assign in12281_2 = {c10538};
    Full_Adder FA_12281(s12281, c12281, in12281_1, in12281_2, c10536);
    wire[0:0] s12282, in12282_1, in12282_2;
    wire c12282;
    assign in12282_1 = {c10540};
    assign in12282_2 = {c10541};
    Full_Adder FA_12282(s12282, c12282, in12282_1, in12282_2, c10539);
    wire[0:0] s12283, in12283_1, in12283_2;
    wire c12283;
    assign in12283_1 = {s10543[0]};
    assign in12283_2 = {s10544[0]};
    Full_Adder FA_12283(s12283, c12283, in12283_1, in12283_2, c10542);
    wire[0:0] s12284, in12284_1, in12284_2;
    wire c12284;
    assign in12284_1 = {s10546[0]};
    assign in12284_2 = {s10547[0]};
    Full_Adder FA_12284(s12284, c12284, in12284_1, in12284_2, s10545[0]);
    wire[0:0] s12285, in12285_1, in12285_2;
    wire c12285;
    assign in12285_1 = {s10549[0]};
    assign in12285_2 = {s10550[0]};
    Full_Adder FA_12285(s12285, c12285, in12285_1, in12285_2, s10548[0]);
    wire[0:0] s12286, in12286_1, in12286_2;
    wire c12286;
    assign in12286_1 = {s8013[0]};
    assign in12286_2 = {c10543};
    Full_Adder FA_12286(s12286, c12286, in12286_1, in12286_2, s8012[0]);
    wire[0:0] s12287, in12287_1, in12287_2;
    wire c12287;
    assign in12287_1 = {c10545};
    assign in12287_2 = {c10546};
    Full_Adder FA_12287(s12287, c12287, in12287_1, in12287_2, c10544);
    wire[0:0] s12288, in12288_1, in12288_2;
    wire c12288;
    assign in12288_1 = {c10548};
    assign in12288_2 = {c10549};
    Full_Adder FA_12288(s12288, c12288, in12288_1, in12288_2, c10547);
    wire[0:0] s12289, in12289_1, in12289_2;
    wire c12289;
    assign in12289_1 = {s10551[0]};
    assign in12289_2 = {s10552[0]};
    Full_Adder FA_12289(s12289, c12289, in12289_1, in12289_2, c10550);
    wire[0:0] s12290, in12290_1, in12290_2;
    wire c12290;
    assign in12290_1 = {s10554[0]};
    assign in12290_2 = {s10555[0]};
    Full_Adder FA_12290(s12290, c12290, in12290_1, in12290_2, s10553[0]);
    wire[0:0] s12291, in12291_1, in12291_2;
    wire c12291;
    assign in12291_1 = {s10557[0]};
    assign in12291_2 = {s10558[0]};
    Full_Adder FA_12291(s12291, c12291, in12291_1, in12291_2, s10556[0]);
    wire[0:0] s12292, in12292_1, in12292_2;
    wire c12292;
    assign in12292_1 = {s8016[0]};
    assign in12292_2 = {c10551};
    Full_Adder FA_12292(s12292, c12292, in12292_1, in12292_2, s8015[0]);
    wire[0:0] s12293, in12293_1, in12293_2;
    wire c12293;
    assign in12293_1 = {c10553};
    assign in12293_2 = {c10554};
    Full_Adder FA_12293(s12293, c12293, in12293_1, in12293_2, c10552);
    wire[0:0] s12294, in12294_1, in12294_2;
    wire c12294;
    assign in12294_1 = {c10556};
    assign in12294_2 = {c10557};
    Full_Adder FA_12294(s12294, c12294, in12294_1, in12294_2, c10555);
    wire[0:0] s12295, in12295_1, in12295_2;
    wire c12295;
    assign in12295_1 = {s10559[0]};
    assign in12295_2 = {s10560[0]};
    Full_Adder FA_12295(s12295, c12295, in12295_1, in12295_2, c10558);
    wire[0:0] s12296, in12296_1, in12296_2;
    wire c12296;
    assign in12296_1 = {s10562[0]};
    assign in12296_2 = {s10563[0]};
    Full_Adder FA_12296(s12296, c12296, in12296_1, in12296_2, s10561[0]);
    wire[0:0] s12297, in12297_1, in12297_2;
    wire c12297;
    assign in12297_1 = {s10565[0]};
    assign in12297_2 = {s10566[0]};
    Full_Adder FA_12297(s12297, c12297, in12297_1, in12297_2, s10564[0]);
    wire[0:0] s12298, in12298_1, in12298_2;
    wire c12298;
    assign in12298_1 = {s8020[0]};
    assign in12298_2 = {c10559};
    Full_Adder FA_12298(s12298, c12298, in12298_1, in12298_2, s8019[0]);
    wire[0:0] s12299, in12299_1, in12299_2;
    wire c12299;
    assign in12299_1 = {c10561};
    assign in12299_2 = {c10562};
    Full_Adder FA_12299(s12299, c12299, in12299_1, in12299_2, c10560);
    wire[0:0] s12300, in12300_1, in12300_2;
    wire c12300;
    assign in12300_1 = {c10564};
    assign in12300_2 = {c10565};
    Full_Adder FA_12300(s12300, c12300, in12300_1, in12300_2, c10563);
    wire[0:0] s12301, in12301_1, in12301_2;
    wire c12301;
    assign in12301_1 = {s10567[0]};
    assign in12301_2 = {s10568[0]};
    Full_Adder FA_12301(s12301, c12301, in12301_1, in12301_2, c10566);
    wire[0:0] s12302, in12302_1, in12302_2;
    wire c12302;
    assign in12302_1 = {s10570[0]};
    assign in12302_2 = {s10571[0]};
    Full_Adder FA_12302(s12302, c12302, in12302_1, in12302_2, s10569[0]);
    wire[0:0] s12303, in12303_1, in12303_2;
    wire c12303;
    assign in12303_1 = {s10573[0]};
    assign in12303_2 = {s10574[0]};
    Full_Adder FA_12303(s12303, c12303, in12303_1, in12303_2, s10572[0]);
    wire[0:0] s12304, in12304_1, in12304_2;
    wire c12304;
    assign in12304_1 = {s8025[0]};
    assign in12304_2 = {c10567};
    Full_Adder FA_12304(s12304, c12304, in12304_1, in12304_2, s8024[0]);
    wire[0:0] s12305, in12305_1, in12305_2;
    wire c12305;
    assign in12305_1 = {c10569};
    assign in12305_2 = {c10570};
    Full_Adder FA_12305(s12305, c12305, in12305_1, in12305_2, c10568);
    wire[0:0] s12306, in12306_1, in12306_2;
    wire c12306;
    assign in12306_1 = {c10572};
    assign in12306_2 = {c10573};
    Full_Adder FA_12306(s12306, c12306, in12306_1, in12306_2, c10571);
    wire[0:0] s12307, in12307_1, in12307_2;
    wire c12307;
    assign in12307_1 = {s10575[0]};
    assign in12307_2 = {s10576[0]};
    Full_Adder FA_12307(s12307, c12307, in12307_1, in12307_2, c10574);
    wire[0:0] s12308, in12308_1, in12308_2;
    wire c12308;
    assign in12308_1 = {s10578[0]};
    assign in12308_2 = {s10579[0]};
    Full_Adder FA_12308(s12308, c12308, in12308_1, in12308_2, s10577[0]);
    wire[0:0] s12309, in12309_1, in12309_2;
    wire c12309;
    assign in12309_1 = {s10581[0]};
    assign in12309_2 = {s10582[0]};
    Full_Adder FA_12309(s12309, c12309, in12309_1, in12309_2, s10580[0]);
    wire[0:0] s12310, in12310_1, in12310_2;
    wire c12310;
    assign in12310_1 = {s8031[0]};
    assign in12310_2 = {c10575};
    Full_Adder FA_12310(s12310, c12310, in12310_1, in12310_2, s8030[0]);
    wire[0:0] s12311, in12311_1, in12311_2;
    wire c12311;
    assign in12311_1 = {c10577};
    assign in12311_2 = {c10578};
    Full_Adder FA_12311(s12311, c12311, in12311_1, in12311_2, c10576);
    wire[0:0] s12312, in12312_1, in12312_2;
    wire c12312;
    assign in12312_1 = {c10580};
    assign in12312_2 = {c10581};
    Full_Adder FA_12312(s12312, c12312, in12312_1, in12312_2, c10579);
    wire[0:0] s12313, in12313_1, in12313_2;
    wire c12313;
    assign in12313_1 = {s10583[0]};
    assign in12313_2 = {s10584[0]};
    Full_Adder FA_12313(s12313, c12313, in12313_1, in12313_2, c10582);
    wire[0:0] s12314, in12314_1, in12314_2;
    wire c12314;
    assign in12314_1 = {s10586[0]};
    assign in12314_2 = {s10587[0]};
    Full_Adder FA_12314(s12314, c12314, in12314_1, in12314_2, s10585[0]);
    wire[0:0] s12315, in12315_1, in12315_2;
    wire c12315;
    assign in12315_1 = {s10589[0]};
    assign in12315_2 = {s10590[0]};
    Full_Adder FA_12315(s12315, c12315, in12315_1, in12315_2, s10588[0]);
    wire[0:0] s12316, in12316_1, in12316_2;
    wire c12316;
    assign in12316_1 = {s8038[0]};
    assign in12316_2 = {c10583};
    Full_Adder FA_12316(s12316, c12316, in12316_1, in12316_2, s8037[0]);
    wire[0:0] s12317, in12317_1, in12317_2;
    wire c12317;
    assign in12317_1 = {c10585};
    assign in12317_2 = {c10586};
    Full_Adder FA_12317(s12317, c12317, in12317_1, in12317_2, c10584);
    wire[0:0] s12318, in12318_1, in12318_2;
    wire c12318;
    assign in12318_1 = {c10588};
    assign in12318_2 = {c10589};
    Full_Adder FA_12318(s12318, c12318, in12318_1, in12318_2, c10587);
    wire[0:0] s12319, in12319_1, in12319_2;
    wire c12319;
    assign in12319_1 = {s10591[0]};
    assign in12319_2 = {s10592[0]};
    Full_Adder FA_12319(s12319, c12319, in12319_1, in12319_2, c10590);
    wire[0:0] s12320, in12320_1, in12320_2;
    wire c12320;
    assign in12320_1 = {s10594[0]};
    assign in12320_2 = {s10595[0]};
    Full_Adder FA_12320(s12320, c12320, in12320_1, in12320_2, s10593[0]);
    wire[0:0] s12321, in12321_1, in12321_2;
    wire c12321;
    assign in12321_1 = {s10597[0]};
    assign in12321_2 = {s10598[0]};
    Full_Adder FA_12321(s12321, c12321, in12321_1, in12321_2, s10596[0]);
    wire[0:0] s12322, in12322_1, in12322_2;
    wire c12322;
    assign in12322_1 = {s8046[0]};
    assign in12322_2 = {c10591};
    Full_Adder FA_12322(s12322, c12322, in12322_1, in12322_2, s8045[0]);
    wire[0:0] s12323, in12323_1, in12323_2;
    wire c12323;
    assign in12323_1 = {c10593};
    assign in12323_2 = {c10594};
    Full_Adder FA_12323(s12323, c12323, in12323_1, in12323_2, c10592);
    wire[0:0] s12324, in12324_1, in12324_2;
    wire c12324;
    assign in12324_1 = {c10596};
    assign in12324_2 = {c10597};
    Full_Adder FA_12324(s12324, c12324, in12324_1, in12324_2, c10595);
    wire[0:0] s12325, in12325_1, in12325_2;
    wire c12325;
    assign in12325_1 = {s10599[0]};
    assign in12325_2 = {s10600[0]};
    Full_Adder FA_12325(s12325, c12325, in12325_1, in12325_2, c10598);
    wire[0:0] s12326, in12326_1, in12326_2;
    wire c12326;
    assign in12326_1 = {s10602[0]};
    assign in12326_2 = {s10603[0]};
    Full_Adder FA_12326(s12326, c12326, in12326_1, in12326_2, s10601[0]);
    wire[0:0] s12327, in12327_1, in12327_2;
    wire c12327;
    assign in12327_1 = {s10605[0]};
    assign in12327_2 = {s10606[0]};
    Full_Adder FA_12327(s12327, c12327, in12327_1, in12327_2, s10604[0]);
    wire[0:0] s12328, in12328_1, in12328_2;
    wire c12328;
    assign in12328_1 = {s8055[0]};
    assign in12328_2 = {c10599};
    Full_Adder FA_12328(s12328, c12328, in12328_1, in12328_2, s8054[0]);
    wire[0:0] s12329, in12329_1, in12329_2;
    wire c12329;
    assign in12329_1 = {c10601};
    assign in12329_2 = {c10602};
    Full_Adder FA_12329(s12329, c12329, in12329_1, in12329_2, c10600);
    wire[0:0] s12330, in12330_1, in12330_2;
    wire c12330;
    assign in12330_1 = {c10604};
    assign in12330_2 = {c10605};
    Full_Adder FA_12330(s12330, c12330, in12330_1, in12330_2, c10603);
    wire[0:0] s12331, in12331_1, in12331_2;
    wire c12331;
    assign in12331_1 = {s10607[0]};
    assign in12331_2 = {s10608[0]};
    Full_Adder FA_12331(s12331, c12331, in12331_1, in12331_2, c10606);
    wire[0:0] s12332, in12332_1, in12332_2;
    wire c12332;
    assign in12332_1 = {s10610[0]};
    assign in12332_2 = {s10611[0]};
    Full_Adder FA_12332(s12332, c12332, in12332_1, in12332_2, s10609[0]);
    wire[0:0] s12333, in12333_1, in12333_2;
    wire c12333;
    assign in12333_1 = {s10613[0]};
    assign in12333_2 = {s10614[0]};
    Full_Adder FA_12333(s12333, c12333, in12333_1, in12333_2, s10612[0]);
    wire[0:0] s12334, in12334_1, in12334_2;
    wire c12334;
    assign in12334_1 = {s8065[0]};
    assign in12334_2 = {c10607};
    Full_Adder FA_12334(s12334, c12334, in12334_1, in12334_2, s8064[0]);
    wire[0:0] s12335, in12335_1, in12335_2;
    wire c12335;
    assign in12335_1 = {c10609};
    assign in12335_2 = {c10610};
    Full_Adder FA_12335(s12335, c12335, in12335_1, in12335_2, c10608);
    wire[0:0] s12336, in12336_1, in12336_2;
    wire c12336;
    assign in12336_1 = {c10612};
    assign in12336_2 = {c10613};
    Full_Adder FA_12336(s12336, c12336, in12336_1, in12336_2, c10611);
    wire[0:0] s12337, in12337_1, in12337_2;
    wire c12337;
    assign in12337_1 = {s10615[0]};
    assign in12337_2 = {s10616[0]};
    Full_Adder FA_12337(s12337, c12337, in12337_1, in12337_2, c10614);
    wire[0:0] s12338, in12338_1, in12338_2;
    wire c12338;
    assign in12338_1 = {s10618[0]};
    assign in12338_2 = {s10619[0]};
    Full_Adder FA_12338(s12338, c12338, in12338_1, in12338_2, s10617[0]);
    wire[0:0] s12339, in12339_1, in12339_2;
    wire c12339;
    assign in12339_1 = {s10621[0]};
    assign in12339_2 = {s10622[0]};
    Full_Adder FA_12339(s12339, c12339, in12339_1, in12339_2, s10620[0]);
    wire[0:0] s12340, in12340_1, in12340_2;
    wire c12340;
    assign in12340_1 = {s8076[0]};
    assign in12340_2 = {c10615};
    Full_Adder FA_12340(s12340, c12340, in12340_1, in12340_2, s8075[0]);
    wire[0:0] s12341, in12341_1, in12341_2;
    wire c12341;
    assign in12341_1 = {c10617};
    assign in12341_2 = {c10618};
    Full_Adder FA_12341(s12341, c12341, in12341_1, in12341_2, c10616);
    wire[0:0] s12342, in12342_1, in12342_2;
    wire c12342;
    assign in12342_1 = {c10620};
    assign in12342_2 = {c10621};
    Full_Adder FA_12342(s12342, c12342, in12342_1, in12342_2, c10619);
    wire[0:0] s12343, in12343_1, in12343_2;
    wire c12343;
    assign in12343_1 = {s10623[0]};
    assign in12343_2 = {s10624[0]};
    Full_Adder FA_12343(s12343, c12343, in12343_1, in12343_2, c10622);
    wire[0:0] s12344, in12344_1, in12344_2;
    wire c12344;
    assign in12344_1 = {s10626[0]};
    assign in12344_2 = {s10627[0]};
    Full_Adder FA_12344(s12344, c12344, in12344_1, in12344_2, s10625[0]);
    wire[0:0] s12345, in12345_1, in12345_2;
    wire c12345;
    assign in12345_1 = {s10629[0]};
    assign in12345_2 = {s10630[0]};
    Full_Adder FA_12345(s12345, c12345, in12345_1, in12345_2, s10628[0]);
    wire[0:0] s12346, in12346_1, in12346_2;
    wire c12346;
    assign in12346_1 = {s8088[0]};
    assign in12346_2 = {c10623};
    Full_Adder FA_12346(s12346, c12346, in12346_1, in12346_2, s8087[0]);
    wire[0:0] s12347, in12347_1, in12347_2;
    wire c12347;
    assign in12347_1 = {c10625};
    assign in12347_2 = {c10626};
    Full_Adder FA_12347(s12347, c12347, in12347_1, in12347_2, c10624);
    wire[0:0] s12348, in12348_1, in12348_2;
    wire c12348;
    assign in12348_1 = {c10628};
    assign in12348_2 = {c10629};
    Full_Adder FA_12348(s12348, c12348, in12348_1, in12348_2, c10627);
    wire[0:0] s12349, in12349_1, in12349_2;
    wire c12349;
    assign in12349_1 = {s10631[0]};
    assign in12349_2 = {s10632[0]};
    Full_Adder FA_12349(s12349, c12349, in12349_1, in12349_2, c10630);
    wire[0:0] s12350, in12350_1, in12350_2;
    wire c12350;
    assign in12350_1 = {s10634[0]};
    assign in12350_2 = {s10635[0]};
    Full_Adder FA_12350(s12350, c12350, in12350_1, in12350_2, s10633[0]);
    wire[0:0] s12351, in12351_1, in12351_2;
    wire c12351;
    assign in12351_1 = {s10637[0]};
    assign in12351_2 = {s10638[0]};
    Full_Adder FA_12351(s12351, c12351, in12351_1, in12351_2, s10636[0]);
    wire[0:0] s12352, in12352_1, in12352_2;
    wire c12352;
    assign in12352_1 = {s8101[0]};
    assign in12352_2 = {c10631};
    Full_Adder FA_12352(s12352, c12352, in12352_1, in12352_2, s8100[0]);
    wire[0:0] s12353, in12353_1, in12353_2;
    wire c12353;
    assign in12353_1 = {c10633};
    assign in12353_2 = {c10634};
    Full_Adder FA_12353(s12353, c12353, in12353_1, in12353_2, c10632);
    wire[0:0] s12354, in12354_1, in12354_2;
    wire c12354;
    assign in12354_1 = {c10636};
    assign in12354_2 = {c10637};
    Full_Adder FA_12354(s12354, c12354, in12354_1, in12354_2, c10635);
    wire[0:0] s12355, in12355_1, in12355_2;
    wire c12355;
    assign in12355_1 = {s10639[0]};
    assign in12355_2 = {s10640[0]};
    Full_Adder FA_12355(s12355, c12355, in12355_1, in12355_2, c10638);
    wire[0:0] s12356, in12356_1, in12356_2;
    wire c12356;
    assign in12356_1 = {s10642[0]};
    assign in12356_2 = {s10643[0]};
    Full_Adder FA_12356(s12356, c12356, in12356_1, in12356_2, s10641[0]);
    wire[0:0] s12357, in12357_1, in12357_2;
    wire c12357;
    assign in12357_1 = {s10645[0]};
    assign in12357_2 = {s10646[0]};
    Full_Adder FA_12357(s12357, c12357, in12357_1, in12357_2, s10644[0]);
    wire[0:0] s12358, in12358_1, in12358_2;
    wire c12358;
    assign in12358_1 = {s8114[0]};
    assign in12358_2 = {c10639};
    Full_Adder FA_12358(s12358, c12358, in12358_1, in12358_2, s8113[0]);
    wire[0:0] s12359, in12359_1, in12359_2;
    wire c12359;
    assign in12359_1 = {c10641};
    assign in12359_2 = {c10642};
    Full_Adder FA_12359(s12359, c12359, in12359_1, in12359_2, c10640);
    wire[0:0] s12360, in12360_1, in12360_2;
    wire c12360;
    assign in12360_1 = {c10644};
    assign in12360_2 = {c10645};
    Full_Adder FA_12360(s12360, c12360, in12360_1, in12360_2, c10643);
    wire[0:0] s12361, in12361_1, in12361_2;
    wire c12361;
    assign in12361_1 = {s10647[0]};
    assign in12361_2 = {s10648[0]};
    Full_Adder FA_12361(s12361, c12361, in12361_1, in12361_2, c10646);
    wire[0:0] s12362, in12362_1, in12362_2;
    wire c12362;
    assign in12362_1 = {s10650[0]};
    assign in12362_2 = {s10651[0]};
    Full_Adder FA_12362(s12362, c12362, in12362_1, in12362_2, s10649[0]);
    wire[0:0] s12363, in12363_1, in12363_2;
    wire c12363;
    assign in12363_1 = {s10653[0]};
    assign in12363_2 = {s10654[0]};
    Full_Adder FA_12363(s12363, c12363, in12363_1, in12363_2, s10652[0]);
    wire[0:0] s12364, in12364_1, in12364_2;
    wire c12364;
    assign in12364_1 = {s8127[0]};
    assign in12364_2 = {c10647};
    Full_Adder FA_12364(s12364, c12364, in12364_1, in12364_2, s8126[0]);
    wire[0:0] s12365, in12365_1, in12365_2;
    wire c12365;
    assign in12365_1 = {c10649};
    assign in12365_2 = {c10650};
    Full_Adder FA_12365(s12365, c12365, in12365_1, in12365_2, c10648);
    wire[0:0] s12366, in12366_1, in12366_2;
    wire c12366;
    assign in12366_1 = {c10652};
    assign in12366_2 = {c10653};
    Full_Adder FA_12366(s12366, c12366, in12366_1, in12366_2, c10651);
    wire[0:0] s12367, in12367_1, in12367_2;
    wire c12367;
    assign in12367_1 = {s10655[0]};
    assign in12367_2 = {s10656[0]};
    Full_Adder FA_12367(s12367, c12367, in12367_1, in12367_2, c10654);
    wire[0:0] s12368, in12368_1, in12368_2;
    wire c12368;
    assign in12368_1 = {s10658[0]};
    assign in12368_2 = {s10659[0]};
    Full_Adder FA_12368(s12368, c12368, in12368_1, in12368_2, s10657[0]);
    wire[0:0] s12369, in12369_1, in12369_2;
    wire c12369;
    assign in12369_1 = {s10661[0]};
    assign in12369_2 = {s10662[0]};
    Full_Adder FA_12369(s12369, c12369, in12369_1, in12369_2, s10660[0]);
    wire[0:0] s12370, in12370_1, in12370_2;
    wire c12370;
    assign in12370_1 = {s8140[0]};
    assign in12370_2 = {c10655};
    Full_Adder FA_12370(s12370, c12370, in12370_1, in12370_2, s8139[0]);
    wire[0:0] s12371, in12371_1, in12371_2;
    wire c12371;
    assign in12371_1 = {c10657};
    assign in12371_2 = {c10658};
    Full_Adder FA_12371(s12371, c12371, in12371_1, in12371_2, c10656);
    wire[0:0] s12372, in12372_1, in12372_2;
    wire c12372;
    assign in12372_1 = {c10660};
    assign in12372_2 = {c10661};
    Full_Adder FA_12372(s12372, c12372, in12372_1, in12372_2, c10659);
    wire[0:0] s12373, in12373_1, in12373_2;
    wire c12373;
    assign in12373_1 = {s10663[0]};
    assign in12373_2 = {s10664[0]};
    Full_Adder FA_12373(s12373, c12373, in12373_1, in12373_2, c10662);
    wire[0:0] s12374, in12374_1, in12374_2;
    wire c12374;
    assign in12374_1 = {s10666[0]};
    assign in12374_2 = {s10667[0]};
    Full_Adder FA_12374(s12374, c12374, in12374_1, in12374_2, s10665[0]);
    wire[0:0] s12375, in12375_1, in12375_2;
    wire c12375;
    assign in12375_1 = {s10669[0]};
    assign in12375_2 = {s10670[0]};
    Full_Adder FA_12375(s12375, c12375, in12375_1, in12375_2, s10668[0]);
    wire[0:0] s12376, in12376_1, in12376_2;
    wire c12376;
    assign in12376_1 = {s8153[0]};
    assign in12376_2 = {c10663};
    Full_Adder FA_12376(s12376, c12376, in12376_1, in12376_2, s8152[0]);
    wire[0:0] s12377, in12377_1, in12377_2;
    wire c12377;
    assign in12377_1 = {c10665};
    assign in12377_2 = {c10666};
    Full_Adder FA_12377(s12377, c12377, in12377_1, in12377_2, c10664);
    wire[0:0] s12378, in12378_1, in12378_2;
    wire c12378;
    assign in12378_1 = {c10668};
    assign in12378_2 = {c10669};
    Full_Adder FA_12378(s12378, c12378, in12378_1, in12378_2, c10667);
    wire[0:0] s12379, in12379_1, in12379_2;
    wire c12379;
    assign in12379_1 = {s10671[0]};
    assign in12379_2 = {s10672[0]};
    Full_Adder FA_12379(s12379, c12379, in12379_1, in12379_2, c10670);
    wire[0:0] s12380, in12380_1, in12380_2;
    wire c12380;
    assign in12380_1 = {s10674[0]};
    assign in12380_2 = {s10675[0]};
    Full_Adder FA_12380(s12380, c12380, in12380_1, in12380_2, s10673[0]);
    wire[0:0] s12381, in12381_1, in12381_2;
    wire c12381;
    assign in12381_1 = {s10677[0]};
    assign in12381_2 = {s10678[0]};
    Full_Adder FA_12381(s12381, c12381, in12381_1, in12381_2, s10676[0]);
    wire[0:0] s12382, in12382_1, in12382_2;
    wire c12382;
    assign in12382_1 = {s8166[0]};
    assign in12382_2 = {c10671};
    Full_Adder FA_12382(s12382, c12382, in12382_1, in12382_2, s8165[0]);
    wire[0:0] s12383, in12383_1, in12383_2;
    wire c12383;
    assign in12383_1 = {c10673};
    assign in12383_2 = {c10674};
    Full_Adder FA_12383(s12383, c12383, in12383_1, in12383_2, c10672);
    wire[0:0] s12384, in12384_1, in12384_2;
    wire c12384;
    assign in12384_1 = {c10676};
    assign in12384_2 = {c10677};
    Full_Adder FA_12384(s12384, c12384, in12384_1, in12384_2, c10675);
    wire[0:0] s12385, in12385_1, in12385_2;
    wire c12385;
    assign in12385_1 = {s10679[0]};
    assign in12385_2 = {s10680[0]};
    Full_Adder FA_12385(s12385, c12385, in12385_1, in12385_2, c10678);
    wire[0:0] s12386, in12386_1, in12386_2;
    wire c12386;
    assign in12386_1 = {s10682[0]};
    assign in12386_2 = {s10683[0]};
    Full_Adder FA_12386(s12386, c12386, in12386_1, in12386_2, s10681[0]);
    wire[0:0] s12387, in12387_1, in12387_2;
    wire c12387;
    assign in12387_1 = {s10685[0]};
    assign in12387_2 = {s10686[0]};
    Full_Adder FA_12387(s12387, c12387, in12387_1, in12387_2, s10684[0]);
    wire[0:0] s12388, in12388_1, in12388_2;
    wire c12388;
    assign in12388_1 = {s8179[0]};
    assign in12388_2 = {c10679};
    Full_Adder FA_12388(s12388, c12388, in12388_1, in12388_2, s8178[0]);
    wire[0:0] s12389, in12389_1, in12389_2;
    wire c12389;
    assign in12389_1 = {c10681};
    assign in12389_2 = {c10682};
    Full_Adder FA_12389(s12389, c12389, in12389_1, in12389_2, c10680);
    wire[0:0] s12390, in12390_1, in12390_2;
    wire c12390;
    assign in12390_1 = {c10684};
    assign in12390_2 = {c10685};
    Full_Adder FA_12390(s12390, c12390, in12390_1, in12390_2, c10683);
    wire[0:0] s12391, in12391_1, in12391_2;
    wire c12391;
    assign in12391_1 = {s10687[0]};
    assign in12391_2 = {s10688[0]};
    Full_Adder FA_12391(s12391, c12391, in12391_1, in12391_2, c10686);
    wire[0:0] s12392, in12392_1, in12392_2;
    wire c12392;
    assign in12392_1 = {s10690[0]};
    assign in12392_2 = {s10691[0]};
    Full_Adder FA_12392(s12392, c12392, in12392_1, in12392_2, s10689[0]);
    wire[0:0] s12393, in12393_1, in12393_2;
    wire c12393;
    assign in12393_1 = {s10693[0]};
    assign in12393_2 = {s10694[0]};
    Full_Adder FA_12393(s12393, c12393, in12393_1, in12393_2, s10692[0]);
    wire[0:0] s12394, in12394_1, in12394_2;
    wire c12394;
    assign in12394_1 = {s8192[0]};
    assign in12394_2 = {c10687};
    Full_Adder FA_12394(s12394, c12394, in12394_1, in12394_2, s8191[0]);
    wire[0:0] s12395, in12395_1, in12395_2;
    wire c12395;
    assign in12395_1 = {c10689};
    assign in12395_2 = {c10690};
    Full_Adder FA_12395(s12395, c12395, in12395_1, in12395_2, c10688);
    wire[0:0] s12396, in12396_1, in12396_2;
    wire c12396;
    assign in12396_1 = {c10692};
    assign in12396_2 = {c10693};
    Full_Adder FA_12396(s12396, c12396, in12396_1, in12396_2, c10691);
    wire[0:0] s12397, in12397_1, in12397_2;
    wire c12397;
    assign in12397_1 = {s10695[0]};
    assign in12397_2 = {s10696[0]};
    Full_Adder FA_12397(s12397, c12397, in12397_1, in12397_2, c10694);
    wire[0:0] s12398, in12398_1, in12398_2;
    wire c12398;
    assign in12398_1 = {s10698[0]};
    assign in12398_2 = {s10699[0]};
    Full_Adder FA_12398(s12398, c12398, in12398_1, in12398_2, s10697[0]);
    wire[0:0] s12399, in12399_1, in12399_2;
    wire c12399;
    assign in12399_1 = {s10701[0]};
    assign in12399_2 = {s10702[0]};
    Full_Adder FA_12399(s12399, c12399, in12399_1, in12399_2, s10700[0]);
    wire[0:0] s12400, in12400_1, in12400_2;
    wire c12400;
    assign in12400_1 = {s8205[0]};
    assign in12400_2 = {c10695};
    Full_Adder FA_12400(s12400, c12400, in12400_1, in12400_2, s8204[0]);
    wire[0:0] s12401, in12401_1, in12401_2;
    wire c12401;
    assign in12401_1 = {c10697};
    assign in12401_2 = {c10698};
    Full_Adder FA_12401(s12401, c12401, in12401_1, in12401_2, c10696);
    wire[0:0] s12402, in12402_1, in12402_2;
    wire c12402;
    assign in12402_1 = {c10700};
    assign in12402_2 = {c10701};
    Full_Adder FA_12402(s12402, c12402, in12402_1, in12402_2, c10699);
    wire[0:0] s12403, in12403_1, in12403_2;
    wire c12403;
    assign in12403_1 = {s10703[0]};
    assign in12403_2 = {s10704[0]};
    Full_Adder FA_12403(s12403, c12403, in12403_1, in12403_2, c10702);
    wire[0:0] s12404, in12404_1, in12404_2;
    wire c12404;
    assign in12404_1 = {s10706[0]};
    assign in12404_2 = {s10707[0]};
    Full_Adder FA_12404(s12404, c12404, in12404_1, in12404_2, s10705[0]);
    wire[0:0] s12405, in12405_1, in12405_2;
    wire c12405;
    assign in12405_1 = {s10709[0]};
    assign in12405_2 = {s10710[0]};
    Full_Adder FA_12405(s12405, c12405, in12405_1, in12405_2, s10708[0]);
    wire[0:0] s12406, in12406_1, in12406_2;
    wire c12406;
    assign in12406_1 = {s8218[0]};
    assign in12406_2 = {c10703};
    Full_Adder FA_12406(s12406, c12406, in12406_1, in12406_2, s8217[0]);
    wire[0:0] s12407, in12407_1, in12407_2;
    wire c12407;
    assign in12407_1 = {c10705};
    assign in12407_2 = {c10706};
    Full_Adder FA_12407(s12407, c12407, in12407_1, in12407_2, c10704);
    wire[0:0] s12408, in12408_1, in12408_2;
    wire c12408;
    assign in12408_1 = {c10708};
    assign in12408_2 = {c10709};
    Full_Adder FA_12408(s12408, c12408, in12408_1, in12408_2, c10707);
    wire[0:0] s12409, in12409_1, in12409_2;
    wire c12409;
    assign in12409_1 = {s10711[0]};
    assign in12409_2 = {s10712[0]};
    Full_Adder FA_12409(s12409, c12409, in12409_1, in12409_2, c10710);
    wire[0:0] s12410, in12410_1, in12410_2;
    wire c12410;
    assign in12410_1 = {s10714[0]};
    assign in12410_2 = {s10715[0]};
    Full_Adder FA_12410(s12410, c12410, in12410_1, in12410_2, s10713[0]);
    wire[0:0] s12411, in12411_1, in12411_2;
    wire c12411;
    assign in12411_1 = {s10717[0]};
    assign in12411_2 = {s10718[0]};
    Full_Adder FA_12411(s12411, c12411, in12411_1, in12411_2, s10716[0]);
    wire[0:0] s12412, in12412_1, in12412_2;
    wire c12412;
    assign in12412_1 = {s8231[0]};
    assign in12412_2 = {c10711};
    Full_Adder FA_12412(s12412, c12412, in12412_1, in12412_2, s8230[0]);
    wire[0:0] s12413, in12413_1, in12413_2;
    wire c12413;
    assign in12413_1 = {c10713};
    assign in12413_2 = {c10714};
    Full_Adder FA_12413(s12413, c12413, in12413_1, in12413_2, c10712);
    wire[0:0] s12414, in12414_1, in12414_2;
    wire c12414;
    assign in12414_1 = {c10716};
    assign in12414_2 = {c10717};
    Full_Adder FA_12414(s12414, c12414, in12414_1, in12414_2, c10715);
    wire[0:0] s12415, in12415_1, in12415_2;
    wire c12415;
    assign in12415_1 = {s10719[0]};
    assign in12415_2 = {s10720[0]};
    Full_Adder FA_12415(s12415, c12415, in12415_1, in12415_2, c10718);
    wire[0:0] s12416, in12416_1, in12416_2;
    wire c12416;
    assign in12416_1 = {s10722[0]};
    assign in12416_2 = {s10723[0]};
    Full_Adder FA_12416(s12416, c12416, in12416_1, in12416_2, s10721[0]);
    wire[0:0] s12417, in12417_1, in12417_2;
    wire c12417;
    assign in12417_1 = {s10725[0]};
    assign in12417_2 = {s10726[0]};
    Full_Adder FA_12417(s12417, c12417, in12417_1, in12417_2, s10724[0]);
    wire[0:0] s12418, in12418_1, in12418_2;
    wire c12418;
    assign in12418_1 = {s8244[0]};
    assign in12418_2 = {c10719};
    Full_Adder FA_12418(s12418, c12418, in12418_1, in12418_2, s8243[0]);
    wire[0:0] s12419, in12419_1, in12419_2;
    wire c12419;
    assign in12419_1 = {c10721};
    assign in12419_2 = {c10722};
    Full_Adder FA_12419(s12419, c12419, in12419_1, in12419_2, c10720);
    wire[0:0] s12420, in12420_1, in12420_2;
    wire c12420;
    assign in12420_1 = {c10724};
    assign in12420_2 = {c10725};
    Full_Adder FA_12420(s12420, c12420, in12420_1, in12420_2, c10723);
    wire[0:0] s12421, in12421_1, in12421_2;
    wire c12421;
    assign in12421_1 = {s10727[0]};
    assign in12421_2 = {s10728[0]};
    Full_Adder FA_12421(s12421, c12421, in12421_1, in12421_2, c10726);
    wire[0:0] s12422, in12422_1, in12422_2;
    wire c12422;
    assign in12422_1 = {s10730[0]};
    assign in12422_2 = {s10731[0]};
    Full_Adder FA_12422(s12422, c12422, in12422_1, in12422_2, s10729[0]);
    wire[0:0] s12423, in12423_1, in12423_2;
    wire c12423;
    assign in12423_1 = {s10733[0]};
    assign in12423_2 = {s10734[0]};
    Full_Adder FA_12423(s12423, c12423, in12423_1, in12423_2, s10732[0]);
    wire[0:0] s12424, in12424_1, in12424_2;
    wire c12424;
    assign in12424_1 = {s8257[0]};
    assign in12424_2 = {c10727};
    Full_Adder FA_12424(s12424, c12424, in12424_1, in12424_2, s8256[0]);
    wire[0:0] s12425, in12425_1, in12425_2;
    wire c12425;
    assign in12425_1 = {c10729};
    assign in12425_2 = {c10730};
    Full_Adder FA_12425(s12425, c12425, in12425_1, in12425_2, c10728);
    wire[0:0] s12426, in12426_1, in12426_2;
    wire c12426;
    assign in12426_1 = {c10732};
    assign in12426_2 = {c10733};
    Full_Adder FA_12426(s12426, c12426, in12426_1, in12426_2, c10731);
    wire[0:0] s12427, in12427_1, in12427_2;
    wire c12427;
    assign in12427_1 = {s10735[0]};
    assign in12427_2 = {s10736[0]};
    Full_Adder FA_12427(s12427, c12427, in12427_1, in12427_2, c10734);
    wire[0:0] s12428, in12428_1, in12428_2;
    wire c12428;
    assign in12428_1 = {s10738[0]};
    assign in12428_2 = {s10739[0]};
    Full_Adder FA_12428(s12428, c12428, in12428_1, in12428_2, s10737[0]);
    wire[0:0] s12429, in12429_1, in12429_2;
    wire c12429;
    assign in12429_1 = {s10741[0]};
    assign in12429_2 = {s10742[0]};
    Full_Adder FA_12429(s12429, c12429, in12429_1, in12429_2, s10740[0]);
    wire[0:0] s12430, in12430_1, in12430_2;
    wire c12430;
    assign in12430_1 = {s8270[0]};
    assign in12430_2 = {c10735};
    Full_Adder FA_12430(s12430, c12430, in12430_1, in12430_2, s8269[0]);
    wire[0:0] s12431, in12431_1, in12431_2;
    wire c12431;
    assign in12431_1 = {c10737};
    assign in12431_2 = {c10738};
    Full_Adder FA_12431(s12431, c12431, in12431_1, in12431_2, c10736);
    wire[0:0] s12432, in12432_1, in12432_2;
    wire c12432;
    assign in12432_1 = {c10740};
    assign in12432_2 = {c10741};
    Full_Adder FA_12432(s12432, c12432, in12432_1, in12432_2, c10739);
    wire[0:0] s12433, in12433_1, in12433_2;
    wire c12433;
    assign in12433_1 = {s10743[0]};
    assign in12433_2 = {s10744[0]};
    Full_Adder FA_12433(s12433, c12433, in12433_1, in12433_2, c10742);
    wire[0:0] s12434, in12434_1, in12434_2;
    wire c12434;
    assign in12434_1 = {s10746[0]};
    assign in12434_2 = {s10747[0]};
    Full_Adder FA_12434(s12434, c12434, in12434_1, in12434_2, s10745[0]);
    wire[0:0] s12435, in12435_1, in12435_2;
    wire c12435;
    assign in12435_1 = {s10749[0]};
    assign in12435_2 = {s10750[0]};
    Full_Adder FA_12435(s12435, c12435, in12435_1, in12435_2, s10748[0]);
    wire[0:0] s12436, in12436_1, in12436_2;
    wire c12436;
    assign in12436_1 = {s8283[0]};
    assign in12436_2 = {c10743};
    Full_Adder FA_12436(s12436, c12436, in12436_1, in12436_2, s8282[0]);
    wire[0:0] s12437, in12437_1, in12437_2;
    wire c12437;
    assign in12437_1 = {c10745};
    assign in12437_2 = {c10746};
    Full_Adder FA_12437(s12437, c12437, in12437_1, in12437_2, c10744);
    wire[0:0] s12438, in12438_1, in12438_2;
    wire c12438;
    assign in12438_1 = {c10748};
    assign in12438_2 = {c10749};
    Full_Adder FA_12438(s12438, c12438, in12438_1, in12438_2, c10747);
    wire[0:0] s12439, in12439_1, in12439_2;
    wire c12439;
    assign in12439_1 = {s10751[0]};
    assign in12439_2 = {s10752[0]};
    Full_Adder FA_12439(s12439, c12439, in12439_1, in12439_2, c10750);
    wire[0:0] s12440, in12440_1, in12440_2;
    wire c12440;
    assign in12440_1 = {s10754[0]};
    assign in12440_2 = {s10755[0]};
    Full_Adder FA_12440(s12440, c12440, in12440_1, in12440_2, s10753[0]);
    wire[0:0] s12441, in12441_1, in12441_2;
    wire c12441;
    assign in12441_1 = {s10757[0]};
    assign in12441_2 = {s10758[0]};
    Full_Adder FA_12441(s12441, c12441, in12441_1, in12441_2, s10756[0]);
    wire[0:0] s12442, in12442_1, in12442_2;
    wire c12442;
    assign in12442_1 = {s8296[0]};
    assign in12442_2 = {c10751};
    Full_Adder FA_12442(s12442, c12442, in12442_1, in12442_2, s8295[0]);
    wire[0:0] s12443, in12443_1, in12443_2;
    wire c12443;
    assign in12443_1 = {c10753};
    assign in12443_2 = {c10754};
    Full_Adder FA_12443(s12443, c12443, in12443_1, in12443_2, c10752);
    wire[0:0] s12444, in12444_1, in12444_2;
    wire c12444;
    assign in12444_1 = {c10756};
    assign in12444_2 = {c10757};
    Full_Adder FA_12444(s12444, c12444, in12444_1, in12444_2, c10755);
    wire[0:0] s12445, in12445_1, in12445_2;
    wire c12445;
    assign in12445_1 = {s10759[0]};
    assign in12445_2 = {s10760[0]};
    Full_Adder FA_12445(s12445, c12445, in12445_1, in12445_2, c10758);
    wire[0:0] s12446, in12446_1, in12446_2;
    wire c12446;
    assign in12446_1 = {s10762[0]};
    assign in12446_2 = {s10763[0]};
    Full_Adder FA_12446(s12446, c12446, in12446_1, in12446_2, s10761[0]);
    wire[0:0] s12447, in12447_1, in12447_2;
    wire c12447;
    assign in12447_1 = {s10765[0]};
    assign in12447_2 = {s10766[0]};
    Full_Adder FA_12447(s12447, c12447, in12447_1, in12447_2, s10764[0]);
    wire[0:0] s12448, in12448_1, in12448_2;
    wire c12448;
    assign in12448_1 = {s8309[0]};
    assign in12448_2 = {c10759};
    Full_Adder FA_12448(s12448, c12448, in12448_1, in12448_2, s8308[0]);
    wire[0:0] s12449, in12449_1, in12449_2;
    wire c12449;
    assign in12449_1 = {c10761};
    assign in12449_2 = {c10762};
    Full_Adder FA_12449(s12449, c12449, in12449_1, in12449_2, c10760);
    wire[0:0] s12450, in12450_1, in12450_2;
    wire c12450;
    assign in12450_1 = {c10764};
    assign in12450_2 = {c10765};
    Full_Adder FA_12450(s12450, c12450, in12450_1, in12450_2, c10763);
    wire[0:0] s12451, in12451_1, in12451_2;
    wire c12451;
    assign in12451_1 = {s10767[0]};
    assign in12451_2 = {s10768[0]};
    Full_Adder FA_12451(s12451, c12451, in12451_1, in12451_2, c10766);
    wire[0:0] s12452, in12452_1, in12452_2;
    wire c12452;
    assign in12452_1 = {s10770[0]};
    assign in12452_2 = {s10771[0]};
    Full_Adder FA_12452(s12452, c12452, in12452_1, in12452_2, s10769[0]);
    wire[0:0] s12453, in12453_1, in12453_2;
    wire c12453;
    assign in12453_1 = {s10773[0]};
    assign in12453_2 = {s10774[0]};
    Full_Adder FA_12453(s12453, c12453, in12453_1, in12453_2, s10772[0]);
    wire[0:0] s12454, in12454_1, in12454_2;
    wire c12454;
    assign in12454_1 = {s8322[0]};
    assign in12454_2 = {c10767};
    Full_Adder FA_12454(s12454, c12454, in12454_1, in12454_2, s8321[0]);
    wire[0:0] s12455, in12455_1, in12455_2;
    wire c12455;
    assign in12455_1 = {c10769};
    assign in12455_2 = {c10770};
    Full_Adder FA_12455(s12455, c12455, in12455_1, in12455_2, c10768);
    wire[0:0] s12456, in12456_1, in12456_2;
    wire c12456;
    assign in12456_1 = {c10772};
    assign in12456_2 = {c10773};
    Full_Adder FA_12456(s12456, c12456, in12456_1, in12456_2, c10771);
    wire[0:0] s12457, in12457_1, in12457_2;
    wire c12457;
    assign in12457_1 = {s10775[0]};
    assign in12457_2 = {s10776[0]};
    Full_Adder FA_12457(s12457, c12457, in12457_1, in12457_2, c10774);
    wire[0:0] s12458, in12458_1, in12458_2;
    wire c12458;
    assign in12458_1 = {s10778[0]};
    assign in12458_2 = {s10779[0]};
    Full_Adder FA_12458(s12458, c12458, in12458_1, in12458_2, s10777[0]);
    wire[0:0] s12459, in12459_1, in12459_2;
    wire c12459;
    assign in12459_1 = {s10781[0]};
    assign in12459_2 = {s10782[0]};
    Full_Adder FA_12459(s12459, c12459, in12459_1, in12459_2, s10780[0]);
    wire[0:0] s12460, in12460_1, in12460_2;
    wire c12460;
    assign in12460_1 = {s8335[0]};
    assign in12460_2 = {c10775};
    Full_Adder FA_12460(s12460, c12460, in12460_1, in12460_2, s8334[0]);
    wire[0:0] s12461, in12461_1, in12461_2;
    wire c12461;
    assign in12461_1 = {c10777};
    assign in12461_2 = {c10778};
    Full_Adder FA_12461(s12461, c12461, in12461_1, in12461_2, c10776);
    wire[0:0] s12462, in12462_1, in12462_2;
    wire c12462;
    assign in12462_1 = {c10780};
    assign in12462_2 = {c10781};
    Full_Adder FA_12462(s12462, c12462, in12462_1, in12462_2, c10779);
    wire[0:0] s12463, in12463_1, in12463_2;
    wire c12463;
    assign in12463_1 = {s10783[0]};
    assign in12463_2 = {s10784[0]};
    Full_Adder FA_12463(s12463, c12463, in12463_1, in12463_2, c10782);
    wire[0:0] s12464, in12464_1, in12464_2;
    wire c12464;
    assign in12464_1 = {s10786[0]};
    assign in12464_2 = {s10787[0]};
    Full_Adder FA_12464(s12464, c12464, in12464_1, in12464_2, s10785[0]);
    wire[0:0] s12465, in12465_1, in12465_2;
    wire c12465;
    assign in12465_1 = {s10789[0]};
    assign in12465_2 = {s10790[0]};
    Full_Adder FA_12465(s12465, c12465, in12465_1, in12465_2, s10788[0]);
    wire[0:0] s12466, in12466_1, in12466_2;
    wire c12466;
    assign in12466_1 = {s8348[0]};
    assign in12466_2 = {c10783};
    Full_Adder FA_12466(s12466, c12466, in12466_1, in12466_2, s8347[0]);
    wire[0:0] s12467, in12467_1, in12467_2;
    wire c12467;
    assign in12467_1 = {c10785};
    assign in12467_2 = {c10786};
    Full_Adder FA_12467(s12467, c12467, in12467_1, in12467_2, c10784);
    wire[0:0] s12468, in12468_1, in12468_2;
    wire c12468;
    assign in12468_1 = {c10788};
    assign in12468_2 = {c10789};
    Full_Adder FA_12468(s12468, c12468, in12468_1, in12468_2, c10787);
    wire[0:0] s12469, in12469_1, in12469_2;
    wire c12469;
    assign in12469_1 = {s10791[0]};
    assign in12469_2 = {s10792[0]};
    Full_Adder FA_12469(s12469, c12469, in12469_1, in12469_2, c10790);
    wire[0:0] s12470, in12470_1, in12470_2;
    wire c12470;
    assign in12470_1 = {s10794[0]};
    assign in12470_2 = {s10795[0]};
    Full_Adder FA_12470(s12470, c12470, in12470_1, in12470_2, s10793[0]);
    wire[0:0] s12471, in12471_1, in12471_2;
    wire c12471;
    assign in12471_1 = {s10797[0]};
    assign in12471_2 = {s10798[0]};
    Full_Adder FA_12471(s12471, c12471, in12471_1, in12471_2, s10796[0]);
    wire[0:0] s12472, in12472_1, in12472_2;
    wire c12472;
    assign in12472_1 = {s8361[0]};
    assign in12472_2 = {c10791};
    Full_Adder FA_12472(s12472, c12472, in12472_1, in12472_2, s8360[0]);
    wire[0:0] s12473, in12473_1, in12473_2;
    wire c12473;
    assign in12473_1 = {c10793};
    assign in12473_2 = {c10794};
    Full_Adder FA_12473(s12473, c12473, in12473_1, in12473_2, c10792);
    wire[0:0] s12474, in12474_1, in12474_2;
    wire c12474;
    assign in12474_1 = {c10796};
    assign in12474_2 = {c10797};
    Full_Adder FA_12474(s12474, c12474, in12474_1, in12474_2, c10795);
    wire[0:0] s12475, in12475_1, in12475_2;
    wire c12475;
    assign in12475_1 = {s10799[0]};
    assign in12475_2 = {s10800[0]};
    Full_Adder FA_12475(s12475, c12475, in12475_1, in12475_2, c10798);
    wire[0:0] s12476, in12476_1, in12476_2;
    wire c12476;
    assign in12476_1 = {s10802[0]};
    assign in12476_2 = {s10803[0]};
    Full_Adder FA_12476(s12476, c12476, in12476_1, in12476_2, s10801[0]);
    wire[0:0] s12477, in12477_1, in12477_2;
    wire c12477;
    assign in12477_1 = {s10805[0]};
    assign in12477_2 = {s10806[0]};
    Full_Adder FA_12477(s12477, c12477, in12477_1, in12477_2, s10804[0]);
    wire[0:0] s12478, in12478_1, in12478_2;
    wire c12478;
    assign in12478_1 = {s8374[0]};
    assign in12478_2 = {c10799};
    Full_Adder FA_12478(s12478, c12478, in12478_1, in12478_2, s8373[0]);
    wire[0:0] s12479, in12479_1, in12479_2;
    wire c12479;
    assign in12479_1 = {c10801};
    assign in12479_2 = {c10802};
    Full_Adder FA_12479(s12479, c12479, in12479_1, in12479_2, c10800);
    wire[0:0] s12480, in12480_1, in12480_2;
    wire c12480;
    assign in12480_1 = {c10804};
    assign in12480_2 = {c10805};
    Full_Adder FA_12480(s12480, c12480, in12480_1, in12480_2, c10803);
    wire[0:0] s12481, in12481_1, in12481_2;
    wire c12481;
    assign in12481_1 = {s10807[0]};
    assign in12481_2 = {s10808[0]};
    Full_Adder FA_12481(s12481, c12481, in12481_1, in12481_2, c10806);
    wire[0:0] s12482, in12482_1, in12482_2;
    wire c12482;
    assign in12482_1 = {s10810[0]};
    assign in12482_2 = {s10811[0]};
    Full_Adder FA_12482(s12482, c12482, in12482_1, in12482_2, s10809[0]);
    wire[0:0] s12483, in12483_1, in12483_2;
    wire c12483;
    assign in12483_1 = {s10813[0]};
    assign in12483_2 = {s10814[0]};
    Full_Adder FA_12483(s12483, c12483, in12483_1, in12483_2, s10812[0]);
    wire[0:0] s12484, in12484_1, in12484_2;
    wire c12484;
    assign in12484_1 = {s8387[0]};
    assign in12484_2 = {c10807};
    Full_Adder FA_12484(s12484, c12484, in12484_1, in12484_2, s8386[0]);
    wire[0:0] s12485, in12485_1, in12485_2;
    wire c12485;
    assign in12485_1 = {c10809};
    assign in12485_2 = {c10810};
    Full_Adder FA_12485(s12485, c12485, in12485_1, in12485_2, c10808);
    wire[0:0] s12486, in12486_1, in12486_2;
    wire c12486;
    assign in12486_1 = {c10812};
    assign in12486_2 = {c10813};
    Full_Adder FA_12486(s12486, c12486, in12486_1, in12486_2, c10811);
    wire[0:0] s12487, in12487_1, in12487_2;
    wire c12487;
    assign in12487_1 = {s10815[0]};
    assign in12487_2 = {s10816[0]};
    Full_Adder FA_12487(s12487, c12487, in12487_1, in12487_2, c10814);
    wire[0:0] s12488, in12488_1, in12488_2;
    wire c12488;
    assign in12488_1 = {s10818[0]};
    assign in12488_2 = {s10819[0]};
    Full_Adder FA_12488(s12488, c12488, in12488_1, in12488_2, s10817[0]);
    wire[0:0] s12489, in12489_1, in12489_2;
    wire c12489;
    assign in12489_1 = {s10821[0]};
    assign in12489_2 = {s10822[0]};
    Full_Adder FA_12489(s12489, c12489, in12489_1, in12489_2, s10820[0]);
    wire[0:0] s12490, in12490_1, in12490_2;
    wire c12490;
    assign in12490_1 = {s8400[0]};
    assign in12490_2 = {c10815};
    Full_Adder FA_12490(s12490, c12490, in12490_1, in12490_2, s8399[0]);
    wire[0:0] s12491, in12491_1, in12491_2;
    wire c12491;
    assign in12491_1 = {c10817};
    assign in12491_2 = {c10818};
    Full_Adder FA_12491(s12491, c12491, in12491_1, in12491_2, c10816);
    wire[0:0] s12492, in12492_1, in12492_2;
    wire c12492;
    assign in12492_1 = {c10820};
    assign in12492_2 = {c10821};
    Full_Adder FA_12492(s12492, c12492, in12492_1, in12492_2, c10819);
    wire[0:0] s12493, in12493_1, in12493_2;
    wire c12493;
    assign in12493_1 = {s10823[0]};
    assign in12493_2 = {s10824[0]};
    Full_Adder FA_12493(s12493, c12493, in12493_1, in12493_2, c10822);
    wire[0:0] s12494, in12494_1, in12494_2;
    wire c12494;
    assign in12494_1 = {s10826[0]};
    assign in12494_2 = {s10827[0]};
    Full_Adder FA_12494(s12494, c12494, in12494_1, in12494_2, s10825[0]);
    wire[0:0] s12495, in12495_1, in12495_2;
    wire c12495;
    assign in12495_1 = {s10829[0]};
    assign in12495_2 = {s10830[0]};
    Full_Adder FA_12495(s12495, c12495, in12495_1, in12495_2, s10828[0]);
    wire[0:0] s12496, in12496_1, in12496_2;
    wire c12496;
    assign in12496_1 = {s8413[0]};
    assign in12496_2 = {c10823};
    Full_Adder FA_12496(s12496, c12496, in12496_1, in12496_2, s8412[0]);
    wire[0:0] s12497, in12497_1, in12497_2;
    wire c12497;
    assign in12497_1 = {c10825};
    assign in12497_2 = {c10826};
    Full_Adder FA_12497(s12497, c12497, in12497_1, in12497_2, c10824);
    wire[0:0] s12498, in12498_1, in12498_2;
    wire c12498;
    assign in12498_1 = {c10828};
    assign in12498_2 = {c10829};
    Full_Adder FA_12498(s12498, c12498, in12498_1, in12498_2, c10827);
    wire[0:0] s12499, in12499_1, in12499_2;
    wire c12499;
    assign in12499_1 = {s10831[0]};
    assign in12499_2 = {s10832[0]};
    Full_Adder FA_12499(s12499, c12499, in12499_1, in12499_2, c10830);
    wire[0:0] s12500, in12500_1, in12500_2;
    wire c12500;
    assign in12500_1 = {s10834[0]};
    assign in12500_2 = {s10835[0]};
    Full_Adder FA_12500(s12500, c12500, in12500_1, in12500_2, s10833[0]);
    wire[0:0] s12501, in12501_1, in12501_2;
    wire c12501;
    assign in12501_1 = {s10837[0]};
    assign in12501_2 = {s10838[0]};
    Full_Adder FA_12501(s12501, c12501, in12501_1, in12501_2, s10836[0]);
    wire[0:0] s12502, in12502_1, in12502_2;
    wire c12502;
    assign in12502_1 = {s8426[0]};
    assign in12502_2 = {c10831};
    Full_Adder FA_12502(s12502, c12502, in12502_1, in12502_2, s8425[0]);
    wire[0:0] s12503, in12503_1, in12503_2;
    wire c12503;
    assign in12503_1 = {c10833};
    assign in12503_2 = {c10834};
    Full_Adder FA_12503(s12503, c12503, in12503_1, in12503_2, c10832);
    wire[0:0] s12504, in12504_1, in12504_2;
    wire c12504;
    assign in12504_1 = {c10836};
    assign in12504_2 = {c10837};
    Full_Adder FA_12504(s12504, c12504, in12504_1, in12504_2, c10835);
    wire[0:0] s12505, in12505_1, in12505_2;
    wire c12505;
    assign in12505_1 = {s10839[0]};
    assign in12505_2 = {s10840[0]};
    Full_Adder FA_12505(s12505, c12505, in12505_1, in12505_2, c10838);
    wire[0:0] s12506, in12506_1, in12506_2;
    wire c12506;
    assign in12506_1 = {s10842[0]};
    assign in12506_2 = {s10843[0]};
    Full_Adder FA_12506(s12506, c12506, in12506_1, in12506_2, s10841[0]);
    wire[0:0] s12507, in12507_1, in12507_2;
    wire c12507;
    assign in12507_1 = {s10845[0]};
    assign in12507_2 = {s10846[0]};
    Full_Adder FA_12507(s12507, c12507, in12507_1, in12507_2, s10844[0]);
    wire[0:0] s12508, in12508_1, in12508_2;
    wire c12508;
    assign in12508_1 = {s8439[0]};
    assign in12508_2 = {c10839};
    Full_Adder FA_12508(s12508, c12508, in12508_1, in12508_2, s8438[0]);
    wire[0:0] s12509, in12509_1, in12509_2;
    wire c12509;
    assign in12509_1 = {c10841};
    assign in12509_2 = {c10842};
    Full_Adder FA_12509(s12509, c12509, in12509_1, in12509_2, c10840);
    wire[0:0] s12510, in12510_1, in12510_2;
    wire c12510;
    assign in12510_1 = {c10844};
    assign in12510_2 = {c10845};
    Full_Adder FA_12510(s12510, c12510, in12510_1, in12510_2, c10843);
    wire[0:0] s12511, in12511_1, in12511_2;
    wire c12511;
    assign in12511_1 = {s10847[0]};
    assign in12511_2 = {s10848[0]};
    Full_Adder FA_12511(s12511, c12511, in12511_1, in12511_2, c10846);
    wire[0:0] s12512, in12512_1, in12512_2;
    wire c12512;
    assign in12512_1 = {s10850[0]};
    assign in12512_2 = {s10851[0]};
    Full_Adder FA_12512(s12512, c12512, in12512_1, in12512_2, s10849[0]);
    wire[0:0] s12513, in12513_1, in12513_2;
    wire c12513;
    assign in12513_1 = {s10853[0]};
    assign in12513_2 = {s10854[0]};
    Full_Adder FA_12513(s12513, c12513, in12513_1, in12513_2, s10852[0]);
    wire[0:0] s12514, in12514_1, in12514_2;
    wire c12514;
    assign in12514_1 = {s8452[0]};
    assign in12514_2 = {c10847};
    Full_Adder FA_12514(s12514, c12514, in12514_1, in12514_2, s8451[0]);
    wire[0:0] s12515, in12515_1, in12515_2;
    wire c12515;
    assign in12515_1 = {c10849};
    assign in12515_2 = {c10850};
    Full_Adder FA_12515(s12515, c12515, in12515_1, in12515_2, c10848);
    wire[0:0] s12516, in12516_1, in12516_2;
    wire c12516;
    assign in12516_1 = {c10852};
    assign in12516_2 = {c10853};
    Full_Adder FA_12516(s12516, c12516, in12516_1, in12516_2, c10851);
    wire[0:0] s12517, in12517_1, in12517_2;
    wire c12517;
    assign in12517_1 = {s10855[0]};
    assign in12517_2 = {s10856[0]};
    Full_Adder FA_12517(s12517, c12517, in12517_1, in12517_2, c10854);
    wire[0:0] s12518, in12518_1, in12518_2;
    wire c12518;
    assign in12518_1 = {s10858[0]};
    assign in12518_2 = {s10859[0]};
    Full_Adder FA_12518(s12518, c12518, in12518_1, in12518_2, s10857[0]);
    wire[0:0] s12519, in12519_1, in12519_2;
    wire c12519;
    assign in12519_1 = {s10861[0]};
    assign in12519_2 = {s10862[0]};
    Full_Adder FA_12519(s12519, c12519, in12519_1, in12519_2, s10860[0]);
    wire[0:0] s12520, in12520_1, in12520_2;
    wire c12520;
    assign in12520_1 = {s8465[0]};
    assign in12520_2 = {c10855};
    Full_Adder FA_12520(s12520, c12520, in12520_1, in12520_2, s8464[0]);
    wire[0:0] s12521, in12521_1, in12521_2;
    wire c12521;
    assign in12521_1 = {c10857};
    assign in12521_2 = {c10858};
    Full_Adder FA_12521(s12521, c12521, in12521_1, in12521_2, c10856);
    wire[0:0] s12522, in12522_1, in12522_2;
    wire c12522;
    assign in12522_1 = {c10860};
    assign in12522_2 = {c10861};
    Full_Adder FA_12522(s12522, c12522, in12522_1, in12522_2, c10859);
    wire[0:0] s12523, in12523_1, in12523_2;
    wire c12523;
    assign in12523_1 = {s10863[0]};
    assign in12523_2 = {s10864[0]};
    Full_Adder FA_12523(s12523, c12523, in12523_1, in12523_2, c10862);
    wire[0:0] s12524, in12524_1, in12524_2;
    wire c12524;
    assign in12524_1 = {s10866[0]};
    assign in12524_2 = {s10867[0]};
    Full_Adder FA_12524(s12524, c12524, in12524_1, in12524_2, s10865[0]);
    wire[0:0] s12525, in12525_1, in12525_2;
    wire c12525;
    assign in12525_1 = {s10869[0]};
    assign in12525_2 = {s10870[0]};
    Full_Adder FA_12525(s12525, c12525, in12525_1, in12525_2, s10868[0]);
    wire[0:0] s12526, in12526_1, in12526_2;
    wire c12526;
    assign in12526_1 = {s8478[0]};
    assign in12526_2 = {c10863};
    Full_Adder FA_12526(s12526, c12526, in12526_1, in12526_2, s8477[0]);
    wire[0:0] s12527, in12527_1, in12527_2;
    wire c12527;
    assign in12527_1 = {c10865};
    assign in12527_2 = {c10866};
    Full_Adder FA_12527(s12527, c12527, in12527_1, in12527_2, c10864);
    wire[0:0] s12528, in12528_1, in12528_2;
    wire c12528;
    assign in12528_1 = {c10868};
    assign in12528_2 = {c10869};
    Full_Adder FA_12528(s12528, c12528, in12528_1, in12528_2, c10867);
    wire[0:0] s12529, in12529_1, in12529_2;
    wire c12529;
    assign in12529_1 = {s10871[0]};
    assign in12529_2 = {s10872[0]};
    Full_Adder FA_12529(s12529, c12529, in12529_1, in12529_2, c10870);
    wire[0:0] s12530, in12530_1, in12530_2;
    wire c12530;
    assign in12530_1 = {s10874[0]};
    assign in12530_2 = {s10875[0]};
    Full_Adder FA_12530(s12530, c12530, in12530_1, in12530_2, s10873[0]);
    wire[0:0] s12531, in12531_1, in12531_2;
    wire c12531;
    assign in12531_1 = {s10877[0]};
    assign in12531_2 = {s10878[0]};
    Full_Adder FA_12531(s12531, c12531, in12531_1, in12531_2, s10876[0]);
    wire[0:0] s12532, in12532_1, in12532_2;
    wire c12532;
    assign in12532_1 = {s8491[0]};
    assign in12532_2 = {c10871};
    Full_Adder FA_12532(s12532, c12532, in12532_1, in12532_2, s8490[0]);
    wire[0:0] s12533, in12533_1, in12533_2;
    wire c12533;
    assign in12533_1 = {c10873};
    assign in12533_2 = {c10874};
    Full_Adder FA_12533(s12533, c12533, in12533_1, in12533_2, c10872);
    wire[0:0] s12534, in12534_1, in12534_2;
    wire c12534;
    assign in12534_1 = {c10876};
    assign in12534_2 = {c10877};
    Full_Adder FA_12534(s12534, c12534, in12534_1, in12534_2, c10875);
    wire[0:0] s12535, in12535_1, in12535_2;
    wire c12535;
    assign in12535_1 = {s10879[0]};
    assign in12535_2 = {s10880[0]};
    Full_Adder FA_12535(s12535, c12535, in12535_1, in12535_2, c10878);
    wire[0:0] s12536, in12536_1, in12536_2;
    wire c12536;
    assign in12536_1 = {s10882[0]};
    assign in12536_2 = {s10883[0]};
    Full_Adder FA_12536(s12536, c12536, in12536_1, in12536_2, s10881[0]);
    wire[0:0] s12537, in12537_1, in12537_2;
    wire c12537;
    assign in12537_1 = {s10885[0]};
    assign in12537_2 = {s10886[0]};
    Full_Adder FA_12537(s12537, c12537, in12537_1, in12537_2, s10884[0]);
    wire[0:0] s12538, in12538_1, in12538_2;
    wire c12538;
    assign in12538_1 = {s8504[0]};
    assign in12538_2 = {c10879};
    Full_Adder FA_12538(s12538, c12538, in12538_1, in12538_2, s8503[0]);
    wire[0:0] s12539, in12539_1, in12539_2;
    wire c12539;
    assign in12539_1 = {c10881};
    assign in12539_2 = {c10882};
    Full_Adder FA_12539(s12539, c12539, in12539_1, in12539_2, c10880);
    wire[0:0] s12540, in12540_1, in12540_2;
    wire c12540;
    assign in12540_1 = {c10884};
    assign in12540_2 = {c10885};
    Full_Adder FA_12540(s12540, c12540, in12540_1, in12540_2, c10883);
    wire[0:0] s12541, in12541_1, in12541_2;
    wire c12541;
    assign in12541_1 = {s10887[0]};
    assign in12541_2 = {s10888[0]};
    Full_Adder FA_12541(s12541, c12541, in12541_1, in12541_2, c10886);
    wire[0:0] s12542, in12542_1, in12542_2;
    wire c12542;
    assign in12542_1 = {s10890[0]};
    assign in12542_2 = {s10891[0]};
    Full_Adder FA_12542(s12542, c12542, in12542_1, in12542_2, s10889[0]);
    wire[0:0] s12543, in12543_1, in12543_2;
    wire c12543;
    assign in12543_1 = {s10893[0]};
    assign in12543_2 = {s10894[0]};
    Full_Adder FA_12543(s12543, c12543, in12543_1, in12543_2, s10892[0]);
    wire[0:0] s12544, in12544_1, in12544_2;
    wire c12544;
    assign in12544_1 = {s8517[0]};
    assign in12544_2 = {c10887};
    Full_Adder FA_12544(s12544, c12544, in12544_1, in12544_2, s8516[0]);
    wire[0:0] s12545, in12545_1, in12545_2;
    wire c12545;
    assign in12545_1 = {c10889};
    assign in12545_2 = {c10890};
    Full_Adder FA_12545(s12545, c12545, in12545_1, in12545_2, c10888);
    wire[0:0] s12546, in12546_1, in12546_2;
    wire c12546;
    assign in12546_1 = {c10892};
    assign in12546_2 = {c10893};
    Full_Adder FA_12546(s12546, c12546, in12546_1, in12546_2, c10891);
    wire[0:0] s12547, in12547_1, in12547_2;
    wire c12547;
    assign in12547_1 = {s10895[0]};
    assign in12547_2 = {s10896[0]};
    Full_Adder FA_12547(s12547, c12547, in12547_1, in12547_2, c10894);
    wire[0:0] s12548, in12548_1, in12548_2;
    wire c12548;
    assign in12548_1 = {s10898[0]};
    assign in12548_2 = {s10899[0]};
    Full_Adder FA_12548(s12548, c12548, in12548_1, in12548_2, s10897[0]);
    wire[0:0] s12549, in12549_1, in12549_2;
    wire c12549;
    assign in12549_1 = {s10901[0]};
    assign in12549_2 = {s10902[0]};
    Full_Adder FA_12549(s12549, c12549, in12549_1, in12549_2, s10900[0]);
    wire[0:0] s12550, in12550_1, in12550_2;
    wire c12550;
    assign in12550_1 = {s8530[0]};
    assign in12550_2 = {c10895};
    Full_Adder FA_12550(s12550, c12550, in12550_1, in12550_2, s8529[0]);
    wire[0:0] s12551, in12551_1, in12551_2;
    wire c12551;
    assign in12551_1 = {c10897};
    assign in12551_2 = {c10898};
    Full_Adder FA_12551(s12551, c12551, in12551_1, in12551_2, c10896);
    wire[0:0] s12552, in12552_1, in12552_2;
    wire c12552;
    assign in12552_1 = {c10900};
    assign in12552_2 = {c10901};
    Full_Adder FA_12552(s12552, c12552, in12552_1, in12552_2, c10899);
    wire[0:0] s12553, in12553_1, in12553_2;
    wire c12553;
    assign in12553_1 = {s10903[0]};
    assign in12553_2 = {s10904[0]};
    Full_Adder FA_12553(s12553, c12553, in12553_1, in12553_2, c10902);
    wire[0:0] s12554, in12554_1, in12554_2;
    wire c12554;
    assign in12554_1 = {s10906[0]};
    assign in12554_2 = {s10907[0]};
    Full_Adder FA_12554(s12554, c12554, in12554_1, in12554_2, s10905[0]);
    wire[0:0] s12555, in12555_1, in12555_2;
    wire c12555;
    assign in12555_1 = {s10909[0]};
    assign in12555_2 = {s10910[0]};
    Full_Adder FA_12555(s12555, c12555, in12555_1, in12555_2, s10908[0]);
    wire[0:0] s12556, in12556_1, in12556_2;
    wire c12556;
    assign in12556_1 = {s8543[0]};
    assign in12556_2 = {c10903};
    Full_Adder FA_12556(s12556, c12556, in12556_1, in12556_2, s8542[0]);
    wire[0:0] s12557, in12557_1, in12557_2;
    wire c12557;
    assign in12557_1 = {c10905};
    assign in12557_2 = {c10906};
    Full_Adder FA_12557(s12557, c12557, in12557_1, in12557_2, c10904);
    wire[0:0] s12558, in12558_1, in12558_2;
    wire c12558;
    assign in12558_1 = {c10908};
    assign in12558_2 = {c10909};
    Full_Adder FA_12558(s12558, c12558, in12558_1, in12558_2, c10907);
    wire[0:0] s12559, in12559_1, in12559_2;
    wire c12559;
    assign in12559_1 = {s10911[0]};
    assign in12559_2 = {s10912[0]};
    Full_Adder FA_12559(s12559, c12559, in12559_1, in12559_2, c10910);
    wire[0:0] s12560, in12560_1, in12560_2;
    wire c12560;
    assign in12560_1 = {s10914[0]};
    assign in12560_2 = {s10915[0]};
    Full_Adder FA_12560(s12560, c12560, in12560_1, in12560_2, s10913[0]);
    wire[0:0] s12561, in12561_1, in12561_2;
    wire c12561;
    assign in12561_1 = {s10917[0]};
    assign in12561_2 = {s10918[0]};
    Full_Adder FA_12561(s12561, c12561, in12561_1, in12561_2, s10916[0]);
    wire[0:0] s12562, in12562_1, in12562_2;
    wire c12562;
    assign in12562_1 = {s8556[0]};
    assign in12562_2 = {c10911};
    Full_Adder FA_12562(s12562, c12562, in12562_1, in12562_2, s8555[0]);
    wire[0:0] s12563, in12563_1, in12563_2;
    wire c12563;
    assign in12563_1 = {c10913};
    assign in12563_2 = {c10914};
    Full_Adder FA_12563(s12563, c12563, in12563_1, in12563_2, c10912);
    wire[0:0] s12564, in12564_1, in12564_2;
    wire c12564;
    assign in12564_1 = {c10916};
    assign in12564_2 = {c10917};
    Full_Adder FA_12564(s12564, c12564, in12564_1, in12564_2, c10915);
    wire[0:0] s12565, in12565_1, in12565_2;
    wire c12565;
    assign in12565_1 = {s10919[0]};
    assign in12565_2 = {s10920[0]};
    Full_Adder FA_12565(s12565, c12565, in12565_1, in12565_2, c10918);
    wire[0:0] s12566, in12566_1, in12566_2;
    wire c12566;
    assign in12566_1 = {s10922[0]};
    assign in12566_2 = {s10923[0]};
    Full_Adder FA_12566(s12566, c12566, in12566_1, in12566_2, s10921[0]);
    wire[0:0] s12567, in12567_1, in12567_2;
    wire c12567;
    assign in12567_1 = {s10925[0]};
    assign in12567_2 = {s10926[0]};
    Full_Adder FA_12567(s12567, c12567, in12567_1, in12567_2, s10924[0]);
    wire[0:0] s12568, in12568_1, in12568_2;
    wire c12568;
    assign in12568_1 = {s8569[0]};
    assign in12568_2 = {c10919};
    Full_Adder FA_12568(s12568, c12568, in12568_1, in12568_2, s8568[0]);
    wire[0:0] s12569, in12569_1, in12569_2;
    wire c12569;
    assign in12569_1 = {c10921};
    assign in12569_2 = {c10922};
    Full_Adder FA_12569(s12569, c12569, in12569_1, in12569_2, c10920);
    wire[0:0] s12570, in12570_1, in12570_2;
    wire c12570;
    assign in12570_1 = {c10924};
    assign in12570_2 = {c10925};
    Full_Adder FA_12570(s12570, c12570, in12570_1, in12570_2, c10923);
    wire[0:0] s12571, in12571_1, in12571_2;
    wire c12571;
    assign in12571_1 = {s10927[0]};
    assign in12571_2 = {s10928[0]};
    Full_Adder FA_12571(s12571, c12571, in12571_1, in12571_2, c10926);
    wire[0:0] s12572, in12572_1, in12572_2;
    wire c12572;
    assign in12572_1 = {s10930[0]};
    assign in12572_2 = {s10931[0]};
    Full_Adder FA_12572(s12572, c12572, in12572_1, in12572_2, s10929[0]);
    wire[0:0] s12573, in12573_1, in12573_2;
    wire c12573;
    assign in12573_1 = {s10933[0]};
    assign in12573_2 = {s10934[0]};
    Full_Adder FA_12573(s12573, c12573, in12573_1, in12573_2, s10932[0]);
    wire[0:0] s12574, in12574_1, in12574_2;
    wire c12574;
    assign in12574_1 = {s8582[0]};
    assign in12574_2 = {c10927};
    Full_Adder FA_12574(s12574, c12574, in12574_1, in12574_2, s8581[0]);
    wire[0:0] s12575, in12575_1, in12575_2;
    wire c12575;
    assign in12575_1 = {c10929};
    assign in12575_2 = {c10930};
    Full_Adder FA_12575(s12575, c12575, in12575_1, in12575_2, c10928);
    wire[0:0] s12576, in12576_1, in12576_2;
    wire c12576;
    assign in12576_1 = {c10932};
    assign in12576_2 = {c10933};
    Full_Adder FA_12576(s12576, c12576, in12576_1, in12576_2, c10931);
    wire[0:0] s12577, in12577_1, in12577_2;
    wire c12577;
    assign in12577_1 = {s10935[0]};
    assign in12577_2 = {s10936[0]};
    Full_Adder FA_12577(s12577, c12577, in12577_1, in12577_2, c10934);
    wire[0:0] s12578, in12578_1, in12578_2;
    wire c12578;
    assign in12578_1 = {s10938[0]};
    assign in12578_2 = {s10939[0]};
    Full_Adder FA_12578(s12578, c12578, in12578_1, in12578_2, s10937[0]);
    wire[0:0] s12579, in12579_1, in12579_2;
    wire c12579;
    assign in12579_1 = {s10941[0]};
    assign in12579_2 = {s10942[0]};
    Full_Adder FA_12579(s12579, c12579, in12579_1, in12579_2, s10940[0]);
    wire[0:0] s12580, in12580_1, in12580_2;
    wire c12580;
    assign in12580_1 = {s8595[0]};
    assign in12580_2 = {c10935};
    Full_Adder FA_12580(s12580, c12580, in12580_1, in12580_2, s8594[0]);
    wire[0:0] s12581, in12581_1, in12581_2;
    wire c12581;
    assign in12581_1 = {c10937};
    assign in12581_2 = {c10938};
    Full_Adder FA_12581(s12581, c12581, in12581_1, in12581_2, c10936);
    wire[0:0] s12582, in12582_1, in12582_2;
    wire c12582;
    assign in12582_1 = {c10940};
    assign in12582_2 = {c10941};
    Full_Adder FA_12582(s12582, c12582, in12582_1, in12582_2, c10939);
    wire[0:0] s12583, in12583_1, in12583_2;
    wire c12583;
    assign in12583_1 = {s10943[0]};
    assign in12583_2 = {s10944[0]};
    Full_Adder FA_12583(s12583, c12583, in12583_1, in12583_2, c10942);
    wire[0:0] s12584, in12584_1, in12584_2;
    wire c12584;
    assign in12584_1 = {s10946[0]};
    assign in12584_2 = {s10947[0]};
    Full_Adder FA_12584(s12584, c12584, in12584_1, in12584_2, s10945[0]);
    wire[0:0] s12585, in12585_1, in12585_2;
    wire c12585;
    assign in12585_1 = {s10949[0]};
    assign in12585_2 = {s10950[0]};
    Full_Adder FA_12585(s12585, c12585, in12585_1, in12585_2, s10948[0]);
    wire[0:0] s12586, in12586_1, in12586_2;
    wire c12586;
    assign in12586_1 = {s8608[0]};
    assign in12586_2 = {c10943};
    Full_Adder FA_12586(s12586, c12586, in12586_1, in12586_2, s8607[0]);
    wire[0:0] s12587, in12587_1, in12587_2;
    wire c12587;
    assign in12587_1 = {c10945};
    assign in12587_2 = {c10946};
    Full_Adder FA_12587(s12587, c12587, in12587_1, in12587_2, c10944);
    wire[0:0] s12588, in12588_1, in12588_2;
    wire c12588;
    assign in12588_1 = {c10948};
    assign in12588_2 = {c10949};
    Full_Adder FA_12588(s12588, c12588, in12588_1, in12588_2, c10947);
    wire[0:0] s12589, in12589_1, in12589_2;
    wire c12589;
    assign in12589_1 = {s10951[0]};
    assign in12589_2 = {s10952[0]};
    Full_Adder FA_12589(s12589, c12589, in12589_1, in12589_2, c10950);
    wire[0:0] s12590, in12590_1, in12590_2;
    wire c12590;
    assign in12590_1 = {s10954[0]};
    assign in12590_2 = {s10955[0]};
    Full_Adder FA_12590(s12590, c12590, in12590_1, in12590_2, s10953[0]);
    wire[0:0] s12591, in12591_1, in12591_2;
    wire c12591;
    assign in12591_1 = {s10957[0]};
    assign in12591_2 = {s10958[0]};
    Full_Adder FA_12591(s12591, c12591, in12591_1, in12591_2, s10956[0]);
    wire[0:0] s12592, in12592_1, in12592_2;
    wire c12592;
    assign in12592_1 = {s8621[0]};
    assign in12592_2 = {c10951};
    Full_Adder FA_12592(s12592, c12592, in12592_1, in12592_2, s8620[0]);
    wire[0:0] s12593, in12593_1, in12593_2;
    wire c12593;
    assign in12593_1 = {c10953};
    assign in12593_2 = {c10954};
    Full_Adder FA_12593(s12593, c12593, in12593_1, in12593_2, c10952);
    wire[0:0] s12594, in12594_1, in12594_2;
    wire c12594;
    assign in12594_1 = {c10956};
    assign in12594_2 = {c10957};
    Full_Adder FA_12594(s12594, c12594, in12594_1, in12594_2, c10955);
    wire[0:0] s12595, in12595_1, in12595_2;
    wire c12595;
    assign in12595_1 = {s10959[0]};
    assign in12595_2 = {s10960[0]};
    Full_Adder FA_12595(s12595, c12595, in12595_1, in12595_2, c10958);
    wire[0:0] s12596, in12596_1, in12596_2;
    wire c12596;
    assign in12596_1 = {s10962[0]};
    assign in12596_2 = {s10963[0]};
    Full_Adder FA_12596(s12596, c12596, in12596_1, in12596_2, s10961[0]);
    wire[0:0] s12597, in12597_1, in12597_2;
    wire c12597;
    assign in12597_1 = {s10965[0]};
    assign in12597_2 = {s10966[0]};
    Full_Adder FA_12597(s12597, c12597, in12597_1, in12597_2, s10964[0]);
    wire[0:0] s12598, in12598_1, in12598_2;
    wire c12598;
    assign in12598_1 = {s8634[0]};
    assign in12598_2 = {c10959};
    Full_Adder FA_12598(s12598, c12598, in12598_1, in12598_2, s8633[0]);
    wire[0:0] s12599, in12599_1, in12599_2;
    wire c12599;
    assign in12599_1 = {c10961};
    assign in12599_2 = {c10962};
    Full_Adder FA_12599(s12599, c12599, in12599_1, in12599_2, c10960);
    wire[0:0] s12600, in12600_1, in12600_2;
    wire c12600;
    assign in12600_1 = {c10964};
    assign in12600_2 = {c10965};
    Full_Adder FA_12600(s12600, c12600, in12600_1, in12600_2, c10963);
    wire[0:0] s12601, in12601_1, in12601_2;
    wire c12601;
    assign in12601_1 = {s10967[0]};
    assign in12601_2 = {s10968[0]};
    Full_Adder FA_12601(s12601, c12601, in12601_1, in12601_2, c10966);
    wire[0:0] s12602, in12602_1, in12602_2;
    wire c12602;
    assign in12602_1 = {s10970[0]};
    assign in12602_2 = {s10971[0]};
    Full_Adder FA_12602(s12602, c12602, in12602_1, in12602_2, s10969[0]);
    wire[0:0] s12603, in12603_1, in12603_2;
    wire c12603;
    assign in12603_1 = {s10973[0]};
    assign in12603_2 = {s10974[0]};
    Full_Adder FA_12603(s12603, c12603, in12603_1, in12603_2, s10972[0]);
    wire[0:0] s12604, in12604_1, in12604_2;
    wire c12604;
    assign in12604_1 = {s8647[0]};
    assign in12604_2 = {c10967};
    Full_Adder FA_12604(s12604, c12604, in12604_1, in12604_2, s8646[0]);
    wire[0:0] s12605, in12605_1, in12605_2;
    wire c12605;
    assign in12605_1 = {c10969};
    assign in12605_2 = {c10970};
    Full_Adder FA_12605(s12605, c12605, in12605_1, in12605_2, c10968);
    wire[0:0] s12606, in12606_1, in12606_2;
    wire c12606;
    assign in12606_1 = {c10972};
    assign in12606_2 = {c10973};
    Full_Adder FA_12606(s12606, c12606, in12606_1, in12606_2, c10971);
    wire[0:0] s12607, in12607_1, in12607_2;
    wire c12607;
    assign in12607_1 = {s10975[0]};
    assign in12607_2 = {s10976[0]};
    Full_Adder FA_12607(s12607, c12607, in12607_1, in12607_2, c10974);
    wire[0:0] s12608, in12608_1, in12608_2;
    wire c12608;
    assign in12608_1 = {s10978[0]};
    assign in12608_2 = {s10979[0]};
    Full_Adder FA_12608(s12608, c12608, in12608_1, in12608_2, s10977[0]);
    wire[0:0] s12609, in12609_1, in12609_2;
    wire c12609;
    assign in12609_1 = {s10981[0]};
    assign in12609_2 = {s10982[0]};
    Full_Adder FA_12609(s12609, c12609, in12609_1, in12609_2, s10980[0]);
    wire[0:0] s12610, in12610_1, in12610_2;
    wire c12610;
    assign in12610_1 = {s8660[0]};
    assign in12610_2 = {c10975};
    Full_Adder FA_12610(s12610, c12610, in12610_1, in12610_2, s8659[0]);
    wire[0:0] s12611, in12611_1, in12611_2;
    wire c12611;
    assign in12611_1 = {c10977};
    assign in12611_2 = {c10978};
    Full_Adder FA_12611(s12611, c12611, in12611_1, in12611_2, c10976);
    wire[0:0] s12612, in12612_1, in12612_2;
    wire c12612;
    assign in12612_1 = {c10980};
    assign in12612_2 = {c10981};
    Full_Adder FA_12612(s12612, c12612, in12612_1, in12612_2, c10979);
    wire[0:0] s12613, in12613_1, in12613_2;
    wire c12613;
    assign in12613_1 = {s10983[0]};
    assign in12613_2 = {s10984[0]};
    Full_Adder FA_12613(s12613, c12613, in12613_1, in12613_2, c10982);
    wire[0:0] s12614, in12614_1, in12614_2;
    wire c12614;
    assign in12614_1 = {s10986[0]};
    assign in12614_2 = {s10987[0]};
    Full_Adder FA_12614(s12614, c12614, in12614_1, in12614_2, s10985[0]);
    wire[0:0] s12615, in12615_1, in12615_2;
    wire c12615;
    assign in12615_1 = {s10989[0]};
    assign in12615_2 = {s10990[0]};
    Full_Adder FA_12615(s12615, c12615, in12615_1, in12615_2, s10988[0]);
    wire[0:0] s12616, in12616_1, in12616_2;
    wire c12616;
    assign in12616_1 = {s8673[0]};
    assign in12616_2 = {c10983};
    Full_Adder FA_12616(s12616, c12616, in12616_1, in12616_2, s8672[0]);
    wire[0:0] s12617, in12617_1, in12617_2;
    wire c12617;
    assign in12617_1 = {c10985};
    assign in12617_2 = {c10986};
    Full_Adder FA_12617(s12617, c12617, in12617_1, in12617_2, c10984);
    wire[0:0] s12618, in12618_1, in12618_2;
    wire c12618;
    assign in12618_1 = {c10988};
    assign in12618_2 = {c10989};
    Full_Adder FA_12618(s12618, c12618, in12618_1, in12618_2, c10987);
    wire[0:0] s12619, in12619_1, in12619_2;
    wire c12619;
    assign in12619_1 = {s10991[0]};
    assign in12619_2 = {s10992[0]};
    Full_Adder FA_12619(s12619, c12619, in12619_1, in12619_2, c10990);
    wire[0:0] s12620, in12620_1, in12620_2;
    wire c12620;
    assign in12620_1 = {s10994[0]};
    assign in12620_2 = {s10995[0]};
    Full_Adder FA_12620(s12620, c12620, in12620_1, in12620_2, s10993[0]);
    wire[0:0] s12621, in12621_1, in12621_2;
    wire c12621;
    assign in12621_1 = {s10997[0]};
    assign in12621_2 = {s10998[0]};
    Full_Adder FA_12621(s12621, c12621, in12621_1, in12621_2, s10996[0]);
    wire[0:0] s12622, in12622_1, in12622_2;
    wire c12622;
    assign in12622_1 = {s8686[0]};
    assign in12622_2 = {c10991};
    Full_Adder FA_12622(s12622, c12622, in12622_1, in12622_2, s8685[0]);
    wire[0:0] s12623, in12623_1, in12623_2;
    wire c12623;
    assign in12623_1 = {c10993};
    assign in12623_2 = {c10994};
    Full_Adder FA_12623(s12623, c12623, in12623_1, in12623_2, c10992);
    wire[0:0] s12624, in12624_1, in12624_2;
    wire c12624;
    assign in12624_1 = {c10996};
    assign in12624_2 = {c10997};
    Full_Adder FA_12624(s12624, c12624, in12624_1, in12624_2, c10995);
    wire[0:0] s12625, in12625_1, in12625_2;
    wire c12625;
    assign in12625_1 = {s10999[0]};
    assign in12625_2 = {s11000[0]};
    Full_Adder FA_12625(s12625, c12625, in12625_1, in12625_2, c10998);
    wire[0:0] s12626, in12626_1, in12626_2;
    wire c12626;
    assign in12626_1 = {s11002[0]};
    assign in12626_2 = {s11003[0]};
    Full_Adder FA_12626(s12626, c12626, in12626_1, in12626_2, s11001[0]);
    wire[0:0] s12627, in12627_1, in12627_2;
    wire c12627;
    assign in12627_1 = {s11005[0]};
    assign in12627_2 = {s11006[0]};
    Full_Adder FA_12627(s12627, c12627, in12627_1, in12627_2, s11004[0]);
    wire[0:0] s12628, in12628_1, in12628_2;
    wire c12628;
    assign in12628_1 = {s8699[0]};
    assign in12628_2 = {c10999};
    Full_Adder FA_12628(s12628, c12628, in12628_1, in12628_2, s8698[0]);
    wire[0:0] s12629, in12629_1, in12629_2;
    wire c12629;
    assign in12629_1 = {c11001};
    assign in12629_2 = {c11002};
    Full_Adder FA_12629(s12629, c12629, in12629_1, in12629_2, c11000);
    wire[0:0] s12630, in12630_1, in12630_2;
    wire c12630;
    assign in12630_1 = {c11004};
    assign in12630_2 = {c11005};
    Full_Adder FA_12630(s12630, c12630, in12630_1, in12630_2, c11003);
    wire[0:0] s12631, in12631_1, in12631_2;
    wire c12631;
    assign in12631_1 = {s11007[0]};
    assign in12631_2 = {s11008[0]};
    Full_Adder FA_12631(s12631, c12631, in12631_1, in12631_2, c11006);
    wire[0:0] s12632, in12632_1, in12632_2;
    wire c12632;
    assign in12632_1 = {s11010[0]};
    assign in12632_2 = {s11011[0]};
    Full_Adder FA_12632(s12632, c12632, in12632_1, in12632_2, s11009[0]);
    wire[0:0] s12633, in12633_1, in12633_2;
    wire c12633;
    assign in12633_1 = {s11013[0]};
    assign in12633_2 = {s11014[0]};
    Full_Adder FA_12633(s12633, c12633, in12633_1, in12633_2, s11012[0]);
    wire[0:0] s12634, in12634_1, in12634_2;
    wire c12634;
    assign in12634_1 = {s8712[0]};
    assign in12634_2 = {c11007};
    Full_Adder FA_12634(s12634, c12634, in12634_1, in12634_2, s8711[0]);
    wire[0:0] s12635, in12635_1, in12635_2;
    wire c12635;
    assign in12635_1 = {c11009};
    assign in12635_2 = {c11010};
    Full_Adder FA_12635(s12635, c12635, in12635_1, in12635_2, c11008);
    wire[0:0] s12636, in12636_1, in12636_2;
    wire c12636;
    assign in12636_1 = {c11012};
    assign in12636_2 = {c11013};
    Full_Adder FA_12636(s12636, c12636, in12636_1, in12636_2, c11011);
    wire[0:0] s12637, in12637_1, in12637_2;
    wire c12637;
    assign in12637_1 = {s11015[0]};
    assign in12637_2 = {s11016[0]};
    Full_Adder FA_12637(s12637, c12637, in12637_1, in12637_2, c11014);
    wire[0:0] s12638, in12638_1, in12638_2;
    wire c12638;
    assign in12638_1 = {s11018[0]};
    assign in12638_2 = {s11019[0]};
    Full_Adder FA_12638(s12638, c12638, in12638_1, in12638_2, s11017[0]);
    wire[0:0] s12639, in12639_1, in12639_2;
    wire c12639;
    assign in12639_1 = {s11021[0]};
    assign in12639_2 = {s11022[0]};
    Full_Adder FA_12639(s12639, c12639, in12639_1, in12639_2, s11020[0]);
    wire[0:0] s12640, in12640_1, in12640_2;
    wire c12640;
    assign in12640_1 = {s8725[0]};
    assign in12640_2 = {c11015};
    Full_Adder FA_12640(s12640, c12640, in12640_1, in12640_2, s8724[0]);
    wire[0:0] s12641, in12641_1, in12641_2;
    wire c12641;
    assign in12641_1 = {c11017};
    assign in12641_2 = {c11018};
    Full_Adder FA_12641(s12641, c12641, in12641_1, in12641_2, c11016);
    wire[0:0] s12642, in12642_1, in12642_2;
    wire c12642;
    assign in12642_1 = {c11020};
    assign in12642_2 = {c11021};
    Full_Adder FA_12642(s12642, c12642, in12642_1, in12642_2, c11019);
    wire[0:0] s12643, in12643_1, in12643_2;
    wire c12643;
    assign in12643_1 = {s11023[0]};
    assign in12643_2 = {s11024[0]};
    Full_Adder FA_12643(s12643, c12643, in12643_1, in12643_2, c11022);
    wire[0:0] s12644, in12644_1, in12644_2;
    wire c12644;
    assign in12644_1 = {s11026[0]};
    assign in12644_2 = {s11027[0]};
    Full_Adder FA_12644(s12644, c12644, in12644_1, in12644_2, s11025[0]);
    wire[0:0] s12645, in12645_1, in12645_2;
    wire c12645;
    assign in12645_1 = {s11029[0]};
    assign in12645_2 = {s11030[0]};
    Full_Adder FA_12645(s12645, c12645, in12645_1, in12645_2, s11028[0]);
    wire[0:0] s12646, in12646_1, in12646_2;
    wire c12646;
    assign in12646_1 = {s8738[0]};
    assign in12646_2 = {c11023};
    Full_Adder FA_12646(s12646, c12646, in12646_1, in12646_2, s8737[0]);
    wire[0:0] s12647, in12647_1, in12647_2;
    wire c12647;
    assign in12647_1 = {c11025};
    assign in12647_2 = {c11026};
    Full_Adder FA_12647(s12647, c12647, in12647_1, in12647_2, c11024);
    wire[0:0] s12648, in12648_1, in12648_2;
    wire c12648;
    assign in12648_1 = {c11028};
    assign in12648_2 = {c11029};
    Full_Adder FA_12648(s12648, c12648, in12648_1, in12648_2, c11027);
    wire[0:0] s12649, in12649_1, in12649_2;
    wire c12649;
    assign in12649_1 = {s11031[0]};
    assign in12649_2 = {s11032[0]};
    Full_Adder FA_12649(s12649, c12649, in12649_1, in12649_2, c11030);
    wire[0:0] s12650, in12650_1, in12650_2;
    wire c12650;
    assign in12650_1 = {s11034[0]};
    assign in12650_2 = {s11035[0]};
    Full_Adder FA_12650(s12650, c12650, in12650_1, in12650_2, s11033[0]);
    wire[0:0] s12651, in12651_1, in12651_2;
    wire c12651;
    assign in12651_1 = {s11037[0]};
    assign in12651_2 = {s11038[0]};
    Full_Adder FA_12651(s12651, c12651, in12651_1, in12651_2, s11036[0]);
    wire[0:0] s12652, in12652_1, in12652_2;
    wire c12652;
    assign in12652_1 = {s8751[0]};
    assign in12652_2 = {c11031};
    Full_Adder FA_12652(s12652, c12652, in12652_1, in12652_2, s8750[0]);
    wire[0:0] s12653, in12653_1, in12653_2;
    wire c12653;
    assign in12653_1 = {c11033};
    assign in12653_2 = {c11034};
    Full_Adder FA_12653(s12653, c12653, in12653_1, in12653_2, c11032);
    wire[0:0] s12654, in12654_1, in12654_2;
    wire c12654;
    assign in12654_1 = {c11036};
    assign in12654_2 = {c11037};
    Full_Adder FA_12654(s12654, c12654, in12654_1, in12654_2, c11035);
    wire[0:0] s12655, in12655_1, in12655_2;
    wire c12655;
    assign in12655_1 = {s11039[0]};
    assign in12655_2 = {s11040[0]};
    Full_Adder FA_12655(s12655, c12655, in12655_1, in12655_2, c11038);
    wire[0:0] s12656, in12656_1, in12656_2;
    wire c12656;
    assign in12656_1 = {s11042[0]};
    assign in12656_2 = {s11043[0]};
    Full_Adder FA_12656(s12656, c12656, in12656_1, in12656_2, s11041[0]);
    wire[0:0] s12657, in12657_1, in12657_2;
    wire c12657;
    assign in12657_1 = {s11045[0]};
    assign in12657_2 = {s11046[0]};
    Full_Adder FA_12657(s12657, c12657, in12657_1, in12657_2, s11044[0]);
    wire[0:0] s12658, in12658_1, in12658_2;
    wire c12658;
    assign in12658_1 = {s8764[0]};
    assign in12658_2 = {c11039};
    Full_Adder FA_12658(s12658, c12658, in12658_1, in12658_2, s8763[0]);
    wire[0:0] s12659, in12659_1, in12659_2;
    wire c12659;
    assign in12659_1 = {c11041};
    assign in12659_2 = {c11042};
    Full_Adder FA_12659(s12659, c12659, in12659_1, in12659_2, c11040);
    wire[0:0] s12660, in12660_1, in12660_2;
    wire c12660;
    assign in12660_1 = {c11044};
    assign in12660_2 = {c11045};
    Full_Adder FA_12660(s12660, c12660, in12660_1, in12660_2, c11043);
    wire[0:0] s12661, in12661_1, in12661_2;
    wire c12661;
    assign in12661_1 = {s11047[0]};
    assign in12661_2 = {s11048[0]};
    Full_Adder FA_12661(s12661, c12661, in12661_1, in12661_2, c11046);
    wire[0:0] s12662, in12662_1, in12662_2;
    wire c12662;
    assign in12662_1 = {s11050[0]};
    assign in12662_2 = {s11051[0]};
    Full_Adder FA_12662(s12662, c12662, in12662_1, in12662_2, s11049[0]);
    wire[0:0] s12663, in12663_1, in12663_2;
    wire c12663;
    assign in12663_1 = {s11053[0]};
    assign in12663_2 = {s11054[0]};
    Full_Adder FA_12663(s12663, c12663, in12663_1, in12663_2, s11052[0]);
    wire[0:0] s12664, in12664_1, in12664_2;
    wire c12664;
    assign in12664_1 = {s8777[0]};
    assign in12664_2 = {c11047};
    Full_Adder FA_12664(s12664, c12664, in12664_1, in12664_2, s8776[0]);
    wire[0:0] s12665, in12665_1, in12665_2;
    wire c12665;
    assign in12665_1 = {c11049};
    assign in12665_2 = {c11050};
    Full_Adder FA_12665(s12665, c12665, in12665_1, in12665_2, c11048);
    wire[0:0] s12666, in12666_1, in12666_2;
    wire c12666;
    assign in12666_1 = {c11052};
    assign in12666_2 = {c11053};
    Full_Adder FA_12666(s12666, c12666, in12666_1, in12666_2, c11051);
    wire[0:0] s12667, in12667_1, in12667_2;
    wire c12667;
    assign in12667_1 = {s11055[0]};
    assign in12667_2 = {s11056[0]};
    Full_Adder FA_12667(s12667, c12667, in12667_1, in12667_2, c11054);
    wire[0:0] s12668, in12668_1, in12668_2;
    wire c12668;
    assign in12668_1 = {s11058[0]};
    assign in12668_2 = {s11059[0]};
    Full_Adder FA_12668(s12668, c12668, in12668_1, in12668_2, s11057[0]);
    wire[0:0] s12669, in12669_1, in12669_2;
    wire c12669;
    assign in12669_1 = {s11061[0]};
    assign in12669_2 = {s11062[0]};
    Full_Adder FA_12669(s12669, c12669, in12669_1, in12669_2, s11060[0]);
    wire[0:0] s12670, in12670_1, in12670_2;
    wire c12670;
    assign in12670_1 = {s8790[0]};
    assign in12670_2 = {c11055};
    Full_Adder FA_12670(s12670, c12670, in12670_1, in12670_2, s8789[0]);
    wire[0:0] s12671, in12671_1, in12671_2;
    wire c12671;
    assign in12671_1 = {c11057};
    assign in12671_2 = {c11058};
    Full_Adder FA_12671(s12671, c12671, in12671_1, in12671_2, c11056);
    wire[0:0] s12672, in12672_1, in12672_2;
    wire c12672;
    assign in12672_1 = {c11060};
    assign in12672_2 = {c11061};
    Full_Adder FA_12672(s12672, c12672, in12672_1, in12672_2, c11059);
    wire[0:0] s12673, in12673_1, in12673_2;
    wire c12673;
    assign in12673_1 = {s11063[0]};
    assign in12673_2 = {s11064[0]};
    Full_Adder FA_12673(s12673, c12673, in12673_1, in12673_2, c11062);
    wire[0:0] s12674, in12674_1, in12674_2;
    wire c12674;
    assign in12674_1 = {s11066[0]};
    assign in12674_2 = {s11067[0]};
    Full_Adder FA_12674(s12674, c12674, in12674_1, in12674_2, s11065[0]);
    wire[0:0] s12675, in12675_1, in12675_2;
    wire c12675;
    assign in12675_1 = {s11069[0]};
    assign in12675_2 = {s11070[0]};
    Full_Adder FA_12675(s12675, c12675, in12675_1, in12675_2, s11068[0]);
    wire[0:0] s12676, in12676_1, in12676_2;
    wire c12676;
    assign in12676_1 = {s8803[0]};
    assign in12676_2 = {c11063};
    Full_Adder FA_12676(s12676, c12676, in12676_1, in12676_2, s8802[0]);
    wire[0:0] s12677, in12677_1, in12677_2;
    wire c12677;
    assign in12677_1 = {c11065};
    assign in12677_2 = {c11066};
    Full_Adder FA_12677(s12677, c12677, in12677_1, in12677_2, c11064);
    wire[0:0] s12678, in12678_1, in12678_2;
    wire c12678;
    assign in12678_1 = {c11068};
    assign in12678_2 = {c11069};
    Full_Adder FA_12678(s12678, c12678, in12678_1, in12678_2, c11067);
    wire[0:0] s12679, in12679_1, in12679_2;
    wire c12679;
    assign in12679_1 = {s11071[0]};
    assign in12679_2 = {s11072[0]};
    Full_Adder FA_12679(s12679, c12679, in12679_1, in12679_2, c11070);
    wire[0:0] s12680, in12680_1, in12680_2;
    wire c12680;
    assign in12680_1 = {s11074[0]};
    assign in12680_2 = {s11075[0]};
    Full_Adder FA_12680(s12680, c12680, in12680_1, in12680_2, s11073[0]);
    wire[0:0] s12681, in12681_1, in12681_2;
    wire c12681;
    assign in12681_1 = {s11077[0]};
    assign in12681_2 = {s11078[0]};
    Full_Adder FA_12681(s12681, c12681, in12681_1, in12681_2, s11076[0]);
    wire[0:0] s12682, in12682_1, in12682_2;
    wire c12682;
    assign in12682_1 = {s8816[0]};
    assign in12682_2 = {c11071};
    Full_Adder FA_12682(s12682, c12682, in12682_1, in12682_2, s8815[0]);
    wire[0:0] s12683, in12683_1, in12683_2;
    wire c12683;
    assign in12683_1 = {c11073};
    assign in12683_2 = {c11074};
    Full_Adder FA_12683(s12683, c12683, in12683_1, in12683_2, c11072);
    wire[0:0] s12684, in12684_1, in12684_2;
    wire c12684;
    assign in12684_1 = {c11076};
    assign in12684_2 = {c11077};
    Full_Adder FA_12684(s12684, c12684, in12684_1, in12684_2, c11075);
    wire[0:0] s12685, in12685_1, in12685_2;
    wire c12685;
    assign in12685_1 = {s11079[0]};
    assign in12685_2 = {s11080[0]};
    Full_Adder FA_12685(s12685, c12685, in12685_1, in12685_2, c11078);
    wire[0:0] s12686, in12686_1, in12686_2;
    wire c12686;
    assign in12686_1 = {s11082[0]};
    assign in12686_2 = {s11083[0]};
    Full_Adder FA_12686(s12686, c12686, in12686_1, in12686_2, s11081[0]);
    wire[0:0] s12687, in12687_1, in12687_2;
    wire c12687;
    assign in12687_1 = {s11085[0]};
    assign in12687_2 = {s11086[0]};
    Full_Adder FA_12687(s12687, c12687, in12687_1, in12687_2, s11084[0]);
    wire[0:0] s12688, in12688_1, in12688_2;
    wire c12688;
    assign in12688_1 = {s8829[0]};
    assign in12688_2 = {c11079};
    Full_Adder FA_12688(s12688, c12688, in12688_1, in12688_2, s8828[0]);
    wire[0:0] s12689, in12689_1, in12689_2;
    wire c12689;
    assign in12689_1 = {c11081};
    assign in12689_2 = {c11082};
    Full_Adder FA_12689(s12689, c12689, in12689_1, in12689_2, c11080);
    wire[0:0] s12690, in12690_1, in12690_2;
    wire c12690;
    assign in12690_1 = {c11084};
    assign in12690_2 = {c11085};
    Full_Adder FA_12690(s12690, c12690, in12690_1, in12690_2, c11083);
    wire[0:0] s12691, in12691_1, in12691_2;
    wire c12691;
    assign in12691_1 = {s11087[0]};
    assign in12691_2 = {s11088[0]};
    Full_Adder FA_12691(s12691, c12691, in12691_1, in12691_2, c11086);
    wire[0:0] s12692, in12692_1, in12692_2;
    wire c12692;
    assign in12692_1 = {s11090[0]};
    assign in12692_2 = {s11091[0]};
    Full_Adder FA_12692(s12692, c12692, in12692_1, in12692_2, s11089[0]);
    wire[0:0] s12693, in12693_1, in12693_2;
    wire c12693;
    assign in12693_1 = {s11093[0]};
    assign in12693_2 = {s11094[0]};
    Full_Adder FA_12693(s12693, c12693, in12693_1, in12693_2, s11092[0]);
    wire[0:0] s12694, in12694_1, in12694_2;
    wire c12694;
    assign in12694_1 = {s8842[0]};
    assign in12694_2 = {c11087};
    Full_Adder FA_12694(s12694, c12694, in12694_1, in12694_2, s8841[0]);
    wire[0:0] s12695, in12695_1, in12695_2;
    wire c12695;
    assign in12695_1 = {c11089};
    assign in12695_2 = {c11090};
    Full_Adder FA_12695(s12695, c12695, in12695_1, in12695_2, c11088);
    wire[0:0] s12696, in12696_1, in12696_2;
    wire c12696;
    assign in12696_1 = {c11092};
    assign in12696_2 = {c11093};
    Full_Adder FA_12696(s12696, c12696, in12696_1, in12696_2, c11091);
    wire[0:0] s12697, in12697_1, in12697_2;
    wire c12697;
    assign in12697_1 = {s11095[0]};
    assign in12697_2 = {s11096[0]};
    Full_Adder FA_12697(s12697, c12697, in12697_1, in12697_2, c11094);
    wire[0:0] s12698, in12698_1, in12698_2;
    wire c12698;
    assign in12698_1 = {s11098[0]};
    assign in12698_2 = {s11099[0]};
    Full_Adder FA_12698(s12698, c12698, in12698_1, in12698_2, s11097[0]);
    wire[0:0] s12699, in12699_1, in12699_2;
    wire c12699;
    assign in12699_1 = {s11101[0]};
    assign in12699_2 = {s11102[0]};
    Full_Adder FA_12699(s12699, c12699, in12699_1, in12699_2, s11100[0]);
    wire[0:0] s12700, in12700_1, in12700_2;
    wire c12700;
    assign in12700_1 = {s8855[0]};
    assign in12700_2 = {c11095};
    Full_Adder FA_12700(s12700, c12700, in12700_1, in12700_2, s8854[0]);
    wire[0:0] s12701, in12701_1, in12701_2;
    wire c12701;
    assign in12701_1 = {c11097};
    assign in12701_2 = {c11098};
    Full_Adder FA_12701(s12701, c12701, in12701_1, in12701_2, c11096);
    wire[0:0] s12702, in12702_1, in12702_2;
    wire c12702;
    assign in12702_1 = {c11100};
    assign in12702_2 = {c11101};
    Full_Adder FA_12702(s12702, c12702, in12702_1, in12702_2, c11099);
    wire[0:0] s12703, in12703_1, in12703_2;
    wire c12703;
    assign in12703_1 = {s11103[0]};
    assign in12703_2 = {s11104[0]};
    Full_Adder FA_12703(s12703, c12703, in12703_1, in12703_2, c11102);
    wire[0:0] s12704, in12704_1, in12704_2;
    wire c12704;
    assign in12704_1 = {s11106[0]};
    assign in12704_2 = {s11107[0]};
    Full_Adder FA_12704(s12704, c12704, in12704_1, in12704_2, s11105[0]);
    wire[0:0] s12705, in12705_1, in12705_2;
    wire c12705;
    assign in12705_1 = {s11109[0]};
    assign in12705_2 = {s11110[0]};
    Full_Adder FA_12705(s12705, c12705, in12705_1, in12705_2, s11108[0]);
    wire[0:0] s12706, in12706_1, in12706_2;
    wire c12706;
    assign in12706_1 = {s8868[0]};
    assign in12706_2 = {c11103};
    Full_Adder FA_12706(s12706, c12706, in12706_1, in12706_2, s8867[0]);
    wire[0:0] s12707, in12707_1, in12707_2;
    wire c12707;
    assign in12707_1 = {c11105};
    assign in12707_2 = {c11106};
    Full_Adder FA_12707(s12707, c12707, in12707_1, in12707_2, c11104);
    wire[0:0] s12708, in12708_1, in12708_2;
    wire c12708;
    assign in12708_1 = {c11108};
    assign in12708_2 = {c11109};
    Full_Adder FA_12708(s12708, c12708, in12708_1, in12708_2, c11107);
    wire[0:0] s12709, in12709_1, in12709_2;
    wire c12709;
    assign in12709_1 = {s11111[0]};
    assign in12709_2 = {s11112[0]};
    Full_Adder FA_12709(s12709, c12709, in12709_1, in12709_2, c11110);
    wire[0:0] s12710, in12710_1, in12710_2;
    wire c12710;
    assign in12710_1 = {s11114[0]};
    assign in12710_2 = {s11115[0]};
    Full_Adder FA_12710(s12710, c12710, in12710_1, in12710_2, s11113[0]);
    wire[0:0] s12711, in12711_1, in12711_2;
    wire c12711;
    assign in12711_1 = {s11117[0]};
    assign in12711_2 = {s11118[0]};
    Full_Adder FA_12711(s12711, c12711, in12711_1, in12711_2, s11116[0]);
    wire[0:0] s12712, in12712_1, in12712_2;
    wire c12712;
    assign in12712_1 = {s8881[0]};
    assign in12712_2 = {c11111};
    Full_Adder FA_12712(s12712, c12712, in12712_1, in12712_2, s8880[0]);
    wire[0:0] s12713, in12713_1, in12713_2;
    wire c12713;
    assign in12713_1 = {c11113};
    assign in12713_2 = {c11114};
    Full_Adder FA_12713(s12713, c12713, in12713_1, in12713_2, c11112);
    wire[0:0] s12714, in12714_1, in12714_2;
    wire c12714;
    assign in12714_1 = {c11116};
    assign in12714_2 = {c11117};
    Full_Adder FA_12714(s12714, c12714, in12714_1, in12714_2, c11115);
    wire[0:0] s12715, in12715_1, in12715_2;
    wire c12715;
    assign in12715_1 = {s11119[0]};
    assign in12715_2 = {s11120[0]};
    Full_Adder FA_12715(s12715, c12715, in12715_1, in12715_2, c11118);
    wire[0:0] s12716, in12716_1, in12716_2;
    wire c12716;
    assign in12716_1 = {s11122[0]};
    assign in12716_2 = {s11123[0]};
    Full_Adder FA_12716(s12716, c12716, in12716_1, in12716_2, s11121[0]);
    wire[0:0] s12717, in12717_1, in12717_2;
    wire c12717;
    assign in12717_1 = {s11125[0]};
    assign in12717_2 = {s11126[0]};
    Full_Adder FA_12717(s12717, c12717, in12717_1, in12717_2, s11124[0]);
    wire[0:0] s12718, in12718_1, in12718_2;
    wire c12718;
    assign in12718_1 = {s8894[0]};
    assign in12718_2 = {c11119};
    Full_Adder FA_12718(s12718, c12718, in12718_1, in12718_2, s8893[0]);
    wire[0:0] s12719, in12719_1, in12719_2;
    wire c12719;
    assign in12719_1 = {c11121};
    assign in12719_2 = {c11122};
    Full_Adder FA_12719(s12719, c12719, in12719_1, in12719_2, c11120);
    wire[0:0] s12720, in12720_1, in12720_2;
    wire c12720;
    assign in12720_1 = {c11124};
    assign in12720_2 = {c11125};
    Full_Adder FA_12720(s12720, c12720, in12720_1, in12720_2, c11123);
    wire[0:0] s12721, in12721_1, in12721_2;
    wire c12721;
    assign in12721_1 = {s11127[0]};
    assign in12721_2 = {s11128[0]};
    Full_Adder FA_12721(s12721, c12721, in12721_1, in12721_2, c11126);
    wire[0:0] s12722, in12722_1, in12722_2;
    wire c12722;
    assign in12722_1 = {s11130[0]};
    assign in12722_2 = {s11131[0]};
    Full_Adder FA_12722(s12722, c12722, in12722_1, in12722_2, s11129[0]);
    wire[0:0] s12723, in12723_1, in12723_2;
    wire c12723;
    assign in12723_1 = {s11133[0]};
    assign in12723_2 = {s11134[0]};
    Full_Adder FA_12723(s12723, c12723, in12723_1, in12723_2, s11132[0]);
    wire[0:0] s12724, in12724_1, in12724_2;
    wire c12724;
    assign in12724_1 = {s8907[0]};
    assign in12724_2 = {c11127};
    Full_Adder FA_12724(s12724, c12724, in12724_1, in12724_2, s8906[0]);
    wire[0:0] s12725, in12725_1, in12725_2;
    wire c12725;
    assign in12725_1 = {c11129};
    assign in12725_2 = {c11130};
    Full_Adder FA_12725(s12725, c12725, in12725_1, in12725_2, c11128);
    wire[0:0] s12726, in12726_1, in12726_2;
    wire c12726;
    assign in12726_1 = {c11132};
    assign in12726_2 = {c11133};
    Full_Adder FA_12726(s12726, c12726, in12726_1, in12726_2, c11131);
    wire[0:0] s12727, in12727_1, in12727_2;
    wire c12727;
    assign in12727_1 = {s11135[0]};
    assign in12727_2 = {s11136[0]};
    Full_Adder FA_12727(s12727, c12727, in12727_1, in12727_2, c11134);
    wire[0:0] s12728, in12728_1, in12728_2;
    wire c12728;
    assign in12728_1 = {s11138[0]};
    assign in12728_2 = {s11139[0]};
    Full_Adder FA_12728(s12728, c12728, in12728_1, in12728_2, s11137[0]);
    wire[0:0] s12729, in12729_1, in12729_2;
    wire c12729;
    assign in12729_1 = {s11141[0]};
    assign in12729_2 = {s11142[0]};
    Full_Adder FA_12729(s12729, c12729, in12729_1, in12729_2, s11140[0]);
    wire[0:0] s12730, in12730_1, in12730_2;
    wire c12730;
    assign in12730_1 = {s8920[0]};
    assign in12730_2 = {c11135};
    Full_Adder FA_12730(s12730, c12730, in12730_1, in12730_2, s8919[0]);
    wire[0:0] s12731, in12731_1, in12731_2;
    wire c12731;
    assign in12731_1 = {c11137};
    assign in12731_2 = {c11138};
    Full_Adder FA_12731(s12731, c12731, in12731_1, in12731_2, c11136);
    wire[0:0] s12732, in12732_1, in12732_2;
    wire c12732;
    assign in12732_1 = {c11140};
    assign in12732_2 = {c11141};
    Full_Adder FA_12732(s12732, c12732, in12732_1, in12732_2, c11139);
    wire[0:0] s12733, in12733_1, in12733_2;
    wire c12733;
    assign in12733_1 = {s11143[0]};
    assign in12733_2 = {s11144[0]};
    Full_Adder FA_12733(s12733, c12733, in12733_1, in12733_2, c11142);
    wire[0:0] s12734, in12734_1, in12734_2;
    wire c12734;
    assign in12734_1 = {s11146[0]};
    assign in12734_2 = {s11147[0]};
    Full_Adder FA_12734(s12734, c12734, in12734_1, in12734_2, s11145[0]);
    wire[0:0] s12735, in12735_1, in12735_2;
    wire c12735;
    assign in12735_1 = {s11149[0]};
    assign in12735_2 = {s11150[0]};
    Full_Adder FA_12735(s12735, c12735, in12735_1, in12735_2, s11148[0]);
    wire[0:0] s12736, in12736_1, in12736_2;
    wire c12736;
    assign in12736_1 = {s8933[0]};
    assign in12736_2 = {c11143};
    Full_Adder FA_12736(s12736, c12736, in12736_1, in12736_2, s8932[0]);
    wire[0:0] s12737, in12737_1, in12737_2;
    wire c12737;
    assign in12737_1 = {c11145};
    assign in12737_2 = {c11146};
    Full_Adder FA_12737(s12737, c12737, in12737_1, in12737_2, c11144);
    wire[0:0] s12738, in12738_1, in12738_2;
    wire c12738;
    assign in12738_1 = {c11148};
    assign in12738_2 = {c11149};
    Full_Adder FA_12738(s12738, c12738, in12738_1, in12738_2, c11147);
    wire[0:0] s12739, in12739_1, in12739_2;
    wire c12739;
    assign in12739_1 = {s11151[0]};
    assign in12739_2 = {s11152[0]};
    Full_Adder FA_12739(s12739, c12739, in12739_1, in12739_2, c11150);
    wire[0:0] s12740, in12740_1, in12740_2;
    wire c12740;
    assign in12740_1 = {s11154[0]};
    assign in12740_2 = {s11155[0]};
    Full_Adder FA_12740(s12740, c12740, in12740_1, in12740_2, s11153[0]);
    wire[0:0] s12741, in12741_1, in12741_2;
    wire c12741;
    assign in12741_1 = {s11157[0]};
    assign in12741_2 = {s11158[0]};
    Full_Adder FA_12741(s12741, c12741, in12741_1, in12741_2, s11156[0]);
    wire[0:0] s12742, in12742_1, in12742_2;
    wire c12742;
    assign in12742_1 = {s8946[0]};
    assign in12742_2 = {c11151};
    Full_Adder FA_12742(s12742, c12742, in12742_1, in12742_2, s8945[0]);
    wire[0:0] s12743, in12743_1, in12743_2;
    wire c12743;
    assign in12743_1 = {c11153};
    assign in12743_2 = {c11154};
    Full_Adder FA_12743(s12743, c12743, in12743_1, in12743_2, c11152);
    wire[0:0] s12744, in12744_1, in12744_2;
    wire c12744;
    assign in12744_1 = {c11156};
    assign in12744_2 = {c11157};
    Full_Adder FA_12744(s12744, c12744, in12744_1, in12744_2, c11155);
    wire[0:0] s12745, in12745_1, in12745_2;
    wire c12745;
    assign in12745_1 = {s11159[0]};
    assign in12745_2 = {s11160[0]};
    Full_Adder FA_12745(s12745, c12745, in12745_1, in12745_2, c11158);
    wire[0:0] s12746, in12746_1, in12746_2;
    wire c12746;
    assign in12746_1 = {s11162[0]};
    assign in12746_2 = {s11163[0]};
    Full_Adder FA_12746(s12746, c12746, in12746_1, in12746_2, s11161[0]);
    wire[0:0] s12747, in12747_1, in12747_2;
    wire c12747;
    assign in12747_1 = {s11165[0]};
    assign in12747_2 = {s11166[0]};
    Full_Adder FA_12747(s12747, c12747, in12747_1, in12747_2, s11164[0]);
    wire[0:0] s12748, in12748_1, in12748_2;
    wire c12748;
    assign in12748_1 = {s8959[0]};
    assign in12748_2 = {c11159};
    Full_Adder FA_12748(s12748, c12748, in12748_1, in12748_2, s8958[0]);
    wire[0:0] s12749, in12749_1, in12749_2;
    wire c12749;
    assign in12749_1 = {c11161};
    assign in12749_2 = {c11162};
    Full_Adder FA_12749(s12749, c12749, in12749_1, in12749_2, c11160);
    wire[0:0] s12750, in12750_1, in12750_2;
    wire c12750;
    assign in12750_1 = {c11164};
    assign in12750_2 = {c11165};
    Full_Adder FA_12750(s12750, c12750, in12750_1, in12750_2, c11163);
    wire[0:0] s12751, in12751_1, in12751_2;
    wire c12751;
    assign in12751_1 = {s11167[0]};
    assign in12751_2 = {s11168[0]};
    Full_Adder FA_12751(s12751, c12751, in12751_1, in12751_2, c11166);
    wire[0:0] s12752, in12752_1, in12752_2;
    wire c12752;
    assign in12752_1 = {s11170[0]};
    assign in12752_2 = {s11171[0]};
    Full_Adder FA_12752(s12752, c12752, in12752_1, in12752_2, s11169[0]);
    wire[0:0] s12753, in12753_1, in12753_2;
    wire c12753;
    assign in12753_1 = {s11173[0]};
    assign in12753_2 = {s11174[0]};
    Full_Adder FA_12753(s12753, c12753, in12753_1, in12753_2, s11172[0]);
    wire[0:0] s12754, in12754_1, in12754_2;
    wire c12754;
    assign in12754_1 = {s8972[0]};
    assign in12754_2 = {c11167};
    Full_Adder FA_12754(s12754, c12754, in12754_1, in12754_2, s8971[0]);
    wire[0:0] s12755, in12755_1, in12755_2;
    wire c12755;
    assign in12755_1 = {c11169};
    assign in12755_2 = {c11170};
    Full_Adder FA_12755(s12755, c12755, in12755_1, in12755_2, c11168);
    wire[0:0] s12756, in12756_1, in12756_2;
    wire c12756;
    assign in12756_1 = {c11172};
    assign in12756_2 = {c11173};
    Full_Adder FA_12756(s12756, c12756, in12756_1, in12756_2, c11171);
    wire[0:0] s12757, in12757_1, in12757_2;
    wire c12757;
    assign in12757_1 = {s11175[0]};
    assign in12757_2 = {s11176[0]};
    Full_Adder FA_12757(s12757, c12757, in12757_1, in12757_2, c11174);
    wire[0:0] s12758, in12758_1, in12758_2;
    wire c12758;
    assign in12758_1 = {s11178[0]};
    assign in12758_2 = {s11179[0]};
    Full_Adder FA_12758(s12758, c12758, in12758_1, in12758_2, s11177[0]);
    wire[0:0] s12759, in12759_1, in12759_2;
    wire c12759;
    assign in12759_1 = {s11181[0]};
    assign in12759_2 = {s11182[0]};
    Full_Adder FA_12759(s12759, c12759, in12759_1, in12759_2, s11180[0]);
    wire[0:0] s12760, in12760_1, in12760_2;
    wire c12760;
    assign in12760_1 = {s8985[0]};
    assign in12760_2 = {c11175};
    Full_Adder FA_12760(s12760, c12760, in12760_1, in12760_2, s8984[0]);
    wire[0:0] s12761, in12761_1, in12761_2;
    wire c12761;
    assign in12761_1 = {c11177};
    assign in12761_2 = {c11178};
    Full_Adder FA_12761(s12761, c12761, in12761_1, in12761_2, c11176);
    wire[0:0] s12762, in12762_1, in12762_2;
    wire c12762;
    assign in12762_1 = {c11180};
    assign in12762_2 = {c11181};
    Full_Adder FA_12762(s12762, c12762, in12762_1, in12762_2, c11179);
    wire[0:0] s12763, in12763_1, in12763_2;
    wire c12763;
    assign in12763_1 = {s11183[0]};
    assign in12763_2 = {s11184[0]};
    Full_Adder FA_12763(s12763, c12763, in12763_1, in12763_2, c11182);
    wire[0:0] s12764, in12764_1, in12764_2;
    wire c12764;
    assign in12764_1 = {s11186[0]};
    assign in12764_2 = {s11187[0]};
    Full_Adder FA_12764(s12764, c12764, in12764_1, in12764_2, s11185[0]);
    wire[0:0] s12765, in12765_1, in12765_2;
    wire c12765;
    assign in12765_1 = {s11189[0]};
    assign in12765_2 = {s11190[0]};
    Full_Adder FA_12765(s12765, c12765, in12765_1, in12765_2, s11188[0]);
    wire[0:0] s12766, in12766_1, in12766_2;
    wire c12766;
    assign in12766_1 = {s8998[0]};
    assign in12766_2 = {c11183};
    Full_Adder FA_12766(s12766, c12766, in12766_1, in12766_2, s8997[0]);
    wire[0:0] s12767, in12767_1, in12767_2;
    wire c12767;
    assign in12767_1 = {c11185};
    assign in12767_2 = {c11186};
    Full_Adder FA_12767(s12767, c12767, in12767_1, in12767_2, c11184);
    wire[0:0] s12768, in12768_1, in12768_2;
    wire c12768;
    assign in12768_1 = {c11188};
    assign in12768_2 = {c11189};
    Full_Adder FA_12768(s12768, c12768, in12768_1, in12768_2, c11187);
    wire[0:0] s12769, in12769_1, in12769_2;
    wire c12769;
    assign in12769_1 = {s11191[0]};
    assign in12769_2 = {s11192[0]};
    Full_Adder FA_12769(s12769, c12769, in12769_1, in12769_2, c11190);
    wire[0:0] s12770, in12770_1, in12770_2;
    wire c12770;
    assign in12770_1 = {s11194[0]};
    assign in12770_2 = {s11195[0]};
    Full_Adder FA_12770(s12770, c12770, in12770_1, in12770_2, s11193[0]);
    wire[0:0] s12771, in12771_1, in12771_2;
    wire c12771;
    assign in12771_1 = {s11197[0]};
    assign in12771_2 = {s11198[0]};
    Full_Adder FA_12771(s12771, c12771, in12771_1, in12771_2, s11196[0]);
    wire[0:0] s12772, in12772_1, in12772_2;
    wire c12772;
    assign in12772_1 = {s9011[0]};
    assign in12772_2 = {c11191};
    Full_Adder FA_12772(s12772, c12772, in12772_1, in12772_2, s9010[0]);
    wire[0:0] s12773, in12773_1, in12773_2;
    wire c12773;
    assign in12773_1 = {c11193};
    assign in12773_2 = {c11194};
    Full_Adder FA_12773(s12773, c12773, in12773_1, in12773_2, c11192);
    wire[0:0] s12774, in12774_1, in12774_2;
    wire c12774;
    assign in12774_1 = {c11196};
    assign in12774_2 = {c11197};
    Full_Adder FA_12774(s12774, c12774, in12774_1, in12774_2, c11195);
    wire[0:0] s12775, in12775_1, in12775_2;
    wire c12775;
    assign in12775_1 = {s11199[0]};
    assign in12775_2 = {s11200[0]};
    Full_Adder FA_12775(s12775, c12775, in12775_1, in12775_2, c11198);
    wire[0:0] s12776, in12776_1, in12776_2;
    wire c12776;
    assign in12776_1 = {s11202[0]};
    assign in12776_2 = {s11203[0]};
    Full_Adder FA_12776(s12776, c12776, in12776_1, in12776_2, s11201[0]);
    wire[0:0] s12777, in12777_1, in12777_2;
    wire c12777;
    assign in12777_1 = {s11205[0]};
    assign in12777_2 = {s11206[0]};
    Full_Adder FA_12777(s12777, c12777, in12777_1, in12777_2, s11204[0]);
    wire[0:0] s12778, in12778_1, in12778_2;
    wire c12778;
    assign in12778_1 = {s9024[0]};
    assign in12778_2 = {c11199};
    Full_Adder FA_12778(s12778, c12778, in12778_1, in12778_2, s9023[0]);
    wire[0:0] s12779, in12779_1, in12779_2;
    wire c12779;
    assign in12779_1 = {c11201};
    assign in12779_2 = {c11202};
    Full_Adder FA_12779(s12779, c12779, in12779_1, in12779_2, c11200);
    wire[0:0] s12780, in12780_1, in12780_2;
    wire c12780;
    assign in12780_1 = {c11204};
    assign in12780_2 = {c11205};
    Full_Adder FA_12780(s12780, c12780, in12780_1, in12780_2, c11203);
    wire[0:0] s12781, in12781_1, in12781_2;
    wire c12781;
    assign in12781_1 = {s11207[0]};
    assign in12781_2 = {s11208[0]};
    Full_Adder FA_12781(s12781, c12781, in12781_1, in12781_2, c11206);
    wire[0:0] s12782, in12782_1, in12782_2;
    wire c12782;
    assign in12782_1 = {s11210[0]};
    assign in12782_2 = {s11211[0]};
    Full_Adder FA_12782(s12782, c12782, in12782_1, in12782_2, s11209[0]);
    wire[0:0] s12783, in12783_1, in12783_2;
    wire c12783;
    assign in12783_1 = {s11213[0]};
    assign in12783_2 = {s11214[0]};
    Full_Adder FA_12783(s12783, c12783, in12783_1, in12783_2, s11212[0]);
    wire[0:0] s12784, in12784_1, in12784_2;
    wire c12784;
    assign in12784_1 = {s9037[0]};
    assign in12784_2 = {c11207};
    Full_Adder FA_12784(s12784, c12784, in12784_1, in12784_2, s9036[0]);
    wire[0:0] s12785, in12785_1, in12785_2;
    wire c12785;
    assign in12785_1 = {c11209};
    assign in12785_2 = {c11210};
    Full_Adder FA_12785(s12785, c12785, in12785_1, in12785_2, c11208);
    wire[0:0] s12786, in12786_1, in12786_2;
    wire c12786;
    assign in12786_1 = {c11212};
    assign in12786_2 = {c11213};
    Full_Adder FA_12786(s12786, c12786, in12786_1, in12786_2, c11211);
    wire[0:0] s12787, in12787_1, in12787_2;
    wire c12787;
    assign in12787_1 = {s11215[0]};
    assign in12787_2 = {s11216[0]};
    Full_Adder FA_12787(s12787, c12787, in12787_1, in12787_2, c11214);
    wire[0:0] s12788, in12788_1, in12788_2;
    wire c12788;
    assign in12788_1 = {s11218[0]};
    assign in12788_2 = {s11219[0]};
    Full_Adder FA_12788(s12788, c12788, in12788_1, in12788_2, s11217[0]);
    wire[0:0] s12789, in12789_1, in12789_2;
    wire c12789;
    assign in12789_1 = {s11221[0]};
    assign in12789_2 = {s11222[0]};
    Full_Adder FA_12789(s12789, c12789, in12789_1, in12789_2, s11220[0]);
    wire[0:0] s12790, in12790_1, in12790_2;
    wire c12790;
    assign in12790_1 = {s9050[0]};
    assign in12790_2 = {c11215};
    Full_Adder FA_12790(s12790, c12790, in12790_1, in12790_2, s9049[0]);
    wire[0:0] s12791, in12791_1, in12791_2;
    wire c12791;
    assign in12791_1 = {c11217};
    assign in12791_2 = {c11218};
    Full_Adder FA_12791(s12791, c12791, in12791_1, in12791_2, c11216);
    wire[0:0] s12792, in12792_1, in12792_2;
    wire c12792;
    assign in12792_1 = {c11220};
    assign in12792_2 = {c11221};
    Full_Adder FA_12792(s12792, c12792, in12792_1, in12792_2, c11219);
    wire[0:0] s12793, in12793_1, in12793_2;
    wire c12793;
    assign in12793_1 = {s11223[0]};
    assign in12793_2 = {s11224[0]};
    Full_Adder FA_12793(s12793, c12793, in12793_1, in12793_2, c11222);
    wire[0:0] s12794, in12794_1, in12794_2;
    wire c12794;
    assign in12794_1 = {s11226[0]};
    assign in12794_2 = {s11227[0]};
    Full_Adder FA_12794(s12794, c12794, in12794_1, in12794_2, s11225[0]);
    wire[0:0] s12795, in12795_1, in12795_2;
    wire c12795;
    assign in12795_1 = {s11229[0]};
    assign in12795_2 = {s11230[0]};
    Full_Adder FA_12795(s12795, c12795, in12795_1, in12795_2, s11228[0]);
    wire[0:0] s12796, in12796_1, in12796_2;
    wire c12796;
    assign in12796_1 = {s9063[0]};
    assign in12796_2 = {c11223};
    Full_Adder FA_12796(s12796, c12796, in12796_1, in12796_2, s9062[0]);
    wire[0:0] s12797, in12797_1, in12797_2;
    wire c12797;
    assign in12797_1 = {c11225};
    assign in12797_2 = {c11226};
    Full_Adder FA_12797(s12797, c12797, in12797_1, in12797_2, c11224);
    wire[0:0] s12798, in12798_1, in12798_2;
    wire c12798;
    assign in12798_1 = {c11228};
    assign in12798_2 = {c11229};
    Full_Adder FA_12798(s12798, c12798, in12798_1, in12798_2, c11227);
    wire[0:0] s12799, in12799_1, in12799_2;
    wire c12799;
    assign in12799_1 = {s11231[0]};
    assign in12799_2 = {s11232[0]};
    Full_Adder FA_12799(s12799, c12799, in12799_1, in12799_2, c11230);
    wire[0:0] s12800, in12800_1, in12800_2;
    wire c12800;
    assign in12800_1 = {s11234[0]};
    assign in12800_2 = {s11235[0]};
    Full_Adder FA_12800(s12800, c12800, in12800_1, in12800_2, s11233[0]);
    wire[0:0] s12801, in12801_1, in12801_2;
    wire c12801;
    assign in12801_1 = {s11237[0]};
    assign in12801_2 = {s11238[0]};
    Full_Adder FA_12801(s12801, c12801, in12801_1, in12801_2, s11236[0]);
    wire[0:0] s12802, in12802_1, in12802_2;
    wire c12802;
    assign in12802_1 = {s9076[0]};
    assign in12802_2 = {c11231};
    Full_Adder FA_12802(s12802, c12802, in12802_1, in12802_2, s9075[0]);
    wire[0:0] s12803, in12803_1, in12803_2;
    wire c12803;
    assign in12803_1 = {c11233};
    assign in12803_2 = {c11234};
    Full_Adder FA_12803(s12803, c12803, in12803_1, in12803_2, c11232);
    wire[0:0] s12804, in12804_1, in12804_2;
    wire c12804;
    assign in12804_1 = {c11236};
    assign in12804_2 = {c11237};
    Full_Adder FA_12804(s12804, c12804, in12804_1, in12804_2, c11235);
    wire[0:0] s12805, in12805_1, in12805_2;
    wire c12805;
    assign in12805_1 = {s11239[0]};
    assign in12805_2 = {s11240[0]};
    Full_Adder FA_12805(s12805, c12805, in12805_1, in12805_2, c11238);
    wire[0:0] s12806, in12806_1, in12806_2;
    wire c12806;
    assign in12806_1 = {s11242[0]};
    assign in12806_2 = {s11243[0]};
    Full_Adder FA_12806(s12806, c12806, in12806_1, in12806_2, s11241[0]);
    wire[0:0] s12807, in12807_1, in12807_2;
    wire c12807;
    assign in12807_1 = {s11245[0]};
    assign in12807_2 = {s11246[0]};
    Full_Adder FA_12807(s12807, c12807, in12807_1, in12807_2, s11244[0]);
    wire[0:0] s12808, in12808_1, in12808_2;
    wire c12808;
    assign in12808_1 = {s9089[0]};
    assign in12808_2 = {c11239};
    Full_Adder FA_12808(s12808, c12808, in12808_1, in12808_2, s9088[0]);
    wire[0:0] s12809, in12809_1, in12809_2;
    wire c12809;
    assign in12809_1 = {c11241};
    assign in12809_2 = {c11242};
    Full_Adder FA_12809(s12809, c12809, in12809_1, in12809_2, c11240);
    wire[0:0] s12810, in12810_1, in12810_2;
    wire c12810;
    assign in12810_1 = {c11244};
    assign in12810_2 = {c11245};
    Full_Adder FA_12810(s12810, c12810, in12810_1, in12810_2, c11243);
    wire[0:0] s12811, in12811_1, in12811_2;
    wire c12811;
    assign in12811_1 = {s11247[0]};
    assign in12811_2 = {s11248[0]};
    Full_Adder FA_12811(s12811, c12811, in12811_1, in12811_2, c11246);
    wire[0:0] s12812, in12812_1, in12812_2;
    wire c12812;
    assign in12812_1 = {s11250[0]};
    assign in12812_2 = {s11251[0]};
    Full_Adder FA_12812(s12812, c12812, in12812_1, in12812_2, s11249[0]);
    wire[0:0] s12813, in12813_1, in12813_2;
    wire c12813;
    assign in12813_1 = {s11253[0]};
    assign in12813_2 = {s11254[0]};
    Full_Adder FA_12813(s12813, c12813, in12813_1, in12813_2, s11252[0]);
    wire[0:0] s12814, in12814_1, in12814_2;
    wire c12814;
    assign in12814_1 = {s9102[0]};
    assign in12814_2 = {c11247};
    Full_Adder FA_12814(s12814, c12814, in12814_1, in12814_2, s9101[0]);
    wire[0:0] s12815, in12815_1, in12815_2;
    wire c12815;
    assign in12815_1 = {c11249};
    assign in12815_2 = {c11250};
    Full_Adder FA_12815(s12815, c12815, in12815_1, in12815_2, c11248);
    wire[0:0] s12816, in12816_1, in12816_2;
    wire c12816;
    assign in12816_1 = {c11252};
    assign in12816_2 = {c11253};
    Full_Adder FA_12816(s12816, c12816, in12816_1, in12816_2, c11251);
    wire[0:0] s12817, in12817_1, in12817_2;
    wire c12817;
    assign in12817_1 = {s11255[0]};
    assign in12817_2 = {s11256[0]};
    Full_Adder FA_12817(s12817, c12817, in12817_1, in12817_2, c11254);
    wire[0:0] s12818, in12818_1, in12818_2;
    wire c12818;
    assign in12818_1 = {s11258[0]};
    assign in12818_2 = {s11259[0]};
    Full_Adder FA_12818(s12818, c12818, in12818_1, in12818_2, s11257[0]);
    wire[0:0] s12819, in12819_1, in12819_2;
    wire c12819;
    assign in12819_1 = {s11261[0]};
    assign in12819_2 = {s11262[0]};
    Full_Adder FA_12819(s12819, c12819, in12819_1, in12819_2, s11260[0]);
    wire[0:0] s12820, in12820_1, in12820_2;
    wire c12820;
    assign in12820_1 = {s9115[0]};
    assign in12820_2 = {c11255};
    Full_Adder FA_12820(s12820, c12820, in12820_1, in12820_2, s9114[0]);
    wire[0:0] s12821, in12821_1, in12821_2;
    wire c12821;
    assign in12821_1 = {c11257};
    assign in12821_2 = {c11258};
    Full_Adder FA_12821(s12821, c12821, in12821_1, in12821_2, c11256);
    wire[0:0] s12822, in12822_1, in12822_2;
    wire c12822;
    assign in12822_1 = {c11260};
    assign in12822_2 = {c11261};
    Full_Adder FA_12822(s12822, c12822, in12822_1, in12822_2, c11259);
    wire[0:0] s12823, in12823_1, in12823_2;
    wire c12823;
    assign in12823_1 = {s11263[0]};
    assign in12823_2 = {s11264[0]};
    Full_Adder FA_12823(s12823, c12823, in12823_1, in12823_2, c11262);
    wire[0:0] s12824, in12824_1, in12824_2;
    wire c12824;
    assign in12824_1 = {s11266[0]};
    assign in12824_2 = {s11267[0]};
    Full_Adder FA_12824(s12824, c12824, in12824_1, in12824_2, s11265[0]);
    wire[0:0] s12825, in12825_1, in12825_2;
    wire c12825;
    assign in12825_1 = {s11269[0]};
    assign in12825_2 = {s11270[0]};
    Full_Adder FA_12825(s12825, c12825, in12825_1, in12825_2, s11268[0]);
    wire[0:0] s12826, in12826_1, in12826_2;
    wire c12826;
    assign in12826_1 = {s9128[0]};
    assign in12826_2 = {c11263};
    Full_Adder FA_12826(s12826, c12826, in12826_1, in12826_2, s9127[0]);
    wire[0:0] s12827, in12827_1, in12827_2;
    wire c12827;
    assign in12827_1 = {c11265};
    assign in12827_2 = {c11266};
    Full_Adder FA_12827(s12827, c12827, in12827_1, in12827_2, c11264);
    wire[0:0] s12828, in12828_1, in12828_2;
    wire c12828;
    assign in12828_1 = {c11268};
    assign in12828_2 = {c11269};
    Full_Adder FA_12828(s12828, c12828, in12828_1, in12828_2, c11267);
    wire[0:0] s12829, in12829_1, in12829_2;
    wire c12829;
    assign in12829_1 = {s11271[0]};
    assign in12829_2 = {s11272[0]};
    Full_Adder FA_12829(s12829, c12829, in12829_1, in12829_2, c11270);
    wire[0:0] s12830, in12830_1, in12830_2;
    wire c12830;
    assign in12830_1 = {s11274[0]};
    assign in12830_2 = {s11275[0]};
    Full_Adder FA_12830(s12830, c12830, in12830_1, in12830_2, s11273[0]);
    wire[0:0] s12831, in12831_1, in12831_2;
    wire c12831;
    assign in12831_1 = {s11277[0]};
    assign in12831_2 = {s11278[0]};
    Full_Adder FA_12831(s12831, c12831, in12831_1, in12831_2, s11276[0]);
    wire[0:0] s12832, in12832_1, in12832_2;
    wire c12832;
    assign in12832_1 = {s9141[0]};
    assign in12832_2 = {c11271};
    Full_Adder FA_12832(s12832, c12832, in12832_1, in12832_2, s9140[0]);
    wire[0:0] s12833, in12833_1, in12833_2;
    wire c12833;
    assign in12833_1 = {c11273};
    assign in12833_2 = {c11274};
    Full_Adder FA_12833(s12833, c12833, in12833_1, in12833_2, c11272);
    wire[0:0] s12834, in12834_1, in12834_2;
    wire c12834;
    assign in12834_1 = {c11276};
    assign in12834_2 = {c11277};
    Full_Adder FA_12834(s12834, c12834, in12834_1, in12834_2, c11275);
    wire[0:0] s12835, in12835_1, in12835_2;
    wire c12835;
    assign in12835_1 = {s11279[0]};
    assign in12835_2 = {s11280[0]};
    Full_Adder FA_12835(s12835, c12835, in12835_1, in12835_2, c11278);
    wire[0:0] s12836, in12836_1, in12836_2;
    wire c12836;
    assign in12836_1 = {s11282[0]};
    assign in12836_2 = {s11283[0]};
    Full_Adder FA_12836(s12836, c12836, in12836_1, in12836_2, s11281[0]);
    wire[0:0] s12837, in12837_1, in12837_2;
    wire c12837;
    assign in12837_1 = {s11285[0]};
    assign in12837_2 = {s11286[0]};
    Full_Adder FA_12837(s12837, c12837, in12837_1, in12837_2, s11284[0]);
    wire[0:0] s12838, in12838_1, in12838_2;
    wire c12838;
    assign in12838_1 = {s9154[0]};
    assign in12838_2 = {c11279};
    Full_Adder FA_12838(s12838, c12838, in12838_1, in12838_2, s9153[0]);
    wire[0:0] s12839, in12839_1, in12839_2;
    wire c12839;
    assign in12839_1 = {c11281};
    assign in12839_2 = {c11282};
    Full_Adder FA_12839(s12839, c12839, in12839_1, in12839_2, c11280);
    wire[0:0] s12840, in12840_1, in12840_2;
    wire c12840;
    assign in12840_1 = {c11284};
    assign in12840_2 = {c11285};
    Full_Adder FA_12840(s12840, c12840, in12840_1, in12840_2, c11283);
    wire[0:0] s12841, in12841_1, in12841_2;
    wire c12841;
    assign in12841_1 = {s11287[0]};
    assign in12841_2 = {s11288[0]};
    Full_Adder FA_12841(s12841, c12841, in12841_1, in12841_2, c11286);
    wire[0:0] s12842, in12842_1, in12842_2;
    wire c12842;
    assign in12842_1 = {s11290[0]};
    assign in12842_2 = {s11291[0]};
    Full_Adder FA_12842(s12842, c12842, in12842_1, in12842_2, s11289[0]);
    wire[0:0] s12843, in12843_1, in12843_2;
    wire c12843;
    assign in12843_1 = {s11293[0]};
    assign in12843_2 = {s11294[0]};
    Full_Adder FA_12843(s12843, c12843, in12843_1, in12843_2, s11292[0]);
    wire[0:0] s12844, in12844_1, in12844_2;
    wire c12844;
    assign in12844_1 = {s9167[0]};
    assign in12844_2 = {c11287};
    Full_Adder FA_12844(s12844, c12844, in12844_1, in12844_2, s9166[0]);
    wire[0:0] s12845, in12845_1, in12845_2;
    wire c12845;
    assign in12845_1 = {c11289};
    assign in12845_2 = {c11290};
    Full_Adder FA_12845(s12845, c12845, in12845_1, in12845_2, c11288);
    wire[0:0] s12846, in12846_1, in12846_2;
    wire c12846;
    assign in12846_1 = {c11292};
    assign in12846_2 = {c11293};
    Full_Adder FA_12846(s12846, c12846, in12846_1, in12846_2, c11291);
    wire[0:0] s12847, in12847_1, in12847_2;
    wire c12847;
    assign in12847_1 = {s11295[0]};
    assign in12847_2 = {s11296[0]};
    Full_Adder FA_12847(s12847, c12847, in12847_1, in12847_2, c11294);
    wire[0:0] s12848, in12848_1, in12848_2;
    wire c12848;
    assign in12848_1 = {s11298[0]};
    assign in12848_2 = {s11299[0]};
    Full_Adder FA_12848(s12848, c12848, in12848_1, in12848_2, s11297[0]);
    wire[0:0] s12849, in12849_1, in12849_2;
    wire c12849;
    assign in12849_1 = {s11301[0]};
    assign in12849_2 = {s11302[0]};
    Full_Adder FA_12849(s12849, c12849, in12849_1, in12849_2, s11300[0]);
    wire[0:0] s12850, in12850_1, in12850_2;
    wire c12850;
    assign in12850_1 = {s9180[0]};
    assign in12850_2 = {c11295};
    Full_Adder FA_12850(s12850, c12850, in12850_1, in12850_2, s9179[0]);
    wire[0:0] s12851, in12851_1, in12851_2;
    wire c12851;
    assign in12851_1 = {c11297};
    assign in12851_2 = {c11298};
    Full_Adder FA_12851(s12851, c12851, in12851_1, in12851_2, c11296);
    wire[0:0] s12852, in12852_1, in12852_2;
    wire c12852;
    assign in12852_1 = {c11300};
    assign in12852_2 = {c11301};
    Full_Adder FA_12852(s12852, c12852, in12852_1, in12852_2, c11299);
    wire[0:0] s12853, in12853_1, in12853_2;
    wire c12853;
    assign in12853_1 = {s11303[0]};
    assign in12853_2 = {s11304[0]};
    Full_Adder FA_12853(s12853, c12853, in12853_1, in12853_2, c11302);
    wire[0:0] s12854, in12854_1, in12854_2;
    wire c12854;
    assign in12854_1 = {s11306[0]};
    assign in12854_2 = {s11307[0]};
    Full_Adder FA_12854(s12854, c12854, in12854_1, in12854_2, s11305[0]);
    wire[0:0] s12855, in12855_1, in12855_2;
    wire c12855;
    assign in12855_1 = {s11309[0]};
    assign in12855_2 = {s11310[0]};
    Full_Adder FA_12855(s12855, c12855, in12855_1, in12855_2, s11308[0]);
    wire[0:0] s12856, in12856_1, in12856_2;
    wire c12856;
    assign in12856_1 = {s9193[0]};
    assign in12856_2 = {c11303};
    Full_Adder FA_12856(s12856, c12856, in12856_1, in12856_2, s9192[0]);
    wire[0:0] s12857, in12857_1, in12857_2;
    wire c12857;
    assign in12857_1 = {c11305};
    assign in12857_2 = {c11306};
    Full_Adder FA_12857(s12857, c12857, in12857_1, in12857_2, c11304);
    wire[0:0] s12858, in12858_1, in12858_2;
    wire c12858;
    assign in12858_1 = {c11308};
    assign in12858_2 = {c11309};
    Full_Adder FA_12858(s12858, c12858, in12858_1, in12858_2, c11307);
    wire[0:0] s12859, in12859_1, in12859_2;
    wire c12859;
    assign in12859_1 = {s11311[0]};
    assign in12859_2 = {s11312[0]};
    Full_Adder FA_12859(s12859, c12859, in12859_1, in12859_2, c11310);
    wire[0:0] s12860, in12860_1, in12860_2;
    wire c12860;
    assign in12860_1 = {s11314[0]};
    assign in12860_2 = {s11315[0]};
    Full_Adder FA_12860(s12860, c12860, in12860_1, in12860_2, s11313[0]);
    wire[0:0] s12861, in12861_1, in12861_2;
    wire c12861;
    assign in12861_1 = {s11317[0]};
    assign in12861_2 = {s11318[0]};
    Full_Adder FA_12861(s12861, c12861, in12861_1, in12861_2, s11316[0]);
    wire[0:0] s12862, in12862_1, in12862_2;
    wire c12862;
    assign in12862_1 = {s9206[0]};
    assign in12862_2 = {c11311};
    Full_Adder FA_12862(s12862, c12862, in12862_1, in12862_2, s9205[0]);
    wire[0:0] s12863, in12863_1, in12863_2;
    wire c12863;
    assign in12863_1 = {c11313};
    assign in12863_2 = {c11314};
    Full_Adder FA_12863(s12863, c12863, in12863_1, in12863_2, c11312);
    wire[0:0] s12864, in12864_1, in12864_2;
    wire c12864;
    assign in12864_1 = {c11316};
    assign in12864_2 = {c11317};
    Full_Adder FA_12864(s12864, c12864, in12864_1, in12864_2, c11315);
    wire[0:0] s12865, in12865_1, in12865_2;
    wire c12865;
    assign in12865_1 = {s11319[0]};
    assign in12865_2 = {s11320[0]};
    Full_Adder FA_12865(s12865, c12865, in12865_1, in12865_2, c11318);
    wire[0:0] s12866, in12866_1, in12866_2;
    wire c12866;
    assign in12866_1 = {s11322[0]};
    assign in12866_2 = {s11323[0]};
    Full_Adder FA_12866(s12866, c12866, in12866_1, in12866_2, s11321[0]);
    wire[0:0] s12867, in12867_1, in12867_2;
    wire c12867;
    assign in12867_1 = {s11325[0]};
    assign in12867_2 = {s11326[0]};
    Full_Adder FA_12867(s12867, c12867, in12867_1, in12867_2, s11324[0]);
    wire[0:0] s12868, in12868_1, in12868_2;
    wire c12868;
    assign in12868_1 = {s9219[0]};
    assign in12868_2 = {c11319};
    Full_Adder FA_12868(s12868, c12868, in12868_1, in12868_2, s9218[0]);
    wire[0:0] s12869, in12869_1, in12869_2;
    wire c12869;
    assign in12869_1 = {c11321};
    assign in12869_2 = {c11322};
    Full_Adder FA_12869(s12869, c12869, in12869_1, in12869_2, c11320);
    wire[0:0] s12870, in12870_1, in12870_2;
    wire c12870;
    assign in12870_1 = {c11324};
    assign in12870_2 = {c11325};
    Full_Adder FA_12870(s12870, c12870, in12870_1, in12870_2, c11323);
    wire[0:0] s12871, in12871_1, in12871_2;
    wire c12871;
    assign in12871_1 = {s11327[0]};
    assign in12871_2 = {s11328[0]};
    Full_Adder FA_12871(s12871, c12871, in12871_1, in12871_2, c11326);
    wire[0:0] s12872, in12872_1, in12872_2;
    wire c12872;
    assign in12872_1 = {s11330[0]};
    assign in12872_2 = {s11331[0]};
    Full_Adder FA_12872(s12872, c12872, in12872_1, in12872_2, s11329[0]);
    wire[0:0] s12873, in12873_1, in12873_2;
    wire c12873;
    assign in12873_1 = {s11333[0]};
    assign in12873_2 = {s11334[0]};
    Full_Adder FA_12873(s12873, c12873, in12873_1, in12873_2, s11332[0]);
    wire[0:0] s12874, in12874_1, in12874_2;
    wire c12874;
    assign in12874_1 = {s9232[0]};
    assign in12874_2 = {c11327};
    Full_Adder FA_12874(s12874, c12874, in12874_1, in12874_2, s9231[0]);
    wire[0:0] s12875, in12875_1, in12875_2;
    wire c12875;
    assign in12875_1 = {c11329};
    assign in12875_2 = {c11330};
    Full_Adder FA_12875(s12875, c12875, in12875_1, in12875_2, c11328);
    wire[0:0] s12876, in12876_1, in12876_2;
    wire c12876;
    assign in12876_1 = {c11332};
    assign in12876_2 = {c11333};
    Full_Adder FA_12876(s12876, c12876, in12876_1, in12876_2, c11331);
    wire[0:0] s12877, in12877_1, in12877_2;
    wire c12877;
    assign in12877_1 = {s11335[0]};
    assign in12877_2 = {s11336[0]};
    Full_Adder FA_12877(s12877, c12877, in12877_1, in12877_2, c11334);
    wire[0:0] s12878, in12878_1, in12878_2;
    wire c12878;
    assign in12878_1 = {s11338[0]};
    assign in12878_2 = {s11339[0]};
    Full_Adder FA_12878(s12878, c12878, in12878_1, in12878_2, s11337[0]);
    wire[0:0] s12879, in12879_1, in12879_2;
    wire c12879;
    assign in12879_1 = {s11341[0]};
    assign in12879_2 = {s11342[0]};
    Full_Adder FA_12879(s12879, c12879, in12879_1, in12879_2, s11340[0]);
    wire[0:0] s12880, in12880_1, in12880_2;
    wire c12880;
    assign in12880_1 = {s9245[0]};
    assign in12880_2 = {c11335};
    Full_Adder FA_12880(s12880, c12880, in12880_1, in12880_2, s9244[0]);
    wire[0:0] s12881, in12881_1, in12881_2;
    wire c12881;
    assign in12881_1 = {c11337};
    assign in12881_2 = {c11338};
    Full_Adder FA_12881(s12881, c12881, in12881_1, in12881_2, c11336);
    wire[0:0] s12882, in12882_1, in12882_2;
    wire c12882;
    assign in12882_1 = {c11340};
    assign in12882_2 = {c11341};
    Full_Adder FA_12882(s12882, c12882, in12882_1, in12882_2, c11339);
    wire[0:0] s12883, in12883_1, in12883_2;
    wire c12883;
    assign in12883_1 = {s11343[0]};
    assign in12883_2 = {s11344[0]};
    Full_Adder FA_12883(s12883, c12883, in12883_1, in12883_2, c11342);
    wire[0:0] s12884, in12884_1, in12884_2;
    wire c12884;
    assign in12884_1 = {s11346[0]};
    assign in12884_2 = {s11347[0]};
    Full_Adder FA_12884(s12884, c12884, in12884_1, in12884_2, s11345[0]);
    wire[0:0] s12885, in12885_1, in12885_2;
    wire c12885;
    assign in12885_1 = {s11349[0]};
    assign in12885_2 = {s11350[0]};
    Full_Adder FA_12885(s12885, c12885, in12885_1, in12885_2, s11348[0]);
    wire[0:0] s12886, in12886_1, in12886_2;
    wire c12886;
    assign in12886_1 = {s9258[0]};
    assign in12886_2 = {c11343};
    Full_Adder FA_12886(s12886, c12886, in12886_1, in12886_2, s9257[0]);
    wire[0:0] s12887, in12887_1, in12887_2;
    wire c12887;
    assign in12887_1 = {c11345};
    assign in12887_2 = {c11346};
    Full_Adder FA_12887(s12887, c12887, in12887_1, in12887_2, c11344);
    wire[0:0] s12888, in12888_1, in12888_2;
    wire c12888;
    assign in12888_1 = {c11348};
    assign in12888_2 = {c11349};
    Full_Adder FA_12888(s12888, c12888, in12888_1, in12888_2, c11347);
    wire[0:0] s12889, in12889_1, in12889_2;
    wire c12889;
    assign in12889_1 = {s11351[0]};
    assign in12889_2 = {s11352[0]};
    Full_Adder FA_12889(s12889, c12889, in12889_1, in12889_2, c11350);
    wire[0:0] s12890, in12890_1, in12890_2;
    wire c12890;
    assign in12890_1 = {s11354[0]};
    assign in12890_2 = {s11355[0]};
    Full_Adder FA_12890(s12890, c12890, in12890_1, in12890_2, s11353[0]);
    wire[0:0] s12891, in12891_1, in12891_2;
    wire c12891;
    assign in12891_1 = {s11357[0]};
    assign in12891_2 = {s11358[0]};
    Full_Adder FA_12891(s12891, c12891, in12891_1, in12891_2, s11356[0]);
    wire[0:0] s12892, in12892_1, in12892_2;
    wire c12892;
    assign in12892_1 = {s9271[0]};
    assign in12892_2 = {c11351};
    Full_Adder FA_12892(s12892, c12892, in12892_1, in12892_2, s9270[0]);
    wire[0:0] s12893, in12893_1, in12893_2;
    wire c12893;
    assign in12893_1 = {c11353};
    assign in12893_2 = {c11354};
    Full_Adder FA_12893(s12893, c12893, in12893_1, in12893_2, c11352);
    wire[0:0] s12894, in12894_1, in12894_2;
    wire c12894;
    assign in12894_1 = {c11356};
    assign in12894_2 = {c11357};
    Full_Adder FA_12894(s12894, c12894, in12894_1, in12894_2, c11355);
    wire[0:0] s12895, in12895_1, in12895_2;
    wire c12895;
    assign in12895_1 = {s11359[0]};
    assign in12895_2 = {s11360[0]};
    Full_Adder FA_12895(s12895, c12895, in12895_1, in12895_2, c11358);
    wire[0:0] s12896, in12896_1, in12896_2;
    wire c12896;
    assign in12896_1 = {s11362[0]};
    assign in12896_2 = {s11363[0]};
    Full_Adder FA_12896(s12896, c12896, in12896_1, in12896_2, s11361[0]);
    wire[0:0] s12897, in12897_1, in12897_2;
    wire c12897;
    assign in12897_1 = {s11365[0]};
    assign in12897_2 = {s11366[0]};
    Full_Adder FA_12897(s12897, c12897, in12897_1, in12897_2, s11364[0]);
    wire[0:0] s12898, in12898_1, in12898_2;
    wire c12898;
    assign in12898_1 = {s9284[0]};
    assign in12898_2 = {c11359};
    Full_Adder FA_12898(s12898, c12898, in12898_1, in12898_2, s9283[0]);
    wire[0:0] s12899, in12899_1, in12899_2;
    wire c12899;
    assign in12899_1 = {c11361};
    assign in12899_2 = {c11362};
    Full_Adder FA_12899(s12899, c12899, in12899_1, in12899_2, c11360);
    wire[0:0] s12900, in12900_1, in12900_2;
    wire c12900;
    assign in12900_1 = {c11364};
    assign in12900_2 = {c11365};
    Full_Adder FA_12900(s12900, c12900, in12900_1, in12900_2, c11363);
    wire[0:0] s12901, in12901_1, in12901_2;
    wire c12901;
    assign in12901_1 = {s11367[0]};
    assign in12901_2 = {s11368[0]};
    Full_Adder FA_12901(s12901, c12901, in12901_1, in12901_2, c11366);
    wire[0:0] s12902, in12902_1, in12902_2;
    wire c12902;
    assign in12902_1 = {s11370[0]};
    assign in12902_2 = {s11371[0]};
    Full_Adder FA_12902(s12902, c12902, in12902_1, in12902_2, s11369[0]);
    wire[0:0] s12903, in12903_1, in12903_2;
    wire c12903;
    assign in12903_1 = {s11373[0]};
    assign in12903_2 = {s11374[0]};
    Full_Adder FA_12903(s12903, c12903, in12903_1, in12903_2, s11372[0]);
    wire[0:0] s12904, in12904_1, in12904_2;
    wire c12904;
    assign in12904_1 = {s9297[0]};
    assign in12904_2 = {c11367};
    Full_Adder FA_12904(s12904, c12904, in12904_1, in12904_2, s9296[0]);
    wire[0:0] s12905, in12905_1, in12905_2;
    wire c12905;
    assign in12905_1 = {c11369};
    assign in12905_2 = {c11370};
    Full_Adder FA_12905(s12905, c12905, in12905_1, in12905_2, c11368);
    wire[0:0] s12906, in12906_1, in12906_2;
    wire c12906;
    assign in12906_1 = {c11372};
    assign in12906_2 = {c11373};
    Full_Adder FA_12906(s12906, c12906, in12906_1, in12906_2, c11371);
    wire[0:0] s12907, in12907_1, in12907_2;
    wire c12907;
    assign in12907_1 = {s11375[0]};
    assign in12907_2 = {s11376[0]};
    Full_Adder FA_12907(s12907, c12907, in12907_1, in12907_2, c11374);
    wire[0:0] s12908, in12908_1, in12908_2;
    wire c12908;
    assign in12908_1 = {s11378[0]};
    assign in12908_2 = {s11379[0]};
    Full_Adder FA_12908(s12908, c12908, in12908_1, in12908_2, s11377[0]);
    wire[0:0] s12909, in12909_1, in12909_2;
    wire c12909;
    assign in12909_1 = {s11381[0]};
    assign in12909_2 = {s11382[0]};
    Full_Adder FA_12909(s12909, c12909, in12909_1, in12909_2, s11380[0]);
    wire[0:0] s12910, in12910_1, in12910_2;
    wire c12910;
    assign in12910_1 = {s9310[0]};
    assign in12910_2 = {c11375};
    Full_Adder FA_12910(s12910, c12910, in12910_1, in12910_2, s9309[0]);
    wire[0:0] s12911, in12911_1, in12911_2;
    wire c12911;
    assign in12911_1 = {c11377};
    assign in12911_2 = {c11378};
    Full_Adder FA_12911(s12911, c12911, in12911_1, in12911_2, c11376);
    wire[0:0] s12912, in12912_1, in12912_2;
    wire c12912;
    assign in12912_1 = {c11380};
    assign in12912_2 = {c11381};
    Full_Adder FA_12912(s12912, c12912, in12912_1, in12912_2, c11379);
    wire[0:0] s12913, in12913_1, in12913_2;
    wire c12913;
    assign in12913_1 = {s11383[0]};
    assign in12913_2 = {s11384[0]};
    Full_Adder FA_12913(s12913, c12913, in12913_1, in12913_2, c11382);
    wire[0:0] s12914, in12914_1, in12914_2;
    wire c12914;
    assign in12914_1 = {s11386[0]};
    assign in12914_2 = {s11387[0]};
    Full_Adder FA_12914(s12914, c12914, in12914_1, in12914_2, s11385[0]);
    wire[0:0] s12915, in12915_1, in12915_2;
    wire c12915;
    assign in12915_1 = {s11389[0]};
    assign in12915_2 = {s11390[0]};
    Full_Adder FA_12915(s12915, c12915, in12915_1, in12915_2, s11388[0]);
    wire[0:0] s12916, in12916_1, in12916_2;
    wire c12916;
    assign in12916_1 = {s9323[0]};
    assign in12916_2 = {c11383};
    Full_Adder FA_12916(s12916, c12916, in12916_1, in12916_2, s9322[0]);
    wire[0:0] s12917, in12917_1, in12917_2;
    wire c12917;
    assign in12917_1 = {c11385};
    assign in12917_2 = {c11386};
    Full_Adder FA_12917(s12917, c12917, in12917_1, in12917_2, c11384);
    wire[0:0] s12918, in12918_1, in12918_2;
    wire c12918;
    assign in12918_1 = {c11388};
    assign in12918_2 = {c11389};
    Full_Adder FA_12918(s12918, c12918, in12918_1, in12918_2, c11387);
    wire[0:0] s12919, in12919_1, in12919_2;
    wire c12919;
    assign in12919_1 = {s11391[0]};
    assign in12919_2 = {s11392[0]};
    Full_Adder FA_12919(s12919, c12919, in12919_1, in12919_2, c11390);
    wire[0:0] s12920, in12920_1, in12920_2;
    wire c12920;
    assign in12920_1 = {s11394[0]};
    assign in12920_2 = {s11395[0]};
    Full_Adder FA_12920(s12920, c12920, in12920_1, in12920_2, s11393[0]);
    wire[0:0] s12921, in12921_1, in12921_2;
    wire c12921;
    assign in12921_1 = {s11397[0]};
    assign in12921_2 = {s11398[0]};
    Full_Adder FA_12921(s12921, c12921, in12921_1, in12921_2, s11396[0]);
    wire[0:0] s12922, in12922_1, in12922_2;
    wire c12922;
    assign in12922_1 = {s9336[0]};
    assign in12922_2 = {c11391};
    Full_Adder FA_12922(s12922, c12922, in12922_1, in12922_2, s9335[0]);
    wire[0:0] s12923, in12923_1, in12923_2;
    wire c12923;
    assign in12923_1 = {c11393};
    assign in12923_2 = {c11394};
    Full_Adder FA_12923(s12923, c12923, in12923_1, in12923_2, c11392);
    wire[0:0] s12924, in12924_1, in12924_2;
    wire c12924;
    assign in12924_1 = {c11396};
    assign in12924_2 = {c11397};
    Full_Adder FA_12924(s12924, c12924, in12924_1, in12924_2, c11395);
    wire[0:0] s12925, in12925_1, in12925_2;
    wire c12925;
    assign in12925_1 = {s11399[0]};
    assign in12925_2 = {s11400[0]};
    Full_Adder FA_12925(s12925, c12925, in12925_1, in12925_2, c11398);
    wire[0:0] s12926, in12926_1, in12926_2;
    wire c12926;
    assign in12926_1 = {s11402[0]};
    assign in12926_2 = {s11403[0]};
    Full_Adder FA_12926(s12926, c12926, in12926_1, in12926_2, s11401[0]);
    wire[0:0] s12927, in12927_1, in12927_2;
    wire c12927;
    assign in12927_1 = {s11405[0]};
    assign in12927_2 = {s11406[0]};
    Full_Adder FA_12927(s12927, c12927, in12927_1, in12927_2, s11404[0]);
    wire[0:0] s12928, in12928_1, in12928_2;
    wire c12928;
    assign in12928_1 = {s9349[0]};
    assign in12928_2 = {c11399};
    Full_Adder FA_12928(s12928, c12928, in12928_1, in12928_2, s9348[0]);
    wire[0:0] s12929, in12929_1, in12929_2;
    wire c12929;
    assign in12929_1 = {c11401};
    assign in12929_2 = {c11402};
    Full_Adder FA_12929(s12929, c12929, in12929_1, in12929_2, c11400);
    wire[0:0] s12930, in12930_1, in12930_2;
    wire c12930;
    assign in12930_1 = {c11404};
    assign in12930_2 = {c11405};
    Full_Adder FA_12930(s12930, c12930, in12930_1, in12930_2, c11403);
    wire[0:0] s12931, in12931_1, in12931_2;
    wire c12931;
    assign in12931_1 = {s11407[0]};
    assign in12931_2 = {s11408[0]};
    Full_Adder FA_12931(s12931, c12931, in12931_1, in12931_2, c11406);
    wire[0:0] s12932, in12932_1, in12932_2;
    wire c12932;
    assign in12932_1 = {s11410[0]};
    assign in12932_2 = {s11411[0]};
    Full_Adder FA_12932(s12932, c12932, in12932_1, in12932_2, s11409[0]);
    wire[0:0] s12933, in12933_1, in12933_2;
    wire c12933;
    assign in12933_1 = {s11413[0]};
    assign in12933_2 = {s11414[0]};
    Full_Adder FA_12933(s12933, c12933, in12933_1, in12933_2, s11412[0]);
    wire[0:0] s12934, in12934_1, in12934_2;
    wire c12934;
    assign in12934_1 = {s9362[0]};
    assign in12934_2 = {c11407};
    Full_Adder FA_12934(s12934, c12934, in12934_1, in12934_2, s9361[0]);
    wire[0:0] s12935, in12935_1, in12935_2;
    wire c12935;
    assign in12935_1 = {c11409};
    assign in12935_2 = {c11410};
    Full_Adder FA_12935(s12935, c12935, in12935_1, in12935_2, c11408);
    wire[0:0] s12936, in12936_1, in12936_2;
    wire c12936;
    assign in12936_1 = {c11412};
    assign in12936_2 = {c11413};
    Full_Adder FA_12936(s12936, c12936, in12936_1, in12936_2, c11411);
    wire[0:0] s12937, in12937_1, in12937_2;
    wire c12937;
    assign in12937_1 = {s11415[0]};
    assign in12937_2 = {s11416[0]};
    Full_Adder FA_12937(s12937, c12937, in12937_1, in12937_2, c11414);
    wire[0:0] s12938, in12938_1, in12938_2;
    wire c12938;
    assign in12938_1 = {s11418[0]};
    assign in12938_2 = {s11419[0]};
    Full_Adder FA_12938(s12938, c12938, in12938_1, in12938_2, s11417[0]);
    wire[0:0] s12939, in12939_1, in12939_2;
    wire c12939;
    assign in12939_1 = {s11421[0]};
    assign in12939_2 = {s11422[0]};
    Full_Adder FA_12939(s12939, c12939, in12939_1, in12939_2, s11420[0]);
    wire[0:0] s12940, in12940_1, in12940_2;
    wire c12940;
    assign in12940_1 = {s9375[0]};
    assign in12940_2 = {c11415};
    Full_Adder FA_12940(s12940, c12940, in12940_1, in12940_2, s9374[0]);
    wire[0:0] s12941, in12941_1, in12941_2;
    wire c12941;
    assign in12941_1 = {c11417};
    assign in12941_2 = {c11418};
    Full_Adder FA_12941(s12941, c12941, in12941_1, in12941_2, c11416);
    wire[0:0] s12942, in12942_1, in12942_2;
    wire c12942;
    assign in12942_1 = {c11420};
    assign in12942_2 = {c11421};
    Full_Adder FA_12942(s12942, c12942, in12942_1, in12942_2, c11419);
    wire[0:0] s12943, in12943_1, in12943_2;
    wire c12943;
    assign in12943_1 = {s11423[0]};
    assign in12943_2 = {s11424[0]};
    Full_Adder FA_12943(s12943, c12943, in12943_1, in12943_2, c11422);
    wire[0:0] s12944, in12944_1, in12944_2;
    wire c12944;
    assign in12944_1 = {s11426[0]};
    assign in12944_2 = {s11427[0]};
    Full_Adder FA_12944(s12944, c12944, in12944_1, in12944_2, s11425[0]);
    wire[0:0] s12945, in12945_1, in12945_2;
    wire c12945;
    assign in12945_1 = {s11429[0]};
    assign in12945_2 = {s11430[0]};
    Full_Adder FA_12945(s12945, c12945, in12945_1, in12945_2, s11428[0]);
    wire[0:0] s12946, in12946_1, in12946_2;
    wire c12946;
    assign in12946_1 = {s9388[0]};
    assign in12946_2 = {c11423};
    Full_Adder FA_12946(s12946, c12946, in12946_1, in12946_2, s9387[0]);
    wire[0:0] s12947, in12947_1, in12947_2;
    wire c12947;
    assign in12947_1 = {c11425};
    assign in12947_2 = {c11426};
    Full_Adder FA_12947(s12947, c12947, in12947_1, in12947_2, c11424);
    wire[0:0] s12948, in12948_1, in12948_2;
    wire c12948;
    assign in12948_1 = {c11428};
    assign in12948_2 = {c11429};
    Full_Adder FA_12948(s12948, c12948, in12948_1, in12948_2, c11427);
    wire[0:0] s12949, in12949_1, in12949_2;
    wire c12949;
    assign in12949_1 = {s11431[0]};
    assign in12949_2 = {s11432[0]};
    Full_Adder FA_12949(s12949, c12949, in12949_1, in12949_2, c11430);
    wire[0:0] s12950, in12950_1, in12950_2;
    wire c12950;
    assign in12950_1 = {s11434[0]};
    assign in12950_2 = {s11435[0]};
    Full_Adder FA_12950(s12950, c12950, in12950_1, in12950_2, s11433[0]);
    wire[0:0] s12951, in12951_1, in12951_2;
    wire c12951;
    assign in12951_1 = {s11437[0]};
    assign in12951_2 = {s11438[0]};
    Full_Adder FA_12951(s12951, c12951, in12951_1, in12951_2, s11436[0]);
    wire[0:0] s12952, in12952_1, in12952_2;
    wire c12952;
    assign in12952_1 = {s9401[0]};
    assign in12952_2 = {c11431};
    Full_Adder FA_12952(s12952, c12952, in12952_1, in12952_2, s9400[0]);
    wire[0:0] s12953, in12953_1, in12953_2;
    wire c12953;
    assign in12953_1 = {c11433};
    assign in12953_2 = {c11434};
    Full_Adder FA_12953(s12953, c12953, in12953_1, in12953_2, c11432);
    wire[0:0] s12954, in12954_1, in12954_2;
    wire c12954;
    assign in12954_1 = {c11436};
    assign in12954_2 = {c11437};
    Full_Adder FA_12954(s12954, c12954, in12954_1, in12954_2, c11435);
    wire[0:0] s12955, in12955_1, in12955_2;
    wire c12955;
    assign in12955_1 = {s11439[0]};
    assign in12955_2 = {s11440[0]};
    Full_Adder FA_12955(s12955, c12955, in12955_1, in12955_2, c11438);
    wire[0:0] s12956, in12956_1, in12956_2;
    wire c12956;
    assign in12956_1 = {s11442[0]};
    assign in12956_2 = {s11443[0]};
    Full_Adder FA_12956(s12956, c12956, in12956_1, in12956_2, s11441[0]);
    wire[0:0] s12957, in12957_1, in12957_2;
    wire c12957;
    assign in12957_1 = {s11445[0]};
    assign in12957_2 = {s11446[0]};
    Full_Adder FA_12957(s12957, c12957, in12957_1, in12957_2, s11444[0]);
    wire[0:0] s12958, in12958_1, in12958_2;
    wire c12958;
    assign in12958_1 = {s9414[0]};
    assign in12958_2 = {c11439};
    Full_Adder FA_12958(s12958, c12958, in12958_1, in12958_2, s9413[0]);
    wire[0:0] s12959, in12959_1, in12959_2;
    wire c12959;
    assign in12959_1 = {c11441};
    assign in12959_2 = {c11442};
    Full_Adder FA_12959(s12959, c12959, in12959_1, in12959_2, c11440);
    wire[0:0] s12960, in12960_1, in12960_2;
    wire c12960;
    assign in12960_1 = {c11444};
    assign in12960_2 = {c11445};
    Full_Adder FA_12960(s12960, c12960, in12960_1, in12960_2, c11443);
    wire[0:0] s12961, in12961_1, in12961_2;
    wire c12961;
    assign in12961_1 = {s11447[0]};
    assign in12961_2 = {s11448[0]};
    Full_Adder FA_12961(s12961, c12961, in12961_1, in12961_2, c11446);
    wire[0:0] s12962, in12962_1, in12962_2;
    wire c12962;
    assign in12962_1 = {s11450[0]};
    assign in12962_2 = {s11451[0]};
    Full_Adder FA_12962(s12962, c12962, in12962_1, in12962_2, s11449[0]);
    wire[0:0] s12963, in12963_1, in12963_2;
    wire c12963;
    assign in12963_1 = {s11453[0]};
    assign in12963_2 = {s11454[0]};
    Full_Adder FA_12963(s12963, c12963, in12963_1, in12963_2, s11452[0]);
    wire[0:0] s12964, in12964_1, in12964_2;
    wire c12964;
    assign in12964_1 = {s9427[0]};
    assign in12964_2 = {c11447};
    Full_Adder FA_12964(s12964, c12964, in12964_1, in12964_2, s9426[0]);
    wire[0:0] s12965, in12965_1, in12965_2;
    wire c12965;
    assign in12965_1 = {c11449};
    assign in12965_2 = {c11450};
    Full_Adder FA_12965(s12965, c12965, in12965_1, in12965_2, c11448);
    wire[0:0] s12966, in12966_1, in12966_2;
    wire c12966;
    assign in12966_1 = {c11452};
    assign in12966_2 = {c11453};
    Full_Adder FA_12966(s12966, c12966, in12966_1, in12966_2, c11451);
    wire[0:0] s12967, in12967_1, in12967_2;
    wire c12967;
    assign in12967_1 = {s11455[0]};
    assign in12967_2 = {s11456[0]};
    Full_Adder FA_12967(s12967, c12967, in12967_1, in12967_2, c11454);
    wire[0:0] s12968, in12968_1, in12968_2;
    wire c12968;
    assign in12968_1 = {s11458[0]};
    assign in12968_2 = {s11459[0]};
    Full_Adder FA_12968(s12968, c12968, in12968_1, in12968_2, s11457[0]);
    wire[0:0] s12969, in12969_1, in12969_2;
    wire c12969;
    assign in12969_1 = {s11461[0]};
    assign in12969_2 = {s11462[0]};
    Full_Adder FA_12969(s12969, c12969, in12969_1, in12969_2, s11460[0]);
    wire[0:0] s12970, in12970_1, in12970_2;
    wire c12970;
    assign in12970_1 = {s9440[0]};
    assign in12970_2 = {c11455};
    Full_Adder FA_12970(s12970, c12970, in12970_1, in12970_2, s9439[0]);
    wire[0:0] s12971, in12971_1, in12971_2;
    wire c12971;
    assign in12971_1 = {c11457};
    assign in12971_2 = {c11458};
    Full_Adder FA_12971(s12971, c12971, in12971_1, in12971_2, c11456);
    wire[0:0] s12972, in12972_1, in12972_2;
    wire c12972;
    assign in12972_1 = {c11460};
    assign in12972_2 = {c11461};
    Full_Adder FA_12972(s12972, c12972, in12972_1, in12972_2, c11459);
    wire[0:0] s12973, in12973_1, in12973_2;
    wire c12973;
    assign in12973_1 = {s11463[0]};
    assign in12973_2 = {s11464[0]};
    Full_Adder FA_12973(s12973, c12973, in12973_1, in12973_2, c11462);
    wire[0:0] s12974, in12974_1, in12974_2;
    wire c12974;
    assign in12974_1 = {s11466[0]};
    assign in12974_2 = {s11467[0]};
    Full_Adder FA_12974(s12974, c12974, in12974_1, in12974_2, s11465[0]);
    wire[0:0] s12975, in12975_1, in12975_2;
    wire c12975;
    assign in12975_1 = {s11469[0]};
    assign in12975_2 = {s11470[0]};
    Full_Adder FA_12975(s12975, c12975, in12975_1, in12975_2, s11468[0]);
    wire[0:0] s12976, in12976_1, in12976_2;
    wire c12976;
    assign in12976_1 = {s9453[0]};
    assign in12976_2 = {c11463};
    Full_Adder FA_12976(s12976, c12976, in12976_1, in12976_2, s9452[0]);
    wire[0:0] s12977, in12977_1, in12977_2;
    wire c12977;
    assign in12977_1 = {c11465};
    assign in12977_2 = {c11466};
    Full_Adder FA_12977(s12977, c12977, in12977_1, in12977_2, c11464);
    wire[0:0] s12978, in12978_1, in12978_2;
    wire c12978;
    assign in12978_1 = {c11468};
    assign in12978_2 = {c11469};
    Full_Adder FA_12978(s12978, c12978, in12978_1, in12978_2, c11467);
    wire[0:0] s12979, in12979_1, in12979_2;
    wire c12979;
    assign in12979_1 = {s11471[0]};
    assign in12979_2 = {s11472[0]};
    Full_Adder FA_12979(s12979, c12979, in12979_1, in12979_2, c11470);
    wire[0:0] s12980, in12980_1, in12980_2;
    wire c12980;
    assign in12980_1 = {s11474[0]};
    assign in12980_2 = {s11475[0]};
    Full_Adder FA_12980(s12980, c12980, in12980_1, in12980_2, s11473[0]);
    wire[0:0] s12981, in12981_1, in12981_2;
    wire c12981;
    assign in12981_1 = {s11477[0]};
    assign in12981_2 = {s11478[0]};
    Full_Adder FA_12981(s12981, c12981, in12981_1, in12981_2, s11476[0]);
    wire[0:0] s12982, in12982_1, in12982_2;
    wire c12982;
    assign in12982_1 = {s9466[0]};
    assign in12982_2 = {c11471};
    Full_Adder FA_12982(s12982, c12982, in12982_1, in12982_2, s9465[0]);
    wire[0:0] s12983, in12983_1, in12983_2;
    wire c12983;
    assign in12983_1 = {c11473};
    assign in12983_2 = {c11474};
    Full_Adder FA_12983(s12983, c12983, in12983_1, in12983_2, c11472);
    wire[0:0] s12984, in12984_1, in12984_2;
    wire c12984;
    assign in12984_1 = {c11476};
    assign in12984_2 = {c11477};
    Full_Adder FA_12984(s12984, c12984, in12984_1, in12984_2, c11475);
    wire[0:0] s12985, in12985_1, in12985_2;
    wire c12985;
    assign in12985_1 = {s11479[0]};
    assign in12985_2 = {s11480[0]};
    Full_Adder FA_12985(s12985, c12985, in12985_1, in12985_2, c11478);
    wire[0:0] s12986, in12986_1, in12986_2;
    wire c12986;
    assign in12986_1 = {s11482[0]};
    assign in12986_2 = {s11483[0]};
    Full_Adder FA_12986(s12986, c12986, in12986_1, in12986_2, s11481[0]);
    wire[0:0] s12987, in12987_1, in12987_2;
    wire c12987;
    assign in12987_1 = {s11485[0]};
    assign in12987_2 = {s11486[0]};
    Full_Adder FA_12987(s12987, c12987, in12987_1, in12987_2, s11484[0]);
    wire[0:0] s12988, in12988_1, in12988_2;
    wire c12988;
    assign in12988_1 = {s9479[0]};
    assign in12988_2 = {c11479};
    Full_Adder FA_12988(s12988, c12988, in12988_1, in12988_2, s9478[0]);
    wire[0:0] s12989, in12989_1, in12989_2;
    wire c12989;
    assign in12989_1 = {c11481};
    assign in12989_2 = {c11482};
    Full_Adder FA_12989(s12989, c12989, in12989_1, in12989_2, c11480);
    wire[0:0] s12990, in12990_1, in12990_2;
    wire c12990;
    assign in12990_1 = {c11484};
    assign in12990_2 = {c11485};
    Full_Adder FA_12990(s12990, c12990, in12990_1, in12990_2, c11483);
    wire[0:0] s12991, in12991_1, in12991_2;
    wire c12991;
    assign in12991_1 = {s11487[0]};
    assign in12991_2 = {s11488[0]};
    Full_Adder FA_12991(s12991, c12991, in12991_1, in12991_2, c11486);
    wire[0:0] s12992, in12992_1, in12992_2;
    wire c12992;
    assign in12992_1 = {s11490[0]};
    assign in12992_2 = {s11491[0]};
    Full_Adder FA_12992(s12992, c12992, in12992_1, in12992_2, s11489[0]);
    wire[0:0] s12993, in12993_1, in12993_2;
    wire c12993;
    assign in12993_1 = {s11493[0]};
    assign in12993_2 = {s11494[0]};
    Full_Adder FA_12993(s12993, c12993, in12993_1, in12993_2, s11492[0]);
    wire[0:0] s12994, in12994_1, in12994_2;
    wire c12994;
    assign in12994_1 = {s9492[0]};
    assign in12994_2 = {c11487};
    Full_Adder FA_12994(s12994, c12994, in12994_1, in12994_2, s9491[0]);
    wire[0:0] s12995, in12995_1, in12995_2;
    wire c12995;
    assign in12995_1 = {c11489};
    assign in12995_2 = {c11490};
    Full_Adder FA_12995(s12995, c12995, in12995_1, in12995_2, c11488);
    wire[0:0] s12996, in12996_1, in12996_2;
    wire c12996;
    assign in12996_1 = {c11492};
    assign in12996_2 = {c11493};
    Full_Adder FA_12996(s12996, c12996, in12996_1, in12996_2, c11491);
    wire[0:0] s12997, in12997_1, in12997_2;
    wire c12997;
    assign in12997_1 = {s11495[0]};
    assign in12997_2 = {s11496[0]};
    Full_Adder FA_12997(s12997, c12997, in12997_1, in12997_2, c11494);
    wire[0:0] s12998, in12998_1, in12998_2;
    wire c12998;
    assign in12998_1 = {s11498[0]};
    assign in12998_2 = {s11499[0]};
    Full_Adder FA_12998(s12998, c12998, in12998_1, in12998_2, s11497[0]);
    wire[0:0] s12999, in12999_1, in12999_2;
    wire c12999;
    assign in12999_1 = {s11501[0]};
    assign in12999_2 = {s11502[0]};
    Full_Adder FA_12999(s12999, c12999, in12999_1, in12999_2, s11500[0]);
    wire[0:0] s13000, in13000_1, in13000_2;
    wire c13000;
    assign in13000_1 = {s9505[0]};
    assign in13000_2 = {c11495};
    Full_Adder FA_13000(s13000, c13000, in13000_1, in13000_2, s9504[0]);
    wire[0:0] s13001, in13001_1, in13001_2;
    wire c13001;
    assign in13001_1 = {c11497};
    assign in13001_2 = {c11498};
    Full_Adder FA_13001(s13001, c13001, in13001_1, in13001_2, c11496);
    wire[0:0] s13002, in13002_1, in13002_2;
    wire c13002;
    assign in13002_1 = {c11500};
    assign in13002_2 = {c11501};
    Full_Adder FA_13002(s13002, c13002, in13002_1, in13002_2, c11499);
    wire[0:0] s13003, in13003_1, in13003_2;
    wire c13003;
    assign in13003_1 = {s11503[0]};
    assign in13003_2 = {s11504[0]};
    Full_Adder FA_13003(s13003, c13003, in13003_1, in13003_2, c11502);
    wire[0:0] s13004, in13004_1, in13004_2;
    wire c13004;
    assign in13004_1 = {s11506[0]};
    assign in13004_2 = {s11507[0]};
    Full_Adder FA_13004(s13004, c13004, in13004_1, in13004_2, s11505[0]);
    wire[0:0] s13005, in13005_1, in13005_2;
    wire c13005;
    assign in13005_1 = {s11509[0]};
    assign in13005_2 = {s11510[0]};
    Full_Adder FA_13005(s13005, c13005, in13005_1, in13005_2, s11508[0]);
    wire[0:0] s13006, in13006_1, in13006_2;
    wire c13006;
    assign in13006_1 = {s9518[0]};
    assign in13006_2 = {c11503};
    Full_Adder FA_13006(s13006, c13006, in13006_1, in13006_2, s9517[0]);
    wire[0:0] s13007, in13007_1, in13007_2;
    wire c13007;
    assign in13007_1 = {c11505};
    assign in13007_2 = {c11506};
    Full_Adder FA_13007(s13007, c13007, in13007_1, in13007_2, c11504);
    wire[0:0] s13008, in13008_1, in13008_2;
    wire c13008;
    assign in13008_1 = {c11508};
    assign in13008_2 = {c11509};
    Full_Adder FA_13008(s13008, c13008, in13008_1, in13008_2, c11507);
    wire[0:0] s13009, in13009_1, in13009_2;
    wire c13009;
    assign in13009_1 = {s11511[0]};
    assign in13009_2 = {s11512[0]};
    Full_Adder FA_13009(s13009, c13009, in13009_1, in13009_2, c11510);
    wire[0:0] s13010, in13010_1, in13010_2;
    wire c13010;
    assign in13010_1 = {s11514[0]};
    assign in13010_2 = {s11515[0]};
    Full_Adder FA_13010(s13010, c13010, in13010_1, in13010_2, s11513[0]);
    wire[0:0] s13011, in13011_1, in13011_2;
    wire c13011;
    assign in13011_1 = {s11517[0]};
    assign in13011_2 = {s11518[0]};
    Full_Adder FA_13011(s13011, c13011, in13011_1, in13011_2, s11516[0]);
    wire[0:0] s13012, in13012_1, in13012_2;
    wire c13012;
    assign in13012_1 = {s9531[0]};
    assign in13012_2 = {c11511};
    Full_Adder FA_13012(s13012, c13012, in13012_1, in13012_2, s9530[0]);
    wire[0:0] s13013, in13013_1, in13013_2;
    wire c13013;
    assign in13013_1 = {c11513};
    assign in13013_2 = {c11514};
    Full_Adder FA_13013(s13013, c13013, in13013_1, in13013_2, c11512);
    wire[0:0] s13014, in13014_1, in13014_2;
    wire c13014;
    assign in13014_1 = {c11516};
    assign in13014_2 = {c11517};
    Full_Adder FA_13014(s13014, c13014, in13014_1, in13014_2, c11515);
    wire[0:0] s13015, in13015_1, in13015_2;
    wire c13015;
    assign in13015_1 = {s11519[0]};
    assign in13015_2 = {s11520[0]};
    Full_Adder FA_13015(s13015, c13015, in13015_1, in13015_2, c11518);
    wire[0:0] s13016, in13016_1, in13016_2;
    wire c13016;
    assign in13016_1 = {s11522[0]};
    assign in13016_2 = {s11523[0]};
    Full_Adder FA_13016(s13016, c13016, in13016_1, in13016_2, s11521[0]);
    wire[0:0] s13017, in13017_1, in13017_2;
    wire c13017;
    assign in13017_1 = {s11525[0]};
    assign in13017_2 = {s11526[0]};
    Full_Adder FA_13017(s13017, c13017, in13017_1, in13017_2, s11524[0]);
    wire[0:0] s13018, in13018_1, in13018_2;
    wire c13018;
    assign in13018_1 = {s9544[0]};
    assign in13018_2 = {c11519};
    Full_Adder FA_13018(s13018, c13018, in13018_1, in13018_2, s9543[0]);
    wire[0:0] s13019, in13019_1, in13019_2;
    wire c13019;
    assign in13019_1 = {c11521};
    assign in13019_2 = {c11522};
    Full_Adder FA_13019(s13019, c13019, in13019_1, in13019_2, c11520);
    wire[0:0] s13020, in13020_1, in13020_2;
    wire c13020;
    assign in13020_1 = {c11524};
    assign in13020_2 = {c11525};
    Full_Adder FA_13020(s13020, c13020, in13020_1, in13020_2, c11523);
    wire[0:0] s13021, in13021_1, in13021_2;
    wire c13021;
    assign in13021_1 = {s11527[0]};
    assign in13021_2 = {s11528[0]};
    Full_Adder FA_13021(s13021, c13021, in13021_1, in13021_2, c11526);
    wire[0:0] s13022, in13022_1, in13022_2;
    wire c13022;
    assign in13022_1 = {s11530[0]};
    assign in13022_2 = {s11531[0]};
    Full_Adder FA_13022(s13022, c13022, in13022_1, in13022_2, s11529[0]);
    wire[0:0] s13023, in13023_1, in13023_2;
    wire c13023;
    assign in13023_1 = {s11533[0]};
    assign in13023_2 = {s11534[0]};
    Full_Adder FA_13023(s13023, c13023, in13023_1, in13023_2, s11532[0]);
    wire[0:0] s13024, in13024_1, in13024_2;
    wire c13024;
    assign in13024_1 = {s9557[0]};
    assign in13024_2 = {c11527};
    Full_Adder FA_13024(s13024, c13024, in13024_1, in13024_2, s9556[0]);
    wire[0:0] s13025, in13025_1, in13025_2;
    wire c13025;
    assign in13025_1 = {c11529};
    assign in13025_2 = {c11530};
    Full_Adder FA_13025(s13025, c13025, in13025_1, in13025_2, c11528);
    wire[0:0] s13026, in13026_1, in13026_2;
    wire c13026;
    assign in13026_1 = {c11532};
    assign in13026_2 = {c11533};
    Full_Adder FA_13026(s13026, c13026, in13026_1, in13026_2, c11531);
    wire[0:0] s13027, in13027_1, in13027_2;
    wire c13027;
    assign in13027_1 = {s11535[0]};
    assign in13027_2 = {s11536[0]};
    Full_Adder FA_13027(s13027, c13027, in13027_1, in13027_2, c11534);
    wire[0:0] s13028, in13028_1, in13028_2;
    wire c13028;
    assign in13028_1 = {s11538[0]};
    assign in13028_2 = {s11539[0]};
    Full_Adder FA_13028(s13028, c13028, in13028_1, in13028_2, s11537[0]);
    wire[0:0] s13029, in13029_1, in13029_2;
    wire c13029;
    assign in13029_1 = {s11541[0]};
    assign in13029_2 = {s11542[0]};
    Full_Adder FA_13029(s13029, c13029, in13029_1, in13029_2, s11540[0]);
    wire[0:0] s13030, in13030_1, in13030_2;
    wire c13030;
    assign in13030_1 = {s9570[0]};
    assign in13030_2 = {c11535};
    Full_Adder FA_13030(s13030, c13030, in13030_1, in13030_2, s9569[0]);
    wire[0:0] s13031, in13031_1, in13031_2;
    wire c13031;
    assign in13031_1 = {c11537};
    assign in13031_2 = {c11538};
    Full_Adder FA_13031(s13031, c13031, in13031_1, in13031_2, c11536);
    wire[0:0] s13032, in13032_1, in13032_2;
    wire c13032;
    assign in13032_1 = {c11540};
    assign in13032_2 = {c11541};
    Full_Adder FA_13032(s13032, c13032, in13032_1, in13032_2, c11539);
    wire[0:0] s13033, in13033_1, in13033_2;
    wire c13033;
    assign in13033_1 = {s11543[0]};
    assign in13033_2 = {s11544[0]};
    Full_Adder FA_13033(s13033, c13033, in13033_1, in13033_2, c11542);
    wire[0:0] s13034, in13034_1, in13034_2;
    wire c13034;
    assign in13034_1 = {s11546[0]};
    assign in13034_2 = {s11547[0]};
    Full_Adder FA_13034(s13034, c13034, in13034_1, in13034_2, s11545[0]);
    wire[0:0] s13035, in13035_1, in13035_2;
    wire c13035;
    assign in13035_1 = {s11549[0]};
    assign in13035_2 = {s11550[0]};
    Full_Adder FA_13035(s13035, c13035, in13035_1, in13035_2, s11548[0]);
    wire[0:0] s13036, in13036_1, in13036_2;
    wire c13036;
    assign in13036_1 = {s9583[0]};
    assign in13036_2 = {c11543};
    Full_Adder FA_13036(s13036, c13036, in13036_1, in13036_2, s9582[0]);
    wire[0:0] s13037, in13037_1, in13037_2;
    wire c13037;
    assign in13037_1 = {c11545};
    assign in13037_2 = {c11546};
    Full_Adder FA_13037(s13037, c13037, in13037_1, in13037_2, c11544);
    wire[0:0] s13038, in13038_1, in13038_2;
    wire c13038;
    assign in13038_1 = {c11548};
    assign in13038_2 = {c11549};
    Full_Adder FA_13038(s13038, c13038, in13038_1, in13038_2, c11547);
    wire[0:0] s13039, in13039_1, in13039_2;
    wire c13039;
    assign in13039_1 = {s11551[0]};
    assign in13039_2 = {s11552[0]};
    Full_Adder FA_13039(s13039, c13039, in13039_1, in13039_2, c11550);
    wire[0:0] s13040, in13040_1, in13040_2;
    wire c13040;
    assign in13040_1 = {s11554[0]};
    assign in13040_2 = {s11555[0]};
    Full_Adder FA_13040(s13040, c13040, in13040_1, in13040_2, s11553[0]);
    wire[0:0] s13041, in13041_1, in13041_2;
    wire c13041;
    assign in13041_1 = {s11557[0]};
    assign in13041_2 = {s11558[0]};
    Full_Adder FA_13041(s13041, c13041, in13041_1, in13041_2, s11556[0]);
    wire[0:0] s13042, in13042_1, in13042_2;
    wire c13042;
    assign in13042_1 = {s9596[0]};
    assign in13042_2 = {c11551};
    Full_Adder FA_13042(s13042, c13042, in13042_1, in13042_2, s9595[0]);
    wire[0:0] s13043, in13043_1, in13043_2;
    wire c13043;
    assign in13043_1 = {c11553};
    assign in13043_2 = {c11554};
    Full_Adder FA_13043(s13043, c13043, in13043_1, in13043_2, c11552);
    wire[0:0] s13044, in13044_1, in13044_2;
    wire c13044;
    assign in13044_1 = {c11556};
    assign in13044_2 = {c11557};
    Full_Adder FA_13044(s13044, c13044, in13044_1, in13044_2, c11555);
    wire[0:0] s13045, in13045_1, in13045_2;
    wire c13045;
    assign in13045_1 = {s11559[0]};
    assign in13045_2 = {s11560[0]};
    Full_Adder FA_13045(s13045, c13045, in13045_1, in13045_2, c11558);
    wire[0:0] s13046, in13046_1, in13046_2;
    wire c13046;
    assign in13046_1 = {s11562[0]};
    assign in13046_2 = {s11563[0]};
    Full_Adder FA_13046(s13046, c13046, in13046_1, in13046_2, s11561[0]);
    wire[0:0] s13047, in13047_1, in13047_2;
    wire c13047;
    assign in13047_1 = {s11565[0]};
    assign in13047_2 = {s11566[0]};
    Full_Adder FA_13047(s13047, c13047, in13047_1, in13047_2, s11564[0]);
    wire[0:0] s13048, in13048_1, in13048_2;
    wire c13048;
    assign in13048_1 = {s9609[0]};
    assign in13048_2 = {c11559};
    Full_Adder FA_13048(s13048, c13048, in13048_1, in13048_2, s9608[0]);
    wire[0:0] s13049, in13049_1, in13049_2;
    wire c13049;
    assign in13049_1 = {c11561};
    assign in13049_2 = {c11562};
    Full_Adder FA_13049(s13049, c13049, in13049_1, in13049_2, c11560);
    wire[0:0] s13050, in13050_1, in13050_2;
    wire c13050;
    assign in13050_1 = {c11564};
    assign in13050_2 = {c11565};
    Full_Adder FA_13050(s13050, c13050, in13050_1, in13050_2, c11563);
    wire[0:0] s13051, in13051_1, in13051_2;
    wire c13051;
    assign in13051_1 = {s11567[0]};
    assign in13051_2 = {s11568[0]};
    Full_Adder FA_13051(s13051, c13051, in13051_1, in13051_2, c11566);
    wire[0:0] s13052, in13052_1, in13052_2;
    wire c13052;
    assign in13052_1 = {s11570[0]};
    assign in13052_2 = {s11571[0]};
    Full_Adder FA_13052(s13052, c13052, in13052_1, in13052_2, s11569[0]);
    wire[0:0] s13053, in13053_1, in13053_2;
    wire c13053;
    assign in13053_1 = {s11573[0]};
    assign in13053_2 = {s11574[0]};
    Full_Adder FA_13053(s13053, c13053, in13053_1, in13053_2, s11572[0]);
    wire[0:0] s13054, in13054_1, in13054_2;
    wire c13054;
    assign in13054_1 = {s9622[0]};
    assign in13054_2 = {c11567};
    Full_Adder FA_13054(s13054, c13054, in13054_1, in13054_2, s9621[0]);
    wire[0:0] s13055, in13055_1, in13055_2;
    wire c13055;
    assign in13055_1 = {c11569};
    assign in13055_2 = {c11570};
    Full_Adder FA_13055(s13055, c13055, in13055_1, in13055_2, c11568);
    wire[0:0] s13056, in13056_1, in13056_2;
    wire c13056;
    assign in13056_1 = {c11572};
    assign in13056_2 = {c11573};
    Full_Adder FA_13056(s13056, c13056, in13056_1, in13056_2, c11571);
    wire[0:0] s13057, in13057_1, in13057_2;
    wire c13057;
    assign in13057_1 = {s11575[0]};
    assign in13057_2 = {s11576[0]};
    Full_Adder FA_13057(s13057, c13057, in13057_1, in13057_2, c11574);
    wire[0:0] s13058, in13058_1, in13058_2;
    wire c13058;
    assign in13058_1 = {s11578[0]};
    assign in13058_2 = {s11579[0]};
    Full_Adder FA_13058(s13058, c13058, in13058_1, in13058_2, s11577[0]);
    wire[0:0] s13059, in13059_1, in13059_2;
    wire c13059;
    assign in13059_1 = {s11581[0]};
    assign in13059_2 = {s11582[0]};
    Full_Adder FA_13059(s13059, c13059, in13059_1, in13059_2, s11580[0]);
    wire[0:0] s13060, in13060_1, in13060_2;
    wire c13060;
    assign in13060_1 = {s9635[0]};
    assign in13060_2 = {c11575};
    Full_Adder FA_13060(s13060, c13060, in13060_1, in13060_2, s9634[0]);
    wire[0:0] s13061, in13061_1, in13061_2;
    wire c13061;
    assign in13061_1 = {c11577};
    assign in13061_2 = {c11578};
    Full_Adder FA_13061(s13061, c13061, in13061_1, in13061_2, c11576);
    wire[0:0] s13062, in13062_1, in13062_2;
    wire c13062;
    assign in13062_1 = {c11580};
    assign in13062_2 = {c11581};
    Full_Adder FA_13062(s13062, c13062, in13062_1, in13062_2, c11579);
    wire[0:0] s13063, in13063_1, in13063_2;
    wire c13063;
    assign in13063_1 = {s11583[0]};
    assign in13063_2 = {s11584[0]};
    Full_Adder FA_13063(s13063, c13063, in13063_1, in13063_2, c11582);
    wire[0:0] s13064, in13064_1, in13064_2;
    wire c13064;
    assign in13064_1 = {s11586[0]};
    assign in13064_2 = {s11587[0]};
    Full_Adder FA_13064(s13064, c13064, in13064_1, in13064_2, s11585[0]);
    wire[0:0] s13065, in13065_1, in13065_2;
    wire c13065;
    assign in13065_1 = {s11589[0]};
    assign in13065_2 = {s11590[0]};
    Full_Adder FA_13065(s13065, c13065, in13065_1, in13065_2, s11588[0]);
    wire[0:0] s13066, in13066_1, in13066_2;
    wire c13066;
    assign in13066_1 = {s9648[0]};
    assign in13066_2 = {c11583};
    Full_Adder FA_13066(s13066, c13066, in13066_1, in13066_2, s9647[0]);
    wire[0:0] s13067, in13067_1, in13067_2;
    wire c13067;
    assign in13067_1 = {c11585};
    assign in13067_2 = {c11586};
    Full_Adder FA_13067(s13067, c13067, in13067_1, in13067_2, c11584);
    wire[0:0] s13068, in13068_1, in13068_2;
    wire c13068;
    assign in13068_1 = {c11588};
    assign in13068_2 = {c11589};
    Full_Adder FA_13068(s13068, c13068, in13068_1, in13068_2, c11587);
    wire[0:0] s13069, in13069_1, in13069_2;
    wire c13069;
    assign in13069_1 = {s11591[0]};
    assign in13069_2 = {s11592[0]};
    Full_Adder FA_13069(s13069, c13069, in13069_1, in13069_2, c11590);
    wire[0:0] s13070, in13070_1, in13070_2;
    wire c13070;
    assign in13070_1 = {s11594[0]};
    assign in13070_2 = {s11595[0]};
    Full_Adder FA_13070(s13070, c13070, in13070_1, in13070_2, s11593[0]);
    wire[0:0] s13071, in13071_1, in13071_2;
    wire c13071;
    assign in13071_1 = {s11597[0]};
    assign in13071_2 = {s11598[0]};
    Full_Adder FA_13071(s13071, c13071, in13071_1, in13071_2, s11596[0]);
    wire[0:0] s13072, in13072_1, in13072_2;
    wire c13072;
    assign in13072_1 = {s9661[0]};
    assign in13072_2 = {c11591};
    Full_Adder FA_13072(s13072, c13072, in13072_1, in13072_2, s9660[0]);
    wire[0:0] s13073, in13073_1, in13073_2;
    wire c13073;
    assign in13073_1 = {c11593};
    assign in13073_2 = {c11594};
    Full_Adder FA_13073(s13073, c13073, in13073_1, in13073_2, c11592);
    wire[0:0] s13074, in13074_1, in13074_2;
    wire c13074;
    assign in13074_1 = {c11596};
    assign in13074_2 = {c11597};
    Full_Adder FA_13074(s13074, c13074, in13074_1, in13074_2, c11595);
    wire[0:0] s13075, in13075_1, in13075_2;
    wire c13075;
    assign in13075_1 = {s11599[0]};
    assign in13075_2 = {s11600[0]};
    Full_Adder FA_13075(s13075, c13075, in13075_1, in13075_2, c11598);
    wire[0:0] s13076, in13076_1, in13076_2;
    wire c13076;
    assign in13076_1 = {s11602[0]};
    assign in13076_2 = {s11603[0]};
    Full_Adder FA_13076(s13076, c13076, in13076_1, in13076_2, s11601[0]);
    wire[0:0] s13077, in13077_1, in13077_2;
    wire c13077;
    assign in13077_1 = {s11605[0]};
    assign in13077_2 = {s11606[0]};
    Full_Adder FA_13077(s13077, c13077, in13077_1, in13077_2, s11604[0]);
    wire[0:0] s13078, in13078_1, in13078_2;
    wire c13078;
    assign in13078_1 = {s9674[0]};
    assign in13078_2 = {c11599};
    Full_Adder FA_13078(s13078, c13078, in13078_1, in13078_2, s9673[0]);
    wire[0:0] s13079, in13079_1, in13079_2;
    wire c13079;
    assign in13079_1 = {c11601};
    assign in13079_2 = {c11602};
    Full_Adder FA_13079(s13079, c13079, in13079_1, in13079_2, c11600);
    wire[0:0] s13080, in13080_1, in13080_2;
    wire c13080;
    assign in13080_1 = {c11604};
    assign in13080_2 = {c11605};
    Full_Adder FA_13080(s13080, c13080, in13080_1, in13080_2, c11603);
    wire[0:0] s13081, in13081_1, in13081_2;
    wire c13081;
    assign in13081_1 = {s11607[0]};
    assign in13081_2 = {s11608[0]};
    Full_Adder FA_13081(s13081, c13081, in13081_1, in13081_2, c11606);
    wire[0:0] s13082, in13082_1, in13082_2;
    wire c13082;
    assign in13082_1 = {s11610[0]};
    assign in13082_2 = {s11611[0]};
    Full_Adder FA_13082(s13082, c13082, in13082_1, in13082_2, s11609[0]);
    wire[0:0] s13083, in13083_1, in13083_2;
    wire c13083;
    assign in13083_1 = {s11613[0]};
    assign in13083_2 = {s11614[0]};
    Full_Adder FA_13083(s13083, c13083, in13083_1, in13083_2, s11612[0]);
    wire[0:0] s13084, in13084_1, in13084_2;
    wire c13084;
    assign in13084_1 = {s9687[0]};
    assign in13084_2 = {c11607};
    Full_Adder FA_13084(s13084, c13084, in13084_1, in13084_2, s9686[0]);
    wire[0:0] s13085, in13085_1, in13085_2;
    wire c13085;
    assign in13085_1 = {c11609};
    assign in13085_2 = {c11610};
    Full_Adder FA_13085(s13085, c13085, in13085_1, in13085_2, c11608);
    wire[0:0] s13086, in13086_1, in13086_2;
    wire c13086;
    assign in13086_1 = {c11612};
    assign in13086_2 = {c11613};
    Full_Adder FA_13086(s13086, c13086, in13086_1, in13086_2, c11611);
    wire[0:0] s13087, in13087_1, in13087_2;
    wire c13087;
    assign in13087_1 = {s11615[0]};
    assign in13087_2 = {s11616[0]};
    Full_Adder FA_13087(s13087, c13087, in13087_1, in13087_2, c11614);
    wire[0:0] s13088, in13088_1, in13088_2;
    wire c13088;
    assign in13088_1 = {s11618[0]};
    assign in13088_2 = {s11619[0]};
    Full_Adder FA_13088(s13088, c13088, in13088_1, in13088_2, s11617[0]);
    wire[0:0] s13089, in13089_1, in13089_2;
    wire c13089;
    assign in13089_1 = {s11621[0]};
    assign in13089_2 = {s11622[0]};
    Full_Adder FA_13089(s13089, c13089, in13089_1, in13089_2, s11620[0]);
    wire[0:0] s13090, in13090_1, in13090_2;
    wire c13090;
    assign in13090_1 = {s9700[0]};
    assign in13090_2 = {c11615};
    Full_Adder FA_13090(s13090, c13090, in13090_1, in13090_2, s9699[0]);
    wire[0:0] s13091, in13091_1, in13091_2;
    wire c13091;
    assign in13091_1 = {c11617};
    assign in13091_2 = {c11618};
    Full_Adder FA_13091(s13091, c13091, in13091_1, in13091_2, c11616);
    wire[0:0] s13092, in13092_1, in13092_2;
    wire c13092;
    assign in13092_1 = {c11620};
    assign in13092_2 = {c11621};
    Full_Adder FA_13092(s13092, c13092, in13092_1, in13092_2, c11619);
    wire[0:0] s13093, in13093_1, in13093_2;
    wire c13093;
    assign in13093_1 = {s11623[0]};
    assign in13093_2 = {s11624[0]};
    Full_Adder FA_13093(s13093, c13093, in13093_1, in13093_2, c11622);
    wire[0:0] s13094, in13094_1, in13094_2;
    wire c13094;
    assign in13094_1 = {s11626[0]};
    assign in13094_2 = {s11627[0]};
    Full_Adder FA_13094(s13094, c13094, in13094_1, in13094_2, s11625[0]);
    wire[0:0] s13095, in13095_1, in13095_2;
    wire c13095;
    assign in13095_1 = {s11629[0]};
    assign in13095_2 = {s11630[0]};
    Full_Adder FA_13095(s13095, c13095, in13095_1, in13095_2, s11628[0]);
    wire[0:0] s13096, in13096_1, in13096_2;
    wire c13096;
    assign in13096_1 = {s9713[0]};
    assign in13096_2 = {c11623};
    Full_Adder FA_13096(s13096, c13096, in13096_1, in13096_2, s9712[0]);
    wire[0:0] s13097, in13097_1, in13097_2;
    wire c13097;
    assign in13097_1 = {c11625};
    assign in13097_2 = {c11626};
    Full_Adder FA_13097(s13097, c13097, in13097_1, in13097_2, c11624);
    wire[0:0] s13098, in13098_1, in13098_2;
    wire c13098;
    assign in13098_1 = {c11628};
    assign in13098_2 = {c11629};
    Full_Adder FA_13098(s13098, c13098, in13098_1, in13098_2, c11627);
    wire[0:0] s13099, in13099_1, in13099_2;
    wire c13099;
    assign in13099_1 = {s11631[0]};
    assign in13099_2 = {s11632[0]};
    Full_Adder FA_13099(s13099, c13099, in13099_1, in13099_2, c11630);
    wire[0:0] s13100, in13100_1, in13100_2;
    wire c13100;
    assign in13100_1 = {s11634[0]};
    assign in13100_2 = {s11635[0]};
    Full_Adder FA_13100(s13100, c13100, in13100_1, in13100_2, s11633[0]);
    wire[0:0] s13101, in13101_1, in13101_2;
    wire c13101;
    assign in13101_1 = {s11637[0]};
    assign in13101_2 = {s11638[0]};
    Full_Adder FA_13101(s13101, c13101, in13101_1, in13101_2, s11636[0]);
    wire[0:0] s13102, in13102_1, in13102_2;
    wire c13102;
    assign in13102_1 = {s9726[0]};
    assign in13102_2 = {c11631};
    Full_Adder FA_13102(s13102, c13102, in13102_1, in13102_2, s9725[0]);
    wire[0:0] s13103, in13103_1, in13103_2;
    wire c13103;
    assign in13103_1 = {c11633};
    assign in13103_2 = {c11634};
    Full_Adder FA_13103(s13103, c13103, in13103_1, in13103_2, c11632);
    wire[0:0] s13104, in13104_1, in13104_2;
    wire c13104;
    assign in13104_1 = {c11636};
    assign in13104_2 = {c11637};
    Full_Adder FA_13104(s13104, c13104, in13104_1, in13104_2, c11635);
    wire[0:0] s13105, in13105_1, in13105_2;
    wire c13105;
    assign in13105_1 = {s11639[0]};
    assign in13105_2 = {s11640[0]};
    Full_Adder FA_13105(s13105, c13105, in13105_1, in13105_2, c11638);
    wire[0:0] s13106, in13106_1, in13106_2;
    wire c13106;
    assign in13106_1 = {s11642[0]};
    assign in13106_2 = {s11643[0]};
    Full_Adder FA_13106(s13106, c13106, in13106_1, in13106_2, s11641[0]);
    wire[0:0] s13107, in13107_1, in13107_2;
    wire c13107;
    assign in13107_1 = {s11645[0]};
    assign in13107_2 = {s11646[0]};
    Full_Adder FA_13107(s13107, c13107, in13107_1, in13107_2, s11644[0]);
    wire[0:0] s13108, in13108_1, in13108_2;
    wire c13108;
    assign in13108_1 = {s9739[0]};
    assign in13108_2 = {c11639};
    Full_Adder FA_13108(s13108, c13108, in13108_1, in13108_2, s9738[0]);
    wire[0:0] s13109, in13109_1, in13109_2;
    wire c13109;
    assign in13109_1 = {c11641};
    assign in13109_2 = {c11642};
    Full_Adder FA_13109(s13109, c13109, in13109_1, in13109_2, c11640);
    wire[0:0] s13110, in13110_1, in13110_2;
    wire c13110;
    assign in13110_1 = {c11644};
    assign in13110_2 = {c11645};
    Full_Adder FA_13110(s13110, c13110, in13110_1, in13110_2, c11643);
    wire[0:0] s13111, in13111_1, in13111_2;
    wire c13111;
    assign in13111_1 = {s11647[0]};
    assign in13111_2 = {s11648[0]};
    Full_Adder FA_13111(s13111, c13111, in13111_1, in13111_2, c11646);
    wire[0:0] s13112, in13112_1, in13112_2;
    wire c13112;
    assign in13112_1 = {s11650[0]};
    assign in13112_2 = {s11651[0]};
    Full_Adder FA_13112(s13112, c13112, in13112_1, in13112_2, s11649[0]);
    wire[0:0] s13113, in13113_1, in13113_2;
    wire c13113;
    assign in13113_1 = {s11653[0]};
    assign in13113_2 = {s11654[0]};
    Full_Adder FA_13113(s13113, c13113, in13113_1, in13113_2, s11652[0]);
    wire[0:0] s13114, in13114_1, in13114_2;
    wire c13114;
    assign in13114_1 = {s9752[0]};
    assign in13114_2 = {c11647};
    Full_Adder FA_13114(s13114, c13114, in13114_1, in13114_2, s9751[0]);
    wire[0:0] s13115, in13115_1, in13115_2;
    wire c13115;
    assign in13115_1 = {c11649};
    assign in13115_2 = {c11650};
    Full_Adder FA_13115(s13115, c13115, in13115_1, in13115_2, c11648);
    wire[0:0] s13116, in13116_1, in13116_2;
    wire c13116;
    assign in13116_1 = {c11652};
    assign in13116_2 = {c11653};
    Full_Adder FA_13116(s13116, c13116, in13116_1, in13116_2, c11651);
    wire[0:0] s13117, in13117_1, in13117_2;
    wire c13117;
    assign in13117_1 = {s11655[0]};
    assign in13117_2 = {s11656[0]};
    Full_Adder FA_13117(s13117, c13117, in13117_1, in13117_2, c11654);
    wire[0:0] s13118, in13118_1, in13118_2;
    wire c13118;
    assign in13118_1 = {s11658[0]};
    assign in13118_2 = {s11659[0]};
    Full_Adder FA_13118(s13118, c13118, in13118_1, in13118_2, s11657[0]);
    wire[0:0] s13119, in13119_1, in13119_2;
    wire c13119;
    assign in13119_1 = {s11661[0]};
    assign in13119_2 = {s11662[0]};
    Full_Adder FA_13119(s13119, c13119, in13119_1, in13119_2, s11660[0]);
    wire[0:0] s13120, in13120_1, in13120_2;
    wire c13120;
    assign in13120_1 = {s9765[0]};
    assign in13120_2 = {c11655};
    Full_Adder FA_13120(s13120, c13120, in13120_1, in13120_2, s9764[0]);
    wire[0:0] s13121, in13121_1, in13121_2;
    wire c13121;
    assign in13121_1 = {c11657};
    assign in13121_2 = {c11658};
    Full_Adder FA_13121(s13121, c13121, in13121_1, in13121_2, c11656);
    wire[0:0] s13122, in13122_1, in13122_2;
    wire c13122;
    assign in13122_1 = {c11660};
    assign in13122_2 = {c11661};
    Full_Adder FA_13122(s13122, c13122, in13122_1, in13122_2, c11659);
    wire[0:0] s13123, in13123_1, in13123_2;
    wire c13123;
    assign in13123_1 = {s11663[0]};
    assign in13123_2 = {s11664[0]};
    Full_Adder FA_13123(s13123, c13123, in13123_1, in13123_2, c11662);
    wire[0:0] s13124, in13124_1, in13124_2;
    wire c13124;
    assign in13124_1 = {s11666[0]};
    assign in13124_2 = {s11667[0]};
    Full_Adder FA_13124(s13124, c13124, in13124_1, in13124_2, s11665[0]);
    wire[0:0] s13125, in13125_1, in13125_2;
    wire c13125;
    assign in13125_1 = {s11669[0]};
    assign in13125_2 = {s11670[0]};
    Full_Adder FA_13125(s13125, c13125, in13125_1, in13125_2, s11668[0]);
    wire[0:0] s13126, in13126_1, in13126_2;
    wire c13126;
    assign in13126_1 = {s9778[0]};
    assign in13126_2 = {c11663};
    Full_Adder FA_13126(s13126, c13126, in13126_1, in13126_2, s9777[0]);
    wire[0:0] s13127, in13127_1, in13127_2;
    wire c13127;
    assign in13127_1 = {c11665};
    assign in13127_2 = {c11666};
    Full_Adder FA_13127(s13127, c13127, in13127_1, in13127_2, c11664);
    wire[0:0] s13128, in13128_1, in13128_2;
    wire c13128;
    assign in13128_1 = {c11668};
    assign in13128_2 = {c11669};
    Full_Adder FA_13128(s13128, c13128, in13128_1, in13128_2, c11667);
    wire[0:0] s13129, in13129_1, in13129_2;
    wire c13129;
    assign in13129_1 = {s11671[0]};
    assign in13129_2 = {s11672[0]};
    Full_Adder FA_13129(s13129, c13129, in13129_1, in13129_2, c11670);
    wire[0:0] s13130, in13130_1, in13130_2;
    wire c13130;
    assign in13130_1 = {s11674[0]};
    assign in13130_2 = {s11675[0]};
    Full_Adder FA_13130(s13130, c13130, in13130_1, in13130_2, s11673[0]);
    wire[0:0] s13131, in13131_1, in13131_2;
    wire c13131;
    assign in13131_1 = {s11677[0]};
    assign in13131_2 = {s11678[0]};
    Full_Adder FA_13131(s13131, c13131, in13131_1, in13131_2, s11676[0]);
    wire[0:0] s13132, in13132_1, in13132_2;
    wire c13132;
    assign in13132_1 = {s9791[0]};
    assign in13132_2 = {c11671};
    Full_Adder FA_13132(s13132, c13132, in13132_1, in13132_2, s9790[0]);
    wire[0:0] s13133, in13133_1, in13133_2;
    wire c13133;
    assign in13133_1 = {c11673};
    assign in13133_2 = {c11674};
    Full_Adder FA_13133(s13133, c13133, in13133_1, in13133_2, c11672);
    wire[0:0] s13134, in13134_1, in13134_2;
    wire c13134;
    assign in13134_1 = {c11676};
    assign in13134_2 = {c11677};
    Full_Adder FA_13134(s13134, c13134, in13134_1, in13134_2, c11675);
    wire[0:0] s13135, in13135_1, in13135_2;
    wire c13135;
    assign in13135_1 = {s11679[0]};
    assign in13135_2 = {s11680[0]};
    Full_Adder FA_13135(s13135, c13135, in13135_1, in13135_2, c11678);
    wire[0:0] s13136, in13136_1, in13136_2;
    wire c13136;
    assign in13136_1 = {s11682[0]};
    assign in13136_2 = {s11683[0]};
    Full_Adder FA_13136(s13136, c13136, in13136_1, in13136_2, s11681[0]);
    wire[0:0] s13137, in13137_1, in13137_2;
    wire c13137;
    assign in13137_1 = {s11685[0]};
    assign in13137_2 = {s11686[0]};
    Full_Adder FA_13137(s13137, c13137, in13137_1, in13137_2, s11684[0]);
    wire[0:0] s13138, in13138_1, in13138_2;
    wire c13138;
    assign in13138_1 = {s9804[0]};
    assign in13138_2 = {c11679};
    Full_Adder FA_13138(s13138, c13138, in13138_1, in13138_2, s9803[0]);
    wire[0:0] s13139, in13139_1, in13139_2;
    wire c13139;
    assign in13139_1 = {c11681};
    assign in13139_2 = {c11682};
    Full_Adder FA_13139(s13139, c13139, in13139_1, in13139_2, c11680);
    wire[0:0] s13140, in13140_1, in13140_2;
    wire c13140;
    assign in13140_1 = {c11684};
    assign in13140_2 = {c11685};
    Full_Adder FA_13140(s13140, c13140, in13140_1, in13140_2, c11683);
    wire[0:0] s13141, in13141_1, in13141_2;
    wire c13141;
    assign in13141_1 = {s11687[0]};
    assign in13141_2 = {s11688[0]};
    Full_Adder FA_13141(s13141, c13141, in13141_1, in13141_2, c11686);
    wire[0:0] s13142, in13142_1, in13142_2;
    wire c13142;
    assign in13142_1 = {s11690[0]};
    assign in13142_2 = {s11691[0]};
    Full_Adder FA_13142(s13142, c13142, in13142_1, in13142_2, s11689[0]);
    wire[0:0] s13143, in13143_1, in13143_2;
    wire c13143;
    assign in13143_1 = {s11693[0]};
    assign in13143_2 = {s11694[0]};
    Full_Adder FA_13143(s13143, c13143, in13143_1, in13143_2, s11692[0]);
    wire[0:0] s13144, in13144_1, in13144_2;
    wire c13144;
    assign in13144_1 = {s9817[0]};
    assign in13144_2 = {c11687};
    Full_Adder FA_13144(s13144, c13144, in13144_1, in13144_2, s9816[0]);
    wire[0:0] s13145, in13145_1, in13145_2;
    wire c13145;
    assign in13145_1 = {c11689};
    assign in13145_2 = {c11690};
    Full_Adder FA_13145(s13145, c13145, in13145_1, in13145_2, c11688);
    wire[0:0] s13146, in13146_1, in13146_2;
    wire c13146;
    assign in13146_1 = {c11692};
    assign in13146_2 = {c11693};
    Full_Adder FA_13146(s13146, c13146, in13146_1, in13146_2, c11691);
    wire[0:0] s13147, in13147_1, in13147_2;
    wire c13147;
    assign in13147_1 = {s11695[0]};
    assign in13147_2 = {s11696[0]};
    Full_Adder FA_13147(s13147, c13147, in13147_1, in13147_2, c11694);
    wire[0:0] s13148, in13148_1, in13148_2;
    wire c13148;
    assign in13148_1 = {s11698[0]};
    assign in13148_2 = {s11699[0]};
    Full_Adder FA_13148(s13148, c13148, in13148_1, in13148_2, s11697[0]);
    wire[0:0] s13149, in13149_1, in13149_2;
    wire c13149;
    assign in13149_1 = {s11701[0]};
    assign in13149_2 = {s11702[0]};
    Full_Adder FA_13149(s13149, c13149, in13149_1, in13149_2, s11700[0]);
    wire[0:0] s13150, in13150_1, in13150_2;
    wire c13150;
    assign in13150_1 = {s9830[0]};
    assign in13150_2 = {c11695};
    Full_Adder FA_13150(s13150, c13150, in13150_1, in13150_2, s9829[0]);
    wire[0:0] s13151, in13151_1, in13151_2;
    wire c13151;
    assign in13151_1 = {c11697};
    assign in13151_2 = {c11698};
    Full_Adder FA_13151(s13151, c13151, in13151_1, in13151_2, c11696);
    wire[0:0] s13152, in13152_1, in13152_2;
    wire c13152;
    assign in13152_1 = {c11700};
    assign in13152_2 = {c11701};
    Full_Adder FA_13152(s13152, c13152, in13152_1, in13152_2, c11699);
    wire[0:0] s13153, in13153_1, in13153_2;
    wire c13153;
    assign in13153_1 = {s11703[0]};
    assign in13153_2 = {s11704[0]};
    Full_Adder FA_13153(s13153, c13153, in13153_1, in13153_2, c11702);
    wire[0:0] s13154, in13154_1, in13154_2;
    wire c13154;
    assign in13154_1 = {s11706[0]};
    assign in13154_2 = {s11707[0]};
    Full_Adder FA_13154(s13154, c13154, in13154_1, in13154_2, s11705[0]);
    wire[0:0] s13155, in13155_1, in13155_2;
    wire c13155;
    assign in13155_1 = {s11709[0]};
    assign in13155_2 = {s11710[0]};
    Full_Adder FA_13155(s13155, c13155, in13155_1, in13155_2, s11708[0]);
    wire[0:0] s13156, in13156_1, in13156_2;
    wire c13156;
    assign in13156_1 = {s9843[0]};
    assign in13156_2 = {c11703};
    Full_Adder FA_13156(s13156, c13156, in13156_1, in13156_2, s9842[0]);
    wire[0:0] s13157, in13157_1, in13157_2;
    wire c13157;
    assign in13157_1 = {c11705};
    assign in13157_2 = {c11706};
    Full_Adder FA_13157(s13157, c13157, in13157_1, in13157_2, c11704);
    wire[0:0] s13158, in13158_1, in13158_2;
    wire c13158;
    assign in13158_1 = {c11708};
    assign in13158_2 = {c11709};
    Full_Adder FA_13158(s13158, c13158, in13158_1, in13158_2, c11707);
    wire[0:0] s13159, in13159_1, in13159_2;
    wire c13159;
    assign in13159_1 = {s11711[0]};
    assign in13159_2 = {s11712[0]};
    Full_Adder FA_13159(s13159, c13159, in13159_1, in13159_2, c11710);
    wire[0:0] s13160, in13160_1, in13160_2;
    wire c13160;
    assign in13160_1 = {s11714[0]};
    assign in13160_2 = {s11715[0]};
    Full_Adder FA_13160(s13160, c13160, in13160_1, in13160_2, s11713[0]);
    wire[0:0] s13161, in13161_1, in13161_2;
    wire c13161;
    assign in13161_1 = {s11717[0]};
    assign in13161_2 = {s11718[0]};
    Full_Adder FA_13161(s13161, c13161, in13161_1, in13161_2, s11716[0]);
    wire[0:0] s13162, in13162_1, in13162_2;
    wire c13162;
    assign in13162_1 = {s9856[0]};
    assign in13162_2 = {c11711};
    Full_Adder FA_13162(s13162, c13162, in13162_1, in13162_2, s9855[0]);
    wire[0:0] s13163, in13163_1, in13163_2;
    wire c13163;
    assign in13163_1 = {c11713};
    assign in13163_2 = {c11714};
    Full_Adder FA_13163(s13163, c13163, in13163_1, in13163_2, c11712);
    wire[0:0] s13164, in13164_1, in13164_2;
    wire c13164;
    assign in13164_1 = {c11716};
    assign in13164_2 = {c11717};
    Full_Adder FA_13164(s13164, c13164, in13164_1, in13164_2, c11715);
    wire[0:0] s13165, in13165_1, in13165_2;
    wire c13165;
    assign in13165_1 = {s11719[0]};
    assign in13165_2 = {s11720[0]};
    Full_Adder FA_13165(s13165, c13165, in13165_1, in13165_2, c11718);
    wire[0:0] s13166, in13166_1, in13166_2;
    wire c13166;
    assign in13166_1 = {s11722[0]};
    assign in13166_2 = {s11723[0]};
    Full_Adder FA_13166(s13166, c13166, in13166_1, in13166_2, s11721[0]);
    wire[0:0] s13167, in13167_1, in13167_2;
    wire c13167;
    assign in13167_1 = {s11725[0]};
    assign in13167_2 = {s11726[0]};
    Full_Adder FA_13167(s13167, c13167, in13167_1, in13167_2, s11724[0]);
    wire[0:0] s13168, in13168_1, in13168_2;
    wire c13168;
    assign in13168_1 = {s9869[0]};
    assign in13168_2 = {c11719};
    Full_Adder FA_13168(s13168, c13168, in13168_1, in13168_2, s9868[0]);
    wire[0:0] s13169, in13169_1, in13169_2;
    wire c13169;
    assign in13169_1 = {c11721};
    assign in13169_2 = {c11722};
    Full_Adder FA_13169(s13169, c13169, in13169_1, in13169_2, c11720);
    wire[0:0] s13170, in13170_1, in13170_2;
    wire c13170;
    assign in13170_1 = {c11724};
    assign in13170_2 = {c11725};
    Full_Adder FA_13170(s13170, c13170, in13170_1, in13170_2, c11723);
    wire[0:0] s13171, in13171_1, in13171_2;
    wire c13171;
    assign in13171_1 = {s11727[0]};
    assign in13171_2 = {s11728[0]};
    Full_Adder FA_13171(s13171, c13171, in13171_1, in13171_2, c11726);
    wire[0:0] s13172, in13172_1, in13172_2;
    wire c13172;
    assign in13172_1 = {s11730[0]};
    assign in13172_2 = {s11731[0]};
    Full_Adder FA_13172(s13172, c13172, in13172_1, in13172_2, s11729[0]);
    wire[0:0] s13173, in13173_1, in13173_2;
    wire c13173;
    assign in13173_1 = {s11733[0]};
    assign in13173_2 = {s11734[0]};
    Full_Adder FA_13173(s13173, c13173, in13173_1, in13173_2, s11732[0]);
    wire[0:0] s13174, in13174_1, in13174_2;
    wire c13174;
    assign in13174_1 = {s9882[0]};
    assign in13174_2 = {c11727};
    Full_Adder FA_13174(s13174, c13174, in13174_1, in13174_2, s9881[0]);
    wire[0:0] s13175, in13175_1, in13175_2;
    wire c13175;
    assign in13175_1 = {c11729};
    assign in13175_2 = {c11730};
    Full_Adder FA_13175(s13175, c13175, in13175_1, in13175_2, c11728);
    wire[0:0] s13176, in13176_1, in13176_2;
    wire c13176;
    assign in13176_1 = {c11732};
    assign in13176_2 = {c11733};
    Full_Adder FA_13176(s13176, c13176, in13176_1, in13176_2, c11731);
    wire[0:0] s13177, in13177_1, in13177_2;
    wire c13177;
    assign in13177_1 = {s11735[0]};
    assign in13177_2 = {s11736[0]};
    Full_Adder FA_13177(s13177, c13177, in13177_1, in13177_2, c11734);
    wire[0:0] s13178, in13178_1, in13178_2;
    wire c13178;
    assign in13178_1 = {s11738[0]};
    assign in13178_2 = {s11739[0]};
    Full_Adder FA_13178(s13178, c13178, in13178_1, in13178_2, s11737[0]);
    wire[0:0] s13179, in13179_1, in13179_2;
    wire c13179;
    assign in13179_1 = {s11741[0]};
    assign in13179_2 = {s11742[0]};
    Full_Adder FA_13179(s13179, c13179, in13179_1, in13179_2, s11740[0]);
    wire[0:0] s13180, in13180_1, in13180_2;
    wire c13180;
    assign in13180_1 = {s9895[0]};
    assign in13180_2 = {c11735};
    Full_Adder FA_13180(s13180, c13180, in13180_1, in13180_2, s9894[0]);
    wire[0:0] s13181, in13181_1, in13181_2;
    wire c13181;
    assign in13181_1 = {c11737};
    assign in13181_2 = {c11738};
    Full_Adder FA_13181(s13181, c13181, in13181_1, in13181_2, c11736);
    wire[0:0] s13182, in13182_1, in13182_2;
    wire c13182;
    assign in13182_1 = {c11740};
    assign in13182_2 = {c11741};
    Full_Adder FA_13182(s13182, c13182, in13182_1, in13182_2, c11739);
    wire[0:0] s13183, in13183_1, in13183_2;
    wire c13183;
    assign in13183_1 = {s11743[0]};
    assign in13183_2 = {s11744[0]};
    Full_Adder FA_13183(s13183, c13183, in13183_1, in13183_2, c11742);
    wire[0:0] s13184, in13184_1, in13184_2;
    wire c13184;
    assign in13184_1 = {s11746[0]};
    assign in13184_2 = {s11747[0]};
    Full_Adder FA_13184(s13184, c13184, in13184_1, in13184_2, s11745[0]);
    wire[0:0] s13185, in13185_1, in13185_2;
    wire c13185;
    assign in13185_1 = {s11749[0]};
    assign in13185_2 = {s11750[0]};
    Full_Adder FA_13185(s13185, c13185, in13185_1, in13185_2, s11748[0]);
    wire[0:0] s13186, in13186_1, in13186_2;
    wire c13186;
    assign in13186_1 = {s9908[0]};
    assign in13186_2 = {c11743};
    Full_Adder FA_13186(s13186, c13186, in13186_1, in13186_2, s9907[0]);
    wire[0:0] s13187, in13187_1, in13187_2;
    wire c13187;
    assign in13187_1 = {c11745};
    assign in13187_2 = {c11746};
    Full_Adder FA_13187(s13187, c13187, in13187_1, in13187_2, c11744);
    wire[0:0] s13188, in13188_1, in13188_2;
    wire c13188;
    assign in13188_1 = {c11748};
    assign in13188_2 = {c11749};
    Full_Adder FA_13188(s13188, c13188, in13188_1, in13188_2, c11747);
    wire[0:0] s13189, in13189_1, in13189_2;
    wire c13189;
    assign in13189_1 = {s11751[0]};
    assign in13189_2 = {s11752[0]};
    Full_Adder FA_13189(s13189, c13189, in13189_1, in13189_2, c11750);
    wire[0:0] s13190, in13190_1, in13190_2;
    wire c13190;
    assign in13190_1 = {s11754[0]};
    assign in13190_2 = {s11755[0]};
    Full_Adder FA_13190(s13190, c13190, in13190_1, in13190_2, s11753[0]);
    wire[0:0] s13191, in13191_1, in13191_2;
    wire c13191;
    assign in13191_1 = {s11757[0]};
    assign in13191_2 = {s11758[0]};
    Full_Adder FA_13191(s13191, c13191, in13191_1, in13191_2, s11756[0]);
    wire[0:0] s13192, in13192_1, in13192_2;
    wire c13192;
    assign in13192_1 = {s9921[0]};
    assign in13192_2 = {c11751};
    Full_Adder FA_13192(s13192, c13192, in13192_1, in13192_2, s9920[0]);
    wire[0:0] s13193, in13193_1, in13193_2;
    wire c13193;
    assign in13193_1 = {c11753};
    assign in13193_2 = {c11754};
    Full_Adder FA_13193(s13193, c13193, in13193_1, in13193_2, c11752);
    wire[0:0] s13194, in13194_1, in13194_2;
    wire c13194;
    assign in13194_1 = {c11756};
    assign in13194_2 = {c11757};
    Full_Adder FA_13194(s13194, c13194, in13194_1, in13194_2, c11755);
    wire[0:0] s13195, in13195_1, in13195_2;
    wire c13195;
    assign in13195_1 = {s11759[0]};
    assign in13195_2 = {s11760[0]};
    Full_Adder FA_13195(s13195, c13195, in13195_1, in13195_2, c11758);
    wire[0:0] s13196, in13196_1, in13196_2;
    wire c13196;
    assign in13196_1 = {s11762[0]};
    assign in13196_2 = {s11763[0]};
    Full_Adder FA_13196(s13196, c13196, in13196_1, in13196_2, s11761[0]);
    wire[0:0] s13197, in13197_1, in13197_2;
    wire c13197;
    assign in13197_1 = {s11765[0]};
    assign in13197_2 = {s11766[0]};
    Full_Adder FA_13197(s13197, c13197, in13197_1, in13197_2, s11764[0]);
    wire[0:0] s13198, in13198_1, in13198_2;
    wire c13198;
    assign in13198_1 = {s9934[0]};
    assign in13198_2 = {c11759};
    Full_Adder FA_13198(s13198, c13198, in13198_1, in13198_2, s9933[0]);
    wire[0:0] s13199, in13199_1, in13199_2;
    wire c13199;
    assign in13199_1 = {c11761};
    assign in13199_2 = {c11762};
    Full_Adder FA_13199(s13199, c13199, in13199_1, in13199_2, c11760);
    wire[0:0] s13200, in13200_1, in13200_2;
    wire c13200;
    assign in13200_1 = {c11764};
    assign in13200_2 = {c11765};
    Full_Adder FA_13200(s13200, c13200, in13200_1, in13200_2, c11763);
    wire[0:0] s13201, in13201_1, in13201_2;
    wire c13201;
    assign in13201_1 = {s11767[0]};
    assign in13201_2 = {s11768[0]};
    Full_Adder FA_13201(s13201, c13201, in13201_1, in13201_2, c11766);
    wire[0:0] s13202, in13202_1, in13202_2;
    wire c13202;
    assign in13202_1 = {s11770[0]};
    assign in13202_2 = {s11771[0]};
    Full_Adder FA_13202(s13202, c13202, in13202_1, in13202_2, s11769[0]);
    wire[0:0] s13203, in13203_1, in13203_2;
    wire c13203;
    assign in13203_1 = {s11773[0]};
    assign in13203_2 = {s11774[0]};
    Full_Adder FA_13203(s13203, c13203, in13203_1, in13203_2, s11772[0]);
    wire[0:0] s13204, in13204_1, in13204_2;
    wire c13204;
    assign in13204_1 = {s9947[0]};
    assign in13204_2 = {c11767};
    Full_Adder FA_13204(s13204, c13204, in13204_1, in13204_2, s9946[0]);
    wire[0:0] s13205, in13205_1, in13205_2;
    wire c13205;
    assign in13205_1 = {c11769};
    assign in13205_2 = {c11770};
    Full_Adder FA_13205(s13205, c13205, in13205_1, in13205_2, c11768);
    wire[0:0] s13206, in13206_1, in13206_2;
    wire c13206;
    assign in13206_1 = {c11772};
    assign in13206_2 = {c11773};
    Full_Adder FA_13206(s13206, c13206, in13206_1, in13206_2, c11771);
    wire[0:0] s13207, in13207_1, in13207_2;
    wire c13207;
    assign in13207_1 = {s11775[0]};
    assign in13207_2 = {s11776[0]};
    Full_Adder FA_13207(s13207, c13207, in13207_1, in13207_2, c11774);
    wire[0:0] s13208, in13208_1, in13208_2;
    wire c13208;
    assign in13208_1 = {s11778[0]};
    assign in13208_2 = {s11779[0]};
    Full_Adder FA_13208(s13208, c13208, in13208_1, in13208_2, s11777[0]);
    wire[0:0] s13209, in13209_1, in13209_2;
    wire c13209;
    assign in13209_1 = {s11781[0]};
    assign in13209_2 = {s11782[0]};
    Full_Adder FA_13209(s13209, c13209, in13209_1, in13209_2, s11780[0]);
    wire[0:0] s13210, in13210_1, in13210_2;
    wire c13210;
    assign in13210_1 = {s9960[0]};
    assign in13210_2 = {c11775};
    Full_Adder FA_13210(s13210, c13210, in13210_1, in13210_2, s9959[0]);
    wire[0:0] s13211, in13211_1, in13211_2;
    wire c13211;
    assign in13211_1 = {c11777};
    assign in13211_2 = {c11778};
    Full_Adder FA_13211(s13211, c13211, in13211_1, in13211_2, c11776);
    wire[0:0] s13212, in13212_1, in13212_2;
    wire c13212;
    assign in13212_1 = {c11780};
    assign in13212_2 = {c11781};
    Full_Adder FA_13212(s13212, c13212, in13212_1, in13212_2, c11779);
    wire[0:0] s13213, in13213_1, in13213_2;
    wire c13213;
    assign in13213_1 = {s11783[0]};
    assign in13213_2 = {s11784[0]};
    Full_Adder FA_13213(s13213, c13213, in13213_1, in13213_2, c11782);
    wire[0:0] s13214, in13214_1, in13214_2;
    wire c13214;
    assign in13214_1 = {s11786[0]};
    assign in13214_2 = {s11787[0]};
    Full_Adder FA_13214(s13214, c13214, in13214_1, in13214_2, s11785[0]);
    wire[0:0] s13215, in13215_1, in13215_2;
    wire c13215;
    assign in13215_1 = {s11789[0]};
    assign in13215_2 = {s11790[0]};
    Full_Adder FA_13215(s13215, c13215, in13215_1, in13215_2, s11788[0]);
    wire[0:0] s13216, in13216_1, in13216_2;
    wire c13216;
    assign in13216_1 = {s9973[0]};
    assign in13216_2 = {c11783};
    Full_Adder FA_13216(s13216, c13216, in13216_1, in13216_2, s9972[0]);
    wire[0:0] s13217, in13217_1, in13217_2;
    wire c13217;
    assign in13217_1 = {c11785};
    assign in13217_2 = {c11786};
    Full_Adder FA_13217(s13217, c13217, in13217_1, in13217_2, c11784);
    wire[0:0] s13218, in13218_1, in13218_2;
    wire c13218;
    assign in13218_1 = {c11788};
    assign in13218_2 = {c11789};
    Full_Adder FA_13218(s13218, c13218, in13218_1, in13218_2, c11787);
    wire[0:0] s13219, in13219_1, in13219_2;
    wire c13219;
    assign in13219_1 = {s11791[0]};
    assign in13219_2 = {s11792[0]};
    Full_Adder FA_13219(s13219, c13219, in13219_1, in13219_2, c11790);
    wire[0:0] s13220, in13220_1, in13220_2;
    wire c13220;
    assign in13220_1 = {s11794[0]};
    assign in13220_2 = {s11795[0]};
    Full_Adder FA_13220(s13220, c13220, in13220_1, in13220_2, s11793[0]);
    wire[0:0] s13221, in13221_1, in13221_2;
    wire c13221;
    assign in13221_1 = {s11797[0]};
    assign in13221_2 = {s11798[0]};
    Full_Adder FA_13221(s13221, c13221, in13221_1, in13221_2, s11796[0]);
    wire[0:0] s13222, in13222_1, in13222_2;
    wire c13222;
    assign in13222_1 = {s9986[0]};
    assign in13222_2 = {c11791};
    Full_Adder FA_13222(s13222, c13222, in13222_1, in13222_2, s9985[0]);
    wire[0:0] s13223, in13223_1, in13223_2;
    wire c13223;
    assign in13223_1 = {c11793};
    assign in13223_2 = {c11794};
    Full_Adder FA_13223(s13223, c13223, in13223_1, in13223_2, c11792);
    wire[0:0] s13224, in13224_1, in13224_2;
    wire c13224;
    assign in13224_1 = {c11796};
    assign in13224_2 = {c11797};
    Full_Adder FA_13224(s13224, c13224, in13224_1, in13224_2, c11795);
    wire[0:0] s13225, in13225_1, in13225_2;
    wire c13225;
    assign in13225_1 = {s11799[0]};
    assign in13225_2 = {s11800[0]};
    Full_Adder FA_13225(s13225, c13225, in13225_1, in13225_2, c11798);
    wire[0:0] s13226, in13226_1, in13226_2;
    wire c13226;
    assign in13226_1 = {s11802[0]};
    assign in13226_2 = {s11803[0]};
    Full_Adder FA_13226(s13226, c13226, in13226_1, in13226_2, s11801[0]);
    wire[0:0] s13227, in13227_1, in13227_2;
    wire c13227;
    assign in13227_1 = {s11805[0]};
    assign in13227_2 = {s11806[0]};
    Full_Adder FA_13227(s13227, c13227, in13227_1, in13227_2, s11804[0]);
    wire[0:0] s13228, in13228_1, in13228_2;
    wire c13228;
    assign in13228_1 = {s9999[0]};
    assign in13228_2 = {c11799};
    Full_Adder FA_13228(s13228, c13228, in13228_1, in13228_2, s9998[0]);
    wire[0:0] s13229, in13229_1, in13229_2;
    wire c13229;
    assign in13229_1 = {c11801};
    assign in13229_2 = {c11802};
    Full_Adder FA_13229(s13229, c13229, in13229_1, in13229_2, c11800);
    wire[0:0] s13230, in13230_1, in13230_2;
    wire c13230;
    assign in13230_1 = {c11804};
    assign in13230_2 = {c11805};
    Full_Adder FA_13230(s13230, c13230, in13230_1, in13230_2, c11803);
    wire[0:0] s13231, in13231_1, in13231_2;
    wire c13231;
    assign in13231_1 = {s11807[0]};
    assign in13231_2 = {s11808[0]};
    Full_Adder FA_13231(s13231, c13231, in13231_1, in13231_2, c11806);
    wire[0:0] s13232, in13232_1, in13232_2;
    wire c13232;
    assign in13232_1 = {s11810[0]};
    assign in13232_2 = {s11811[0]};
    Full_Adder FA_13232(s13232, c13232, in13232_1, in13232_2, s11809[0]);
    wire[0:0] s13233, in13233_1, in13233_2;
    wire c13233;
    assign in13233_1 = {s11813[0]};
    assign in13233_2 = {s11814[0]};
    Full_Adder FA_13233(s13233, c13233, in13233_1, in13233_2, s11812[0]);
    wire[0:0] s13234, in13234_1, in13234_2;
    wire c13234;
    assign in13234_1 = {s10012[0]};
    assign in13234_2 = {c11807};
    Full_Adder FA_13234(s13234, c13234, in13234_1, in13234_2, s10011[0]);
    wire[0:0] s13235, in13235_1, in13235_2;
    wire c13235;
    assign in13235_1 = {c11809};
    assign in13235_2 = {c11810};
    Full_Adder FA_13235(s13235, c13235, in13235_1, in13235_2, c11808);
    wire[0:0] s13236, in13236_1, in13236_2;
    wire c13236;
    assign in13236_1 = {c11812};
    assign in13236_2 = {c11813};
    Full_Adder FA_13236(s13236, c13236, in13236_1, in13236_2, c11811);
    wire[0:0] s13237, in13237_1, in13237_2;
    wire c13237;
    assign in13237_1 = {s11815[0]};
    assign in13237_2 = {s11816[0]};
    Full_Adder FA_13237(s13237, c13237, in13237_1, in13237_2, c11814);
    wire[0:0] s13238, in13238_1, in13238_2;
    wire c13238;
    assign in13238_1 = {s11818[0]};
    assign in13238_2 = {s11819[0]};
    Full_Adder FA_13238(s13238, c13238, in13238_1, in13238_2, s11817[0]);
    wire[0:0] s13239, in13239_1, in13239_2;
    wire c13239;
    assign in13239_1 = {s11821[0]};
    assign in13239_2 = {s11822[0]};
    Full_Adder FA_13239(s13239, c13239, in13239_1, in13239_2, s11820[0]);
    wire[0:0] s13240, in13240_1, in13240_2;
    wire c13240;
    assign in13240_1 = {s10025[0]};
    assign in13240_2 = {c11815};
    Full_Adder FA_13240(s13240, c13240, in13240_1, in13240_2, s10024[0]);
    wire[0:0] s13241, in13241_1, in13241_2;
    wire c13241;
    assign in13241_1 = {c11817};
    assign in13241_2 = {c11818};
    Full_Adder FA_13241(s13241, c13241, in13241_1, in13241_2, c11816);
    wire[0:0] s13242, in13242_1, in13242_2;
    wire c13242;
    assign in13242_1 = {c11820};
    assign in13242_2 = {c11821};
    Full_Adder FA_13242(s13242, c13242, in13242_1, in13242_2, c11819);
    wire[0:0] s13243, in13243_1, in13243_2;
    wire c13243;
    assign in13243_1 = {s11823[0]};
    assign in13243_2 = {s11824[0]};
    Full_Adder FA_13243(s13243, c13243, in13243_1, in13243_2, c11822);
    wire[0:0] s13244, in13244_1, in13244_2;
    wire c13244;
    assign in13244_1 = {s11826[0]};
    assign in13244_2 = {s11827[0]};
    Full_Adder FA_13244(s13244, c13244, in13244_1, in13244_2, s11825[0]);
    wire[0:0] s13245, in13245_1, in13245_2;
    wire c13245;
    assign in13245_1 = {s11829[0]};
    assign in13245_2 = {s11830[0]};
    Full_Adder FA_13245(s13245, c13245, in13245_1, in13245_2, s11828[0]);
    wire[0:0] s13246, in13246_1, in13246_2;
    wire c13246;
    assign in13246_1 = {s10038[0]};
    assign in13246_2 = {c11823};
    Full_Adder FA_13246(s13246, c13246, in13246_1, in13246_2, s10037[0]);
    wire[0:0] s13247, in13247_1, in13247_2;
    wire c13247;
    assign in13247_1 = {c11825};
    assign in13247_2 = {c11826};
    Full_Adder FA_13247(s13247, c13247, in13247_1, in13247_2, c11824);
    wire[0:0] s13248, in13248_1, in13248_2;
    wire c13248;
    assign in13248_1 = {c11828};
    assign in13248_2 = {c11829};
    Full_Adder FA_13248(s13248, c13248, in13248_1, in13248_2, c11827);
    wire[0:0] s13249, in13249_1, in13249_2;
    wire c13249;
    assign in13249_1 = {s11831[0]};
    assign in13249_2 = {s11832[0]};
    Full_Adder FA_13249(s13249, c13249, in13249_1, in13249_2, c11830);
    wire[0:0] s13250, in13250_1, in13250_2;
    wire c13250;
    assign in13250_1 = {s11834[0]};
    assign in13250_2 = {s11835[0]};
    Full_Adder FA_13250(s13250, c13250, in13250_1, in13250_2, s11833[0]);
    wire[0:0] s13251, in13251_1, in13251_2;
    wire c13251;
    assign in13251_1 = {s11837[0]};
    assign in13251_2 = {s11838[0]};
    Full_Adder FA_13251(s13251, c13251, in13251_1, in13251_2, s11836[0]);
    wire[0:0] s13252, in13252_1, in13252_2;
    wire c13252;
    assign in13252_1 = {s10051[0]};
    assign in13252_2 = {c11831};
    Full_Adder FA_13252(s13252, c13252, in13252_1, in13252_2, s10050[0]);
    wire[0:0] s13253, in13253_1, in13253_2;
    wire c13253;
    assign in13253_1 = {c11833};
    assign in13253_2 = {c11834};
    Full_Adder FA_13253(s13253, c13253, in13253_1, in13253_2, c11832);
    wire[0:0] s13254, in13254_1, in13254_2;
    wire c13254;
    assign in13254_1 = {c11836};
    assign in13254_2 = {c11837};
    Full_Adder FA_13254(s13254, c13254, in13254_1, in13254_2, c11835);
    wire[0:0] s13255, in13255_1, in13255_2;
    wire c13255;
    assign in13255_1 = {s11839[0]};
    assign in13255_2 = {s11840[0]};
    Full_Adder FA_13255(s13255, c13255, in13255_1, in13255_2, c11838);
    wire[0:0] s13256, in13256_1, in13256_2;
    wire c13256;
    assign in13256_1 = {s11842[0]};
    assign in13256_2 = {s11843[0]};
    Full_Adder FA_13256(s13256, c13256, in13256_1, in13256_2, s11841[0]);
    wire[0:0] s13257, in13257_1, in13257_2;
    wire c13257;
    assign in13257_1 = {s11845[0]};
    assign in13257_2 = {s11846[0]};
    Full_Adder FA_13257(s13257, c13257, in13257_1, in13257_2, s11844[0]);
    wire[0:0] s13258, in13258_1, in13258_2;
    wire c13258;
    assign in13258_1 = {s10064[0]};
    assign in13258_2 = {c11839};
    Full_Adder FA_13258(s13258, c13258, in13258_1, in13258_2, s10063[0]);
    wire[0:0] s13259, in13259_1, in13259_2;
    wire c13259;
    assign in13259_1 = {c11841};
    assign in13259_2 = {c11842};
    Full_Adder FA_13259(s13259, c13259, in13259_1, in13259_2, c11840);
    wire[0:0] s13260, in13260_1, in13260_2;
    wire c13260;
    assign in13260_1 = {c11844};
    assign in13260_2 = {c11845};
    Full_Adder FA_13260(s13260, c13260, in13260_1, in13260_2, c11843);
    wire[0:0] s13261, in13261_1, in13261_2;
    wire c13261;
    assign in13261_1 = {s11847[0]};
    assign in13261_2 = {s11848[0]};
    Full_Adder FA_13261(s13261, c13261, in13261_1, in13261_2, c11846);
    wire[0:0] s13262, in13262_1, in13262_2;
    wire c13262;
    assign in13262_1 = {s11850[0]};
    assign in13262_2 = {s11851[0]};
    Full_Adder FA_13262(s13262, c13262, in13262_1, in13262_2, s11849[0]);
    wire[0:0] s13263, in13263_1, in13263_2;
    wire c13263;
    assign in13263_1 = {s11853[0]};
    assign in13263_2 = {s11854[0]};
    Full_Adder FA_13263(s13263, c13263, in13263_1, in13263_2, s11852[0]);
    wire[0:0] s13264, in13264_1, in13264_2;
    wire c13264;
    assign in13264_1 = {s10077[0]};
    assign in13264_2 = {c11847};
    Full_Adder FA_13264(s13264, c13264, in13264_1, in13264_2, s10076[0]);
    wire[0:0] s13265, in13265_1, in13265_2;
    wire c13265;
    assign in13265_1 = {c11849};
    assign in13265_2 = {c11850};
    Full_Adder FA_13265(s13265, c13265, in13265_1, in13265_2, c11848);
    wire[0:0] s13266, in13266_1, in13266_2;
    wire c13266;
    assign in13266_1 = {c11852};
    assign in13266_2 = {c11853};
    Full_Adder FA_13266(s13266, c13266, in13266_1, in13266_2, c11851);
    wire[0:0] s13267, in13267_1, in13267_2;
    wire c13267;
    assign in13267_1 = {s11855[0]};
    assign in13267_2 = {s11856[0]};
    Full_Adder FA_13267(s13267, c13267, in13267_1, in13267_2, c11854);
    wire[0:0] s13268, in13268_1, in13268_2;
    wire c13268;
    assign in13268_1 = {s11858[0]};
    assign in13268_2 = {s11859[0]};
    Full_Adder FA_13268(s13268, c13268, in13268_1, in13268_2, s11857[0]);
    wire[0:0] s13269, in13269_1, in13269_2;
    wire c13269;
    assign in13269_1 = {s11861[0]};
    assign in13269_2 = {s11862[0]};
    Full_Adder FA_13269(s13269, c13269, in13269_1, in13269_2, s11860[0]);
    wire[0:0] s13270, in13270_1, in13270_2;
    wire c13270;
    assign in13270_1 = {s10090[0]};
    assign in13270_2 = {c11855};
    Full_Adder FA_13270(s13270, c13270, in13270_1, in13270_2, s10089[0]);
    wire[0:0] s13271, in13271_1, in13271_2;
    wire c13271;
    assign in13271_1 = {c11857};
    assign in13271_2 = {c11858};
    Full_Adder FA_13271(s13271, c13271, in13271_1, in13271_2, c11856);
    wire[0:0] s13272, in13272_1, in13272_2;
    wire c13272;
    assign in13272_1 = {c11860};
    assign in13272_2 = {c11861};
    Full_Adder FA_13272(s13272, c13272, in13272_1, in13272_2, c11859);
    wire[0:0] s13273, in13273_1, in13273_2;
    wire c13273;
    assign in13273_1 = {s11863[0]};
    assign in13273_2 = {s11864[0]};
    Full_Adder FA_13273(s13273, c13273, in13273_1, in13273_2, c11862);
    wire[0:0] s13274, in13274_1, in13274_2;
    wire c13274;
    assign in13274_1 = {s11866[0]};
    assign in13274_2 = {s11867[0]};
    Full_Adder FA_13274(s13274, c13274, in13274_1, in13274_2, s11865[0]);
    wire[0:0] s13275, in13275_1, in13275_2;
    wire c13275;
    assign in13275_1 = {s11869[0]};
    assign in13275_2 = {s11870[0]};
    Full_Adder FA_13275(s13275, c13275, in13275_1, in13275_2, s11868[0]);
    wire[0:0] s13276, in13276_1, in13276_2;
    wire c13276;
    assign in13276_1 = {s10103[0]};
    assign in13276_2 = {c11863};
    Full_Adder FA_13276(s13276, c13276, in13276_1, in13276_2, s10102[0]);
    wire[0:0] s13277, in13277_1, in13277_2;
    wire c13277;
    assign in13277_1 = {c11865};
    assign in13277_2 = {c11866};
    Full_Adder FA_13277(s13277, c13277, in13277_1, in13277_2, c11864);
    wire[0:0] s13278, in13278_1, in13278_2;
    wire c13278;
    assign in13278_1 = {c11868};
    assign in13278_2 = {c11869};
    Full_Adder FA_13278(s13278, c13278, in13278_1, in13278_2, c11867);
    wire[0:0] s13279, in13279_1, in13279_2;
    wire c13279;
    assign in13279_1 = {s11871[0]};
    assign in13279_2 = {s11872[0]};
    Full_Adder FA_13279(s13279, c13279, in13279_1, in13279_2, c11870);
    wire[0:0] s13280, in13280_1, in13280_2;
    wire c13280;
    assign in13280_1 = {s11874[0]};
    assign in13280_2 = {s11875[0]};
    Full_Adder FA_13280(s13280, c13280, in13280_1, in13280_2, s11873[0]);
    wire[0:0] s13281, in13281_1, in13281_2;
    wire c13281;
    assign in13281_1 = {s11877[0]};
    assign in13281_2 = {s11878[0]};
    Full_Adder FA_13281(s13281, c13281, in13281_1, in13281_2, s11876[0]);
    wire[0:0] s13282, in13282_1, in13282_2;
    wire c13282;
    assign in13282_1 = {s10116[0]};
    assign in13282_2 = {c11871};
    Full_Adder FA_13282(s13282, c13282, in13282_1, in13282_2, s10115[0]);
    wire[0:0] s13283, in13283_1, in13283_2;
    wire c13283;
    assign in13283_1 = {c11873};
    assign in13283_2 = {c11874};
    Full_Adder FA_13283(s13283, c13283, in13283_1, in13283_2, c11872);
    wire[0:0] s13284, in13284_1, in13284_2;
    wire c13284;
    assign in13284_1 = {c11876};
    assign in13284_2 = {c11877};
    Full_Adder FA_13284(s13284, c13284, in13284_1, in13284_2, c11875);
    wire[0:0] s13285, in13285_1, in13285_2;
    wire c13285;
    assign in13285_1 = {s11879[0]};
    assign in13285_2 = {s11880[0]};
    Full_Adder FA_13285(s13285, c13285, in13285_1, in13285_2, c11878);
    wire[0:0] s13286, in13286_1, in13286_2;
    wire c13286;
    assign in13286_1 = {s11882[0]};
    assign in13286_2 = {s11883[0]};
    Full_Adder FA_13286(s13286, c13286, in13286_1, in13286_2, s11881[0]);
    wire[0:0] s13287, in13287_1, in13287_2;
    wire c13287;
    assign in13287_1 = {s11885[0]};
    assign in13287_2 = {s11886[0]};
    Full_Adder FA_13287(s13287, c13287, in13287_1, in13287_2, s11884[0]);
    wire[0:0] s13288, in13288_1, in13288_2;
    wire c13288;
    assign in13288_1 = {s10129[0]};
    assign in13288_2 = {c11879};
    Full_Adder FA_13288(s13288, c13288, in13288_1, in13288_2, s10128[0]);
    wire[0:0] s13289, in13289_1, in13289_2;
    wire c13289;
    assign in13289_1 = {c11881};
    assign in13289_2 = {c11882};
    Full_Adder FA_13289(s13289, c13289, in13289_1, in13289_2, c11880);
    wire[0:0] s13290, in13290_1, in13290_2;
    wire c13290;
    assign in13290_1 = {c11884};
    assign in13290_2 = {c11885};
    Full_Adder FA_13290(s13290, c13290, in13290_1, in13290_2, c11883);
    wire[0:0] s13291, in13291_1, in13291_2;
    wire c13291;
    assign in13291_1 = {s11887[0]};
    assign in13291_2 = {s11888[0]};
    Full_Adder FA_13291(s13291, c13291, in13291_1, in13291_2, c11886);
    wire[0:0] s13292, in13292_1, in13292_2;
    wire c13292;
    assign in13292_1 = {s11890[0]};
    assign in13292_2 = {s11891[0]};
    Full_Adder FA_13292(s13292, c13292, in13292_1, in13292_2, s11889[0]);
    wire[0:0] s13293, in13293_1, in13293_2;
    wire c13293;
    assign in13293_1 = {s11893[0]};
    assign in13293_2 = {s11894[0]};
    Full_Adder FA_13293(s13293, c13293, in13293_1, in13293_2, s11892[0]);
    wire[0:0] s13294, in13294_1, in13294_2;
    wire c13294;
    assign in13294_1 = {s10142[0]};
    assign in13294_2 = {c11887};
    Full_Adder FA_13294(s13294, c13294, in13294_1, in13294_2, s10141[0]);
    wire[0:0] s13295, in13295_1, in13295_2;
    wire c13295;
    assign in13295_1 = {c11889};
    assign in13295_2 = {c11890};
    Full_Adder FA_13295(s13295, c13295, in13295_1, in13295_2, c11888);
    wire[0:0] s13296, in13296_1, in13296_2;
    wire c13296;
    assign in13296_1 = {c11892};
    assign in13296_2 = {c11893};
    Full_Adder FA_13296(s13296, c13296, in13296_1, in13296_2, c11891);
    wire[0:0] s13297, in13297_1, in13297_2;
    wire c13297;
    assign in13297_1 = {s11895[0]};
    assign in13297_2 = {s11896[0]};
    Full_Adder FA_13297(s13297, c13297, in13297_1, in13297_2, c11894);
    wire[0:0] s13298, in13298_1, in13298_2;
    wire c13298;
    assign in13298_1 = {s11898[0]};
    assign in13298_2 = {s11899[0]};
    Full_Adder FA_13298(s13298, c13298, in13298_1, in13298_2, s11897[0]);
    wire[0:0] s13299, in13299_1, in13299_2;
    wire c13299;
    assign in13299_1 = {s11901[0]};
    assign in13299_2 = {s11902[0]};
    Full_Adder FA_13299(s13299, c13299, in13299_1, in13299_2, s11900[0]);
    wire[0:0] s13300, in13300_1, in13300_2;
    wire c13300;
    assign in13300_1 = {s10155[0]};
    assign in13300_2 = {c11895};
    Full_Adder FA_13300(s13300, c13300, in13300_1, in13300_2, s10154[0]);
    wire[0:0] s13301, in13301_1, in13301_2;
    wire c13301;
    assign in13301_1 = {c11897};
    assign in13301_2 = {c11898};
    Full_Adder FA_13301(s13301, c13301, in13301_1, in13301_2, c11896);
    wire[0:0] s13302, in13302_1, in13302_2;
    wire c13302;
    assign in13302_1 = {c11900};
    assign in13302_2 = {c11901};
    Full_Adder FA_13302(s13302, c13302, in13302_1, in13302_2, c11899);
    wire[0:0] s13303, in13303_1, in13303_2;
    wire c13303;
    assign in13303_1 = {s11903[0]};
    assign in13303_2 = {s11904[0]};
    Full_Adder FA_13303(s13303, c13303, in13303_1, in13303_2, c11902);
    wire[0:0] s13304, in13304_1, in13304_2;
    wire c13304;
    assign in13304_1 = {s11906[0]};
    assign in13304_2 = {s11907[0]};
    Full_Adder FA_13304(s13304, c13304, in13304_1, in13304_2, s11905[0]);
    wire[0:0] s13305, in13305_1, in13305_2;
    wire c13305;
    assign in13305_1 = {s11909[0]};
    assign in13305_2 = {s11910[0]};
    Full_Adder FA_13305(s13305, c13305, in13305_1, in13305_2, s11908[0]);
    wire[0:0] s13306, in13306_1, in13306_2;
    wire c13306;
    assign in13306_1 = {s10168[0]};
    assign in13306_2 = {c11903};
    Full_Adder FA_13306(s13306, c13306, in13306_1, in13306_2, s10167[0]);
    wire[0:0] s13307, in13307_1, in13307_2;
    wire c13307;
    assign in13307_1 = {c11905};
    assign in13307_2 = {c11906};
    Full_Adder FA_13307(s13307, c13307, in13307_1, in13307_2, c11904);
    wire[0:0] s13308, in13308_1, in13308_2;
    wire c13308;
    assign in13308_1 = {c11908};
    assign in13308_2 = {c11909};
    Full_Adder FA_13308(s13308, c13308, in13308_1, in13308_2, c11907);
    wire[0:0] s13309, in13309_1, in13309_2;
    wire c13309;
    assign in13309_1 = {s11911[0]};
    assign in13309_2 = {s11912[0]};
    Full_Adder FA_13309(s13309, c13309, in13309_1, in13309_2, c11910);
    wire[0:0] s13310, in13310_1, in13310_2;
    wire c13310;
    assign in13310_1 = {s11914[0]};
    assign in13310_2 = {s11915[0]};
    Full_Adder FA_13310(s13310, c13310, in13310_1, in13310_2, s11913[0]);
    wire[0:0] s13311, in13311_1, in13311_2;
    wire c13311;
    assign in13311_1 = {s11917[0]};
    assign in13311_2 = {s11918[0]};
    Full_Adder FA_13311(s13311, c13311, in13311_1, in13311_2, s11916[0]);
    wire[0:0] s13312, in13312_1, in13312_2;
    wire c13312;
    assign in13312_1 = {s10181[0]};
    assign in13312_2 = {c11911};
    Full_Adder FA_13312(s13312, c13312, in13312_1, in13312_2, s10180[0]);
    wire[0:0] s13313, in13313_1, in13313_2;
    wire c13313;
    assign in13313_1 = {c11913};
    assign in13313_2 = {c11914};
    Full_Adder FA_13313(s13313, c13313, in13313_1, in13313_2, c11912);
    wire[0:0] s13314, in13314_1, in13314_2;
    wire c13314;
    assign in13314_1 = {c11916};
    assign in13314_2 = {c11917};
    Full_Adder FA_13314(s13314, c13314, in13314_1, in13314_2, c11915);
    wire[0:0] s13315, in13315_1, in13315_2;
    wire c13315;
    assign in13315_1 = {s11919[0]};
    assign in13315_2 = {s11920[0]};
    Full_Adder FA_13315(s13315, c13315, in13315_1, in13315_2, c11918);
    wire[0:0] s13316, in13316_1, in13316_2;
    wire c13316;
    assign in13316_1 = {s11922[0]};
    assign in13316_2 = {s11923[0]};
    Full_Adder FA_13316(s13316, c13316, in13316_1, in13316_2, s11921[0]);
    wire[0:0] s13317, in13317_1, in13317_2;
    wire c13317;
    assign in13317_1 = {s11925[0]};
    assign in13317_2 = {s11926[0]};
    Full_Adder FA_13317(s13317, c13317, in13317_1, in13317_2, s11924[0]);
    wire[0:0] s13318, in13318_1, in13318_2;
    wire c13318;
    assign in13318_1 = {s10194[0]};
    assign in13318_2 = {c11919};
    Full_Adder FA_13318(s13318, c13318, in13318_1, in13318_2, s10193[0]);
    wire[0:0] s13319, in13319_1, in13319_2;
    wire c13319;
    assign in13319_1 = {c11921};
    assign in13319_2 = {c11922};
    Full_Adder FA_13319(s13319, c13319, in13319_1, in13319_2, c11920);
    wire[0:0] s13320, in13320_1, in13320_2;
    wire c13320;
    assign in13320_1 = {c11924};
    assign in13320_2 = {c11925};
    Full_Adder FA_13320(s13320, c13320, in13320_1, in13320_2, c11923);
    wire[0:0] s13321, in13321_1, in13321_2;
    wire c13321;
    assign in13321_1 = {s11927[0]};
    assign in13321_2 = {s11928[0]};
    Full_Adder FA_13321(s13321, c13321, in13321_1, in13321_2, c11926);
    wire[0:0] s13322, in13322_1, in13322_2;
    wire c13322;
    assign in13322_1 = {s11930[0]};
    assign in13322_2 = {s11931[0]};
    Full_Adder FA_13322(s13322, c13322, in13322_1, in13322_2, s11929[0]);
    wire[0:0] s13323, in13323_1, in13323_2;
    wire c13323;
    assign in13323_1 = {s11933[0]};
    assign in13323_2 = {s11934[0]};
    Full_Adder FA_13323(s13323, c13323, in13323_1, in13323_2, s11932[0]);
    wire[0:0] s13324, in13324_1, in13324_2;
    wire c13324;
    assign in13324_1 = {s10207[0]};
    assign in13324_2 = {c11927};
    Full_Adder FA_13324(s13324, c13324, in13324_1, in13324_2, s10206[0]);
    wire[0:0] s13325, in13325_1, in13325_2;
    wire c13325;
    assign in13325_1 = {c11929};
    assign in13325_2 = {c11930};
    Full_Adder FA_13325(s13325, c13325, in13325_1, in13325_2, c11928);
    wire[0:0] s13326, in13326_1, in13326_2;
    wire c13326;
    assign in13326_1 = {c11932};
    assign in13326_2 = {c11933};
    Full_Adder FA_13326(s13326, c13326, in13326_1, in13326_2, c11931);
    wire[0:0] s13327, in13327_1, in13327_2;
    wire c13327;
    assign in13327_1 = {s11935[0]};
    assign in13327_2 = {s11936[0]};
    Full_Adder FA_13327(s13327, c13327, in13327_1, in13327_2, c11934);
    wire[0:0] s13328, in13328_1, in13328_2;
    wire c13328;
    assign in13328_1 = {s11938[0]};
    assign in13328_2 = {s11939[0]};
    Full_Adder FA_13328(s13328, c13328, in13328_1, in13328_2, s11937[0]);
    wire[0:0] s13329, in13329_1, in13329_2;
    wire c13329;
    assign in13329_1 = {s11941[0]};
    assign in13329_2 = {s11942[0]};
    Full_Adder FA_13329(s13329, c13329, in13329_1, in13329_2, s11940[0]);
    wire[0:0] s13330, in13330_1, in13330_2;
    wire c13330;
    assign in13330_1 = {s10220[0]};
    assign in13330_2 = {c11935};
    Full_Adder FA_13330(s13330, c13330, in13330_1, in13330_2, s10219[0]);
    wire[0:0] s13331, in13331_1, in13331_2;
    wire c13331;
    assign in13331_1 = {c11937};
    assign in13331_2 = {c11938};
    Full_Adder FA_13331(s13331, c13331, in13331_1, in13331_2, c11936);
    wire[0:0] s13332, in13332_1, in13332_2;
    wire c13332;
    assign in13332_1 = {c11940};
    assign in13332_2 = {c11941};
    Full_Adder FA_13332(s13332, c13332, in13332_1, in13332_2, c11939);
    wire[0:0] s13333, in13333_1, in13333_2;
    wire c13333;
    assign in13333_1 = {s11943[0]};
    assign in13333_2 = {s11944[0]};
    Full_Adder FA_13333(s13333, c13333, in13333_1, in13333_2, c11942);
    wire[0:0] s13334, in13334_1, in13334_2;
    wire c13334;
    assign in13334_1 = {s11946[0]};
    assign in13334_2 = {s11947[0]};
    Full_Adder FA_13334(s13334, c13334, in13334_1, in13334_2, s11945[0]);
    wire[0:0] s13335, in13335_1, in13335_2;
    wire c13335;
    assign in13335_1 = {s11949[0]};
    assign in13335_2 = {s11950[0]};
    Full_Adder FA_13335(s13335, c13335, in13335_1, in13335_2, s11948[0]);
    wire[0:0] s13336, in13336_1, in13336_2;
    wire c13336;
    assign in13336_1 = {s10233[0]};
    assign in13336_2 = {c11943};
    Full_Adder FA_13336(s13336, c13336, in13336_1, in13336_2, s10232[0]);
    wire[0:0] s13337, in13337_1, in13337_2;
    wire c13337;
    assign in13337_1 = {c11945};
    assign in13337_2 = {c11946};
    Full_Adder FA_13337(s13337, c13337, in13337_1, in13337_2, c11944);
    wire[0:0] s13338, in13338_1, in13338_2;
    wire c13338;
    assign in13338_1 = {c11948};
    assign in13338_2 = {c11949};
    Full_Adder FA_13338(s13338, c13338, in13338_1, in13338_2, c11947);
    wire[0:0] s13339, in13339_1, in13339_2;
    wire c13339;
    assign in13339_1 = {s11951[0]};
    assign in13339_2 = {s11952[0]};
    Full_Adder FA_13339(s13339, c13339, in13339_1, in13339_2, c11950);
    wire[0:0] s13340, in13340_1, in13340_2;
    wire c13340;
    assign in13340_1 = {s11954[0]};
    assign in13340_2 = {s11955[0]};
    Full_Adder FA_13340(s13340, c13340, in13340_1, in13340_2, s11953[0]);
    wire[0:0] s13341, in13341_1, in13341_2;
    wire c13341;
    assign in13341_1 = {s11957[0]};
    assign in13341_2 = {s11958[0]};
    Full_Adder FA_13341(s13341, c13341, in13341_1, in13341_2, s11956[0]);
    wire[0:0] s13342, in13342_1, in13342_2;
    wire c13342;
    assign in13342_1 = {s10246[0]};
    assign in13342_2 = {c11951};
    Full_Adder FA_13342(s13342, c13342, in13342_1, in13342_2, s10245[0]);
    wire[0:0] s13343, in13343_1, in13343_2;
    wire c13343;
    assign in13343_1 = {c11953};
    assign in13343_2 = {c11954};
    Full_Adder FA_13343(s13343, c13343, in13343_1, in13343_2, c11952);
    wire[0:0] s13344, in13344_1, in13344_2;
    wire c13344;
    assign in13344_1 = {c11956};
    assign in13344_2 = {c11957};
    Full_Adder FA_13344(s13344, c13344, in13344_1, in13344_2, c11955);
    wire[0:0] s13345, in13345_1, in13345_2;
    wire c13345;
    assign in13345_1 = {s11959[0]};
    assign in13345_2 = {s11960[0]};
    Full_Adder FA_13345(s13345, c13345, in13345_1, in13345_2, c11958);
    wire[0:0] s13346, in13346_1, in13346_2;
    wire c13346;
    assign in13346_1 = {s11962[0]};
    assign in13346_2 = {s11963[0]};
    Full_Adder FA_13346(s13346, c13346, in13346_1, in13346_2, s11961[0]);
    wire[0:0] s13347, in13347_1, in13347_2;
    wire c13347;
    assign in13347_1 = {s11965[0]};
    assign in13347_2 = {s11966[0]};
    Full_Adder FA_13347(s13347, c13347, in13347_1, in13347_2, s11964[0]);
    wire[0:0] s13348, in13348_1, in13348_2;
    wire c13348;
    assign in13348_1 = {s10259[0]};
    assign in13348_2 = {c11959};
    Full_Adder FA_13348(s13348, c13348, in13348_1, in13348_2, s10258[0]);
    wire[0:0] s13349, in13349_1, in13349_2;
    wire c13349;
    assign in13349_1 = {c11961};
    assign in13349_2 = {c11962};
    Full_Adder FA_13349(s13349, c13349, in13349_1, in13349_2, c11960);
    wire[0:0] s13350, in13350_1, in13350_2;
    wire c13350;
    assign in13350_1 = {c11964};
    assign in13350_2 = {c11965};
    Full_Adder FA_13350(s13350, c13350, in13350_1, in13350_2, c11963);
    wire[0:0] s13351, in13351_1, in13351_2;
    wire c13351;
    assign in13351_1 = {s11967[0]};
    assign in13351_2 = {s11968[0]};
    Full_Adder FA_13351(s13351, c13351, in13351_1, in13351_2, c11966);
    wire[0:0] s13352, in13352_1, in13352_2;
    wire c13352;
    assign in13352_1 = {s11970[0]};
    assign in13352_2 = {s11971[0]};
    Full_Adder FA_13352(s13352, c13352, in13352_1, in13352_2, s11969[0]);
    wire[0:0] s13353, in13353_1, in13353_2;
    wire c13353;
    assign in13353_1 = {s11973[0]};
    assign in13353_2 = {s11974[0]};
    Full_Adder FA_13353(s13353, c13353, in13353_1, in13353_2, s11972[0]);
    wire[0:0] s13354, in13354_1, in13354_2;
    wire c13354;
    assign in13354_1 = {s10272[0]};
    assign in13354_2 = {c11967};
    Full_Adder FA_13354(s13354, c13354, in13354_1, in13354_2, s10271[0]);
    wire[0:0] s13355, in13355_1, in13355_2;
    wire c13355;
    assign in13355_1 = {c11969};
    assign in13355_2 = {c11970};
    Full_Adder FA_13355(s13355, c13355, in13355_1, in13355_2, c11968);
    wire[0:0] s13356, in13356_1, in13356_2;
    wire c13356;
    assign in13356_1 = {c11972};
    assign in13356_2 = {c11973};
    Full_Adder FA_13356(s13356, c13356, in13356_1, in13356_2, c11971);
    wire[0:0] s13357, in13357_1, in13357_2;
    wire c13357;
    assign in13357_1 = {s11975[0]};
    assign in13357_2 = {s11976[0]};
    Full_Adder FA_13357(s13357, c13357, in13357_1, in13357_2, c11974);
    wire[0:0] s13358, in13358_1, in13358_2;
    wire c13358;
    assign in13358_1 = {s11978[0]};
    assign in13358_2 = {s11979[0]};
    Full_Adder FA_13358(s13358, c13358, in13358_1, in13358_2, s11977[0]);
    wire[0:0] s13359, in13359_1, in13359_2;
    wire c13359;
    assign in13359_1 = {s11981[0]};
    assign in13359_2 = {s11982[0]};
    Full_Adder FA_13359(s13359, c13359, in13359_1, in13359_2, s11980[0]);
    wire[0:0] s13360, in13360_1, in13360_2;
    wire c13360;
    assign in13360_1 = {s10285[0]};
    assign in13360_2 = {c11975};
    Full_Adder FA_13360(s13360, c13360, in13360_1, in13360_2, s10284[0]);
    wire[0:0] s13361, in13361_1, in13361_2;
    wire c13361;
    assign in13361_1 = {c11977};
    assign in13361_2 = {c11978};
    Full_Adder FA_13361(s13361, c13361, in13361_1, in13361_2, c11976);
    wire[0:0] s13362, in13362_1, in13362_2;
    wire c13362;
    assign in13362_1 = {c11980};
    assign in13362_2 = {c11981};
    Full_Adder FA_13362(s13362, c13362, in13362_1, in13362_2, c11979);
    wire[0:0] s13363, in13363_1, in13363_2;
    wire c13363;
    assign in13363_1 = {s11983[0]};
    assign in13363_2 = {s11984[0]};
    Full_Adder FA_13363(s13363, c13363, in13363_1, in13363_2, c11982);
    wire[0:0] s13364, in13364_1, in13364_2;
    wire c13364;
    assign in13364_1 = {s11986[0]};
    assign in13364_2 = {s11987[0]};
    Full_Adder FA_13364(s13364, c13364, in13364_1, in13364_2, s11985[0]);
    wire[0:0] s13365, in13365_1, in13365_2;
    wire c13365;
    assign in13365_1 = {s11989[0]};
    assign in13365_2 = {s11990[0]};
    Full_Adder FA_13365(s13365, c13365, in13365_1, in13365_2, s11988[0]);
    wire[0:0] s13366, in13366_1, in13366_2;
    wire c13366;
    assign in13366_1 = {s10298[0]};
    assign in13366_2 = {c11983};
    Full_Adder FA_13366(s13366, c13366, in13366_1, in13366_2, s10297[0]);
    wire[0:0] s13367, in13367_1, in13367_2;
    wire c13367;
    assign in13367_1 = {c11985};
    assign in13367_2 = {c11986};
    Full_Adder FA_13367(s13367, c13367, in13367_1, in13367_2, c11984);
    wire[0:0] s13368, in13368_1, in13368_2;
    wire c13368;
    assign in13368_1 = {c11988};
    assign in13368_2 = {c11989};
    Full_Adder FA_13368(s13368, c13368, in13368_1, in13368_2, c11987);
    wire[0:0] s13369, in13369_1, in13369_2;
    wire c13369;
    assign in13369_1 = {s11991[0]};
    assign in13369_2 = {s11992[0]};
    Full_Adder FA_13369(s13369, c13369, in13369_1, in13369_2, c11990);
    wire[0:0] s13370, in13370_1, in13370_2;
    wire c13370;
    assign in13370_1 = {s11994[0]};
    assign in13370_2 = {s11995[0]};
    Full_Adder FA_13370(s13370, c13370, in13370_1, in13370_2, s11993[0]);
    wire[0:0] s13371, in13371_1, in13371_2;
    wire c13371;
    assign in13371_1 = {s11997[0]};
    assign in13371_2 = {s11998[0]};
    Full_Adder FA_13371(s13371, c13371, in13371_1, in13371_2, s11996[0]);
    wire[0:0] s13372, in13372_1, in13372_2;
    wire c13372;
    assign in13372_1 = {s10311[0]};
    assign in13372_2 = {c11991};
    Full_Adder FA_13372(s13372, c13372, in13372_1, in13372_2, s10310[0]);
    wire[0:0] s13373, in13373_1, in13373_2;
    wire c13373;
    assign in13373_1 = {c11993};
    assign in13373_2 = {c11994};
    Full_Adder FA_13373(s13373, c13373, in13373_1, in13373_2, c11992);
    wire[0:0] s13374, in13374_1, in13374_2;
    wire c13374;
    assign in13374_1 = {c11996};
    assign in13374_2 = {c11997};
    Full_Adder FA_13374(s13374, c13374, in13374_1, in13374_2, c11995);
    wire[0:0] s13375, in13375_1, in13375_2;
    wire c13375;
    assign in13375_1 = {s11999[0]};
    assign in13375_2 = {s12000[0]};
    Full_Adder FA_13375(s13375, c13375, in13375_1, in13375_2, c11998);
    wire[0:0] s13376, in13376_1, in13376_2;
    wire c13376;
    assign in13376_1 = {s12002[0]};
    assign in13376_2 = {s12003[0]};
    Full_Adder FA_13376(s13376, c13376, in13376_1, in13376_2, s12001[0]);
    wire[0:0] s13377, in13377_1, in13377_2;
    wire c13377;
    assign in13377_1 = {s12005[0]};
    assign in13377_2 = {s12006[0]};
    Full_Adder FA_13377(s13377, c13377, in13377_1, in13377_2, s12004[0]);
    wire[0:0] s13378, in13378_1, in13378_2;
    wire c13378;
    assign in13378_1 = {s10324[0]};
    assign in13378_2 = {c11999};
    Full_Adder FA_13378(s13378, c13378, in13378_1, in13378_2, s10323[0]);
    wire[0:0] s13379, in13379_1, in13379_2;
    wire c13379;
    assign in13379_1 = {c12001};
    assign in13379_2 = {c12002};
    Full_Adder FA_13379(s13379, c13379, in13379_1, in13379_2, c12000);
    wire[0:0] s13380, in13380_1, in13380_2;
    wire c13380;
    assign in13380_1 = {c12004};
    assign in13380_2 = {c12005};
    Full_Adder FA_13380(s13380, c13380, in13380_1, in13380_2, c12003);
    wire[0:0] s13381, in13381_1, in13381_2;
    wire c13381;
    assign in13381_1 = {s12007[0]};
    assign in13381_2 = {s12008[0]};
    Full_Adder FA_13381(s13381, c13381, in13381_1, in13381_2, c12006);
    wire[0:0] s13382, in13382_1, in13382_2;
    wire c13382;
    assign in13382_1 = {s12010[0]};
    assign in13382_2 = {s12011[0]};
    Full_Adder FA_13382(s13382, c13382, in13382_1, in13382_2, s12009[0]);
    wire[0:0] s13383, in13383_1, in13383_2;
    wire c13383;
    assign in13383_1 = {s12013[0]};
    assign in13383_2 = {s12014[0]};
    Full_Adder FA_13383(s13383, c13383, in13383_1, in13383_2, s12012[0]);
    wire[0:0] s13384, in13384_1, in13384_2;
    wire c13384;
    assign in13384_1 = {s10337[0]};
    assign in13384_2 = {c12007};
    Full_Adder FA_13384(s13384, c13384, in13384_1, in13384_2, s10336[0]);
    wire[0:0] s13385, in13385_1, in13385_2;
    wire c13385;
    assign in13385_1 = {c12009};
    assign in13385_2 = {c12010};
    Full_Adder FA_13385(s13385, c13385, in13385_1, in13385_2, c12008);
    wire[0:0] s13386, in13386_1, in13386_2;
    wire c13386;
    assign in13386_1 = {c12012};
    assign in13386_2 = {c12013};
    Full_Adder FA_13386(s13386, c13386, in13386_1, in13386_2, c12011);
    wire[0:0] s13387, in13387_1, in13387_2;
    wire c13387;
    assign in13387_1 = {s12015[0]};
    assign in13387_2 = {s12016[0]};
    Full_Adder FA_13387(s13387, c13387, in13387_1, in13387_2, c12014);
    wire[0:0] s13388, in13388_1, in13388_2;
    wire c13388;
    assign in13388_1 = {s12018[0]};
    assign in13388_2 = {s12019[0]};
    Full_Adder FA_13388(s13388, c13388, in13388_1, in13388_2, s12017[0]);
    wire[0:0] s13389, in13389_1, in13389_2;
    wire c13389;
    assign in13389_1 = {s12021[0]};
    assign in13389_2 = {s12022[0]};
    Full_Adder FA_13389(s13389, c13389, in13389_1, in13389_2, s12020[0]);
    wire[0:0] s13390, in13390_1, in13390_2;
    wire c13390;
    assign in13390_1 = {s10350[0]};
    assign in13390_2 = {c12015};
    Full_Adder FA_13390(s13390, c13390, in13390_1, in13390_2, s10349[0]);
    wire[0:0] s13391, in13391_1, in13391_2;
    wire c13391;
    assign in13391_1 = {c12017};
    assign in13391_2 = {c12018};
    Full_Adder FA_13391(s13391, c13391, in13391_1, in13391_2, c12016);
    wire[0:0] s13392, in13392_1, in13392_2;
    wire c13392;
    assign in13392_1 = {c12020};
    assign in13392_2 = {c12021};
    Full_Adder FA_13392(s13392, c13392, in13392_1, in13392_2, c12019);
    wire[0:0] s13393, in13393_1, in13393_2;
    wire c13393;
    assign in13393_1 = {s12023[0]};
    assign in13393_2 = {s12024[0]};
    Full_Adder FA_13393(s13393, c13393, in13393_1, in13393_2, c12022);
    wire[0:0] s13394, in13394_1, in13394_2;
    wire c13394;
    assign in13394_1 = {s12026[0]};
    assign in13394_2 = {s12027[0]};
    Full_Adder FA_13394(s13394, c13394, in13394_1, in13394_2, s12025[0]);
    wire[0:0] s13395, in13395_1, in13395_2;
    wire c13395;
    assign in13395_1 = {s12029[0]};
    assign in13395_2 = {s12030[0]};
    Full_Adder FA_13395(s13395, c13395, in13395_1, in13395_2, s12028[0]);
    wire[0:0] s13396, in13396_1, in13396_2;
    wire c13396;
    assign in13396_1 = {s10363[0]};
    assign in13396_2 = {c12023};
    Full_Adder FA_13396(s13396, c13396, in13396_1, in13396_2, s10362[0]);
    wire[0:0] s13397, in13397_1, in13397_2;
    wire c13397;
    assign in13397_1 = {c12025};
    assign in13397_2 = {c12026};
    Full_Adder FA_13397(s13397, c13397, in13397_1, in13397_2, c12024);
    wire[0:0] s13398, in13398_1, in13398_2;
    wire c13398;
    assign in13398_1 = {c12028};
    assign in13398_2 = {c12029};
    Full_Adder FA_13398(s13398, c13398, in13398_1, in13398_2, c12027);
    wire[0:0] s13399, in13399_1, in13399_2;
    wire c13399;
    assign in13399_1 = {s12031[0]};
    assign in13399_2 = {s12032[0]};
    Full_Adder FA_13399(s13399, c13399, in13399_1, in13399_2, c12030);
    wire[0:0] s13400, in13400_1, in13400_2;
    wire c13400;
    assign in13400_1 = {s12034[0]};
    assign in13400_2 = {s12035[0]};
    Full_Adder FA_13400(s13400, c13400, in13400_1, in13400_2, s12033[0]);
    wire[0:0] s13401, in13401_1, in13401_2;
    wire c13401;
    assign in13401_1 = {s12037[0]};
    assign in13401_2 = {s12038[0]};
    Full_Adder FA_13401(s13401, c13401, in13401_1, in13401_2, s12036[0]);
    wire[0:0] s13402, in13402_1, in13402_2;
    wire c13402;
    assign in13402_1 = {s10376[0]};
    assign in13402_2 = {c12031};
    Full_Adder FA_13402(s13402, c13402, in13402_1, in13402_2, s10375[0]);
    wire[0:0] s13403, in13403_1, in13403_2;
    wire c13403;
    assign in13403_1 = {c12033};
    assign in13403_2 = {c12034};
    Full_Adder FA_13403(s13403, c13403, in13403_1, in13403_2, c12032);
    wire[0:0] s13404, in13404_1, in13404_2;
    wire c13404;
    assign in13404_1 = {c12036};
    assign in13404_2 = {c12037};
    Full_Adder FA_13404(s13404, c13404, in13404_1, in13404_2, c12035);
    wire[0:0] s13405, in13405_1, in13405_2;
    wire c13405;
    assign in13405_1 = {s12039[0]};
    assign in13405_2 = {s12040[0]};
    Full_Adder FA_13405(s13405, c13405, in13405_1, in13405_2, c12038);
    wire[0:0] s13406, in13406_1, in13406_2;
    wire c13406;
    assign in13406_1 = {s12042[0]};
    assign in13406_2 = {s12043[0]};
    Full_Adder FA_13406(s13406, c13406, in13406_1, in13406_2, s12041[0]);
    wire[0:0] s13407, in13407_1, in13407_2;
    wire c13407;
    assign in13407_1 = {s12045[0]};
    assign in13407_2 = {s12046[0]};
    Full_Adder FA_13407(s13407, c13407, in13407_1, in13407_2, s12044[0]);
    wire[0:0] s13408, in13408_1, in13408_2;
    wire c13408;
    assign in13408_1 = {s10389[0]};
    assign in13408_2 = {c12039};
    Full_Adder FA_13408(s13408, c13408, in13408_1, in13408_2, s10388[0]);
    wire[0:0] s13409, in13409_1, in13409_2;
    wire c13409;
    assign in13409_1 = {c12041};
    assign in13409_2 = {c12042};
    Full_Adder FA_13409(s13409, c13409, in13409_1, in13409_2, c12040);
    wire[0:0] s13410, in13410_1, in13410_2;
    wire c13410;
    assign in13410_1 = {c12044};
    assign in13410_2 = {c12045};
    Full_Adder FA_13410(s13410, c13410, in13410_1, in13410_2, c12043);
    wire[0:0] s13411, in13411_1, in13411_2;
    wire c13411;
    assign in13411_1 = {s12047[0]};
    assign in13411_2 = {s12048[0]};
    Full_Adder FA_13411(s13411, c13411, in13411_1, in13411_2, c12046);
    wire[0:0] s13412, in13412_1, in13412_2;
    wire c13412;
    assign in13412_1 = {s12050[0]};
    assign in13412_2 = {s12051[0]};
    Full_Adder FA_13412(s13412, c13412, in13412_1, in13412_2, s12049[0]);
    wire[0:0] s13413, in13413_1, in13413_2;
    wire c13413;
    assign in13413_1 = {s12053[0]};
    assign in13413_2 = {s12054[0]};
    Full_Adder FA_13413(s13413, c13413, in13413_1, in13413_2, s12052[0]);
    wire[0:0] s13414, in13414_1, in13414_2;
    wire c13414;
    assign in13414_1 = {s10402[0]};
    assign in13414_2 = {c12047};
    Full_Adder FA_13414(s13414, c13414, in13414_1, in13414_2, s10401[0]);
    wire[0:0] s13415, in13415_1, in13415_2;
    wire c13415;
    assign in13415_1 = {c12049};
    assign in13415_2 = {c12050};
    Full_Adder FA_13415(s13415, c13415, in13415_1, in13415_2, c12048);
    wire[0:0] s13416, in13416_1, in13416_2;
    wire c13416;
    assign in13416_1 = {c12052};
    assign in13416_2 = {c12053};
    Full_Adder FA_13416(s13416, c13416, in13416_1, in13416_2, c12051);
    wire[0:0] s13417, in13417_1, in13417_2;
    wire c13417;
    assign in13417_1 = {s12055[0]};
    assign in13417_2 = {s12056[0]};
    Full_Adder FA_13417(s13417, c13417, in13417_1, in13417_2, c12054);
    wire[0:0] s13418, in13418_1, in13418_2;
    wire c13418;
    assign in13418_1 = {s12058[0]};
    assign in13418_2 = {s12059[0]};
    Full_Adder FA_13418(s13418, c13418, in13418_1, in13418_2, s12057[0]);
    wire[0:0] s13419, in13419_1, in13419_2;
    wire c13419;
    assign in13419_1 = {s12061[0]};
    assign in13419_2 = {s12062[0]};
    Full_Adder FA_13419(s13419, c13419, in13419_1, in13419_2, s12060[0]);
    wire[0:0] s13420, in13420_1, in13420_2;
    wire c13420;
    assign in13420_1 = {s10415[0]};
    assign in13420_2 = {c12055};
    Full_Adder FA_13420(s13420, c13420, in13420_1, in13420_2, s10414[0]);
    wire[0:0] s13421, in13421_1, in13421_2;
    wire c13421;
    assign in13421_1 = {c12057};
    assign in13421_2 = {c12058};
    Full_Adder FA_13421(s13421, c13421, in13421_1, in13421_2, c12056);
    wire[0:0] s13422, in13422_1, in13422_2;
    wire c13422;
    assign in13422_1 = {c12060};
    assign in13422_2 = {c12061};
    Full_Adder FA_13422(s13422, c13422, in13422_1, in13422_2, c12059);
    wire[0:0] s13423, in13423_1, in13423_2;
    wire c13423;
    assign in13423_1 = {s12063[0]};
    assign in13423_2 = {s12064[0]};
    Full_Adder FA_13423(s13423, c13423, in13423_1, in13423_2, c12062);
    wire[0:0] s13424, in13424_1, in13424_2;
    wire c13424;
    assign in13424_1 = {s12066[0]};
    assign in13424_2 = {s12067[0]};
    Full_Adder FA_13424(s13424, c13424, in13424_1, in13424_2, s12065[0]);
    wire[0:0] s13425, in13425_1, in13425_2;
    wire c13425;
    assign in13425_1 = {s12069[0]};
    assign in13425_2 = {s12070[0]};
    Full_Adder FA_13425(s13425, c13425, in13425_1, in13425_2, s12068[0]);
    wire[0:0] s13426, in13426_1, in13426_2;
    wire c13426;
    assign in13426_1 = {s10428[0]};
    assign in13426_2 = {c12063};
    Full_Adder FA_13426(s13426, c13426, in13426_1, in13426_2, s10427[0]);
    wire[0:0] s13427, in13427_1, in13427_2;
    wire c13427;
    assign in13427_1 = {c12065};
    assign in13427_2 = {c12066};
    Full_Adder FA_13427(s13427, c13427, in13427_1, in13427_2, c12064);
    wire[0:0] s13428, in13428_1, in13428_2;
    wire c13428;
    assign in13428_1 = {c12068};
    assign in13428_2 = {c12069};
    Full_Adder FA_13428(s13428, c13428, in13428_1, in13428_2, c12067);
    wire[0:0] s13429, in13429_1, in13429_2;
    wire c13429;
    assign in13429_1 = {s12071[0]};
    assign in13429_2 = {s12072[0]};
    Full_Adder FA_13429(s13429, c13429, in13429_1, in13429_2, c12070);
    wire[0:0] s13430, in13430_1, in13430_2;
    wire c13430;
    assign in13430_1 = {s12074[0]};
    assign in13430_2 = {s12075[0]};
    Full_Adder FA_13430(s13430, c13430, in13430_1, in13430_2, s12073[0]);
    wire[0:0] s13431, in13431_1, in13431_2;
    wire c13431;
    assign in13431_1 = {s12077[0]};
    assign in13431_2 = {s12078[0]};
    Full_Adder FA_13431(s13431, c13431, in13431_1, in13431_2, s12076[0]);
    wire[0:0] s13432, in13432_1, in13432_2;
    wire c13432;
    assign in13432_1 = {s10440[0]};
    assign in13432_2 = {c12071};
    Full_Adder FA_13432(s13432, c13432, in13432_1, in13432_2, s10439[0]);
    wire[0:0] s13433, in13433_1, in13433_2;
    wire c13433;
    assign in13433_1 = {c12073};
    assign in13433_2 = {c12074};
    Full_Adder FA_13433(s13433, c13433, in13433_1, in13433_2, c12072);
    wire[0:0] s13434, in13434_1, in13434_2;
    wire c13434;
    assign in13434_1 = {c12076};
    assign in13434_2 = {c12077};
    Full_Adder FA_13434(s13434, c13434, in13434_1, in13434_2, c12075);
    wire[0:0] s13435, in13435_1, in13435_2;
    wire c13435;
    assign in13435_1 = {s12079[0]};
    assign in13435_2 = {s12080[0]};
    Full_Adder FA_13435(s13435, c13435, in13435_1, in13435_2, c12078);
    wire[0:0] s13436, in13436_1, in13436_2;
    wire c13436;
    assign in13436_1 = {s12082[0]};
    assign in13436_2 = {s12083[0]};
    Full_Adder FA_13436(s13436, c13436, in13436_1, in13436_2, s12081[0]);
    wire[0:0] s13437, in13437_1, in13437_2;
    wire c13437;
    assign in13437_1 = {s12085[0]};
    assign in13437_2 = {s12086[0]};
    Full_Adder FA_13437(s13437, c13437, in13437_1, in13437_2, s12084[0]);
    wire[0:0] s13438, in13438_1, in13438_2;
    wire c13438;
    assign in13438_1 = {s10451[0]};
    assign in13438_2 = {c12079};
    Full_Adder FA_13438(s13438, c13438, in13438_1, in13438_2, s10450[0]);
    wire[0:0] s13439, in13439_1, in13439_2;
    wire c13439;
    assign in13439_1 = {c12081};
    assign in13439_2 = {c12082};
    Full_Adder FA_13439(s13439, c13439, in13439_1, in13439_2, c12080);
    wire[0:0] s13440, in13440_1, in13440_2;
    wire c13440;
    assign in13440_1 = {c12084};
    assign in13440_2 = {c12085};
    Full_Adder FA_13440(s13440, c13440, in13440_1, in13440_2, c12083);
    wire[0:0] s13441, in13441_1, in13441_2;
    wire c13441;
    assign in13441_1 = {s12087[0]};
    assign in13441_2 = {s12088[0]};
    Full_Adder FA_13441(s13441, c13441, in13441_1, in13441_2, c12086);
    wire[0:0] s13442, in13442_1, in13442_2;
    wire c13442;
    assign in13442_1 = {s12090[0]};
    assign in13442_2 = {s12091[0]};
    Full_Adder FA_13442(s13442, c13442, in13442_1, in13442_2, s12089[0]);
    wire[0:0] s13443, in13443_1, in13443_2;
    wire c13443;
    assign in13443_1 = {s12093[0]};
    assign in13443_2 = {s12094[0]};
    Full_Adder FA_13443(s13443, c13443, in13443_1, in13443_2, s12092[0]);
    wire[0:0] s13444, in13444_1, in13444_2;
    wire c13444;
    assign in13444_1 = {s10461[0]};
    assign in13444_2 = {c12087};
    Full_Adder FA_13444(s13444, c13444, in13444_1, in13444_2, s10460[0]);
    wire[0:0] s13445, in13445_1, in13445_2;
    wire c13445;
    assign in13445_1 = {c12089};
    assign in13445_2 = {c12090};
    Full_Adder FA_13445(s13445, c13445, in13445_1, in13445_2, c12088);
    wire[0:0] s13446, in13446_1, in13446_2;
    wire c13446;
    assign in13446_1 = {c12092};
    assign in13446_2 = {c12093};
    Full_Adder FA_13446(s13446, c13446, in13446_1, in13446_2, c12091);
    wire[0:0] s13447, in13447_1, in13447_2;
    wire c13447;
    assign in13447_1 = {s12095[0]};
    assign in13447_2 = {s12096[0]};
    Full_Adder FA_13447(s13447, c13447, in13447_1, in13447_2, c12094);
    wire[0:0] s13448, in13448_1, in13448_2;
    wire c13448;
    assign in13448_1 = {s12098[0]};
    assign in13448_2 = {s12099[0]};
    Full_Adder FA_13448(s13448, c13448, in13448_1, in13448_2, s12097[0]);
    wire[0:0] s13449, in13449_1, in13449_2;
    wire c13449;
    assign in13449_1 = {s12101[0]};
    assign in13449_2 = {s12102[0]};
    Full_Adder FA_13449(s13449, c13449, in13449_1, in13449_2, s12100[0]);
    wire[0:0] s13450, in13450_1, in13450_2;
    wire c13450;
    assign in13450_1 = {s10470[0]};
    assign in13450_2 = {c12095};
    Full_Adder FA_13450(s13450, c13450, in13450_1, in13450_2, s10469[0]);
    wire[0:0] s13451, in13451_1, in13451_2;
    wire c13451;
    assign in13451_1 = {c12097};
    assign in13451_2 = {c12098};
    Full_Adder FA_13451(s13451, c13451, in13451_1, in13451_2, c12096);
    wire[0:0] s13452, in13452_1, in13452_2;
    wire c13452;
    assign in13452_1 = {c12100};
    assign in13452_2 = {c12101};
    Full_Adder FA_13452(s13452, c13452, in13452_1, in13452_2, c12099);
    wire[0:0] s13453, in13453_1, in13453_2;
    wire c13453;
    assign in13453_1 = {s12103[0]};
    assign in13453_2 = {s12104[0]};
    Full_Adder FA_13453(s13453, c13453, in13453_1, in13453_2, c12102);
    wire[0:0] s13454, in13454_1, in13454_2;
    wire c13454;
    assign in13454_1 = {s12106[0]};
    assign in13454_2 = {s12107[0]};
    Full_Adder FA_13454(s13454, c13454, in13454_1, in13454_2, s12105[0]);
    wire[0:0] s13455, in13455_1, in13455_2;
    wire c13455;
    assign in13455_1 = {s12109[0]};
    assign in13455_2 = {s12110[0]};
    Full_Adder FA_13455(s13455, c13455, in13455_1, in13455_2, s12108[0]);
    wire[0:0] s13456, in13456_1, in13456_2;
    wire c13456;
    assign in13456_1 = {s10478[0]};
    assign in13456_2 = {c12103};
    Full_Adder FA_13456(s13456, c13456, in13456_1, in13456_2, s10477[0]);
    wire[0:0] s13457, in13457_1, in13457_2;
    wire c13457;
    assign in13457_1 = {c12105};
    assign in13457_2 = {c12106};
    Full_Adder FA_13457(s13457, c13457, in13457_1, in13457_2, c12104);
    wire[0:0] s13458, in13458_1, in13458_2;
    wire c13458;
    assign in13458_1 = {c12108};
    assign in13458_2 = {c12109};
    Full_Adder FA_13458(s13458, c13458, in13458_1, in13458_2, c12107);
    wire[0:0] s13459, in13459_1, in13459_2;
    wire c13459;
    assign in13459_1 = {s12111[0]};
    assign in13459_2 = {s12112[0]};
    Full_Adder FA_13459(s13459, c13459, in13459_1, in13459_2, c12110);
    wire[0:0] s13460, in13460_1, in13460_2;
    wire c13460;
    assign in13460_1 = {s12114[0]};
    assign in13460_2 = {s12115[0]};
    Full_Adder FA_13460(s13460, c13460, in13460_1, in13460_2, s12113[0]);
    wire[0:0] s13461, in13461_1, in13461_2;
    wire c13461;
    assign in13461_1 = {s12117[0]};
    assign in13461_2 = {s12118[0]};
    Full_Adder FA_13461(s13461, c13461, in13461_1, in13461_2, s12116[0]);
    wire[0:0] s13462, in13462_1, in13462_2;
    wire c13462;
    assign in13462_1 = {s10485[0]};
    assign in13462_2 = {c12111};
    Full_Adder FA_13462(s13462, c13462, in13462_1, in13462_2, s10484[0]);
    wire[0:0] s13463, in13463_1, in13463_2;
    wire c13463;
    assign in13463_1 = {c12113};
    assign in13463_2 = {c12114};
    Full_Adder FA_13463(s13463, c13463, in13463_1, in13463_2, c12112);
    wire[0:0] s13464, in13464_1, in13464_2;
    wire c13464;
    assign in13464_1 = {c12116};
    assign in13464_2 = {c12117};
    Full_Adder FA_13464(s13464, c13464, in13464_1, in13464_2, c12115);
    wire[0:0] s13465, in13465_1, in13465_2;
    wire c13465;
    assign in13465_1 = {s12119[0]};
    assign in13465_2 = {s12120[0]};
    Full_Adder FA_13465(s13465, c13465, in13465_1, in13465_2, c12118);
    wire[0:0] s13466, in13466_1, in13466_2;
    wire c13466;
    assign in13466_1 = {s12122[0]};
    assign in13466_2 = {s12123[0]};
    Full_Adder FA_13466(s13466, c13466, in13466_1, in13466_2, s12121[0]);
    wire[0:0] s13467, in13467_1, in13467_2;
    wire c13467;
    assign in13467_1 = {s12125[0]};
    assign in13467_2 = {s12126[0]};
    Full_Adder FA_13467(s13467, c13467, in13467_1, in13467_2, s12124[0]);
    wire[0:0] s13468, in13468_1, in13468_2;
    wire c13468;
    assign in13468_1 = {s10491[0]};
    assign in13468_2 = {c12119};
    Full_Adder FA_13468(s13468, c13468, in13468_1, in13468_2, s10490[0]);
    wire[0:0] s13469, in13469_1, in13469_2;
    wire c13469;
    assign in13469_1 = {c12121};
    assign in13469_2 = {c12122};
    Full_Adder FA_13469(s13469, c13469, in13469_1, in13469_2, c12120);
    wire[0:0] s13470, in13470_1, in13470_2;
    wire c13470;
    assign in13470_1 = {c12124};
    assign in13470_2 = {c12125};
    Full_Adder FA_13470(s13470, c13470, in13470_1, in13470_2, c12123);
    wire[0:0] s13471, in13471_1, in13471_2;
    wire c13471;
    assign in13471_1 = {s12127[0]};
    assign in13471_2 = {s12128[0]};
    Full_Adder FA_13471(s13471, c13471, in13471_1, in13471_2, c12126);
    wire[0:0] s13472, in13472_1, in13472_2;
    wire c13472;
    assign in13472_1 = {s12130[0]};
    assign in13472_2 = {s12131[0]};
    Full_Adder FA_13472(s13472, c13472, in13472_1, in13472_2, s12129[0]);
    wire[0:0] s13473, in13473_1, in13473_2;
    wire c13473;
    assign in13473_1 = {s12133[0]};
    assign in13473_2 = {s12134[0]};
    Full_Adder FA_13473(s13473, c13473, in13473_1, in13473_2, s12132[0]);
    wire[0:0] s13474, in13474_1, in13474_2;
    wire c13474;
    assign in13474_1 = {s10496[0]};
    assign in13474_2 = {c12127};
    Full_Adder FA_13474(s13474, c13474, in13474_1, in13474_2, s10495[0]);
    wire[0:0] s13475, in13475_1, in13475_2;
    wire c13475;
    assign in13475_1 = {c12129};
    assign in13475_2 = {c12130};
    Full_Adder FA_13475(s13475, c13475, in13475_1, in13475_2, c12128);
    wire[0:0] s13476, in13476_1, in13476_2;
    wire c13476;
    assign in13476_1 = {c12132};
    assign in13476_2 = {c12133};
    Full_Adder FA_13476(s13476, c13476, in13476_1, in13476_2, c12131);
    wire[0:0] s13477, in13477_1, in13477_2;
    wire c13477;
    assign in13477_1 = {s12135[0]};
    assign in13477_2 = {s12136[0]};
    Full_Adder FA_13477(s13477, c13477, in13477_1, in13477_2, c12134);
    wire[0:0] s13478, in13478_1, in13478_2;
    wire c13478;
    assign in13478_1 = {s12138[0]};
    assign in13478_2 = {s12139[0]};
    Full_Adder FA_13478(s13478, c13478, in13478_1, in13478_2, s12137[0]);
    wire[0:0] s13479, in13479_1, in13479_2;
    wire c13479;
    assign in13479_1 = {s12141[0]};
    assign in13479_2 = {s12142[0]};
    Full_Adder FA_13479(s13479, c13479, in13479_1, in13479_2, s12140[0]);
    wire[0:0] s13480, in13480_1, in13480_2;
    wire c13480;
    assign in13480_1 = {s10500[0]};
    assign in13480_2 = {c12135};
    Full_Adder FA_13480(s13480, c13480, in13480_1, in13480_2, s10499[0]);
    wire[0:0] s13481, in13481_1, in13481_2;
    wire c13481;
    assign in13481_1 = {c12137};
    assign in13481_2 = {c12138};
    Full_Adder FA_13481(s13481, c13481, in13481_1, in13481_2, c12136);
    wire[0:0] s13482, in13482_1, in13482_2;
    wire c13482;
    assign in13482_1 = {c12140};
    assign in13482_2 = {c12141};
    Full_Adder FA_13482(s13482, c13482, in13482_1, in13482_2, c12139);
    wire[0:0] s13483, in13483_1, in13483_2;
    wire c13483;
    assign in13483_1 = {s12143[0]};
    assign in13483_2 = {s12144[0]};
    Full_Adder FA_13483(s13483, c13483, in13483_1, in13483_2, c12142);
    wire[0:0] s13484, in13484_1, in13484_2;
    wire c13484;
    assign in13484_1 = {s12146[0]};
    assign in13484_2 = {s12147[0]};
    Full_Adder FA_13484(s13484, c13484, in13484_1, in13484_2, s12145[0]);
    wire[0:0] s13485, in13485_1, in13485_2;
    wire c13485;
    assign in13485_1 = {s12149[0]};
    assign in13485_2 = {s12150[0]};
    Full_Adder FA_13485(s13485, c13485, in13485_1, in13485_2, s12148[0]);
    wire[0:0] s13486, in13486_1, in13486_2;
    wire c13486;
    assign in13486_1 = {s10503[0]};
    assign in13486_2 = {c12143};
    Full_Adder FA_13486(s13486, c13486, in13486_1, in13486_2, s10502[0]);
    wire[0:0] s13487, in13487_1, in13487_2;
    wire c13487;
    assign in13487_1 = {c12145};
    assign in13487_2 = {c12146};
    Full_Adder FA_13487(s13487, c13487, in13487_1, in13487_2, c12144);
    wire[0:0] s13488, in13488_1, in13488_2;
    wire c13488;
    assign in13488_1 = {c12148};
    assign in13488_2 = {c12149};
    Full_Adder FA_13488(s13488, c13488, in13488_1, in13488_2, c12147);
    wire[0:0] s13489, in13489_1, in13489_2;
    wire c13489;
    assign in13489_1 = {s12151[0]};
    assign in13489_2 = {s12152[0]};
    Full_Adder FA_13489(s13489, c13489, in13489_1, in13489_2, c12150);
    wire[0:0] s13490, in13490_1, in13490_2;
    wire c13490;
    assign in13490_1 = {s12154[0]};
    assign in13490_2 = {s12155[0]};
    Full_Adder FA_13490(s13490, c13490, in13490_1, in13490_2, s12153[0]);
    wire[0:0] s13491, in13491_1, in13491_2;
    wire c13491;
    assign in13491_1 = {s12157[0]};
    assign in13491_2 = {s12158[0]};
    Full_Adder FA_13491(s13491, c13491, in13491_1, in13491_2, s12156[0]);
    wire[0:0] s13492, in13492_1, in13492_2;
    wire c13492;
    assign in13492_1 = {s10505[0]};
    assign in13492_2 = {c12151};
    Full_Adder FA_13492(s13492, c13492, in13492_1, in13492_2, s10504[0]);
    wire[0:0] s13493, in13493_1, in13493_2;
    wire c13493;
    assign in13493_1 = {c12153};
    assign in13493_2 = {c12154};
    Full_Adder FA_13493(s13493, c13493, in13493_1, in13493_2, c12152);
    wire[0:0] s13494, in13494_1, in13494_2;
    wire c13494;
    assign in13494_1 = {c12156};
    assign in13494_2 = {c12157};
    Full_Adder FA_13494(s13494, c13494, in13494_1, in13494_2, c12155);
    wire[0:0] s13495, in13495_1, in13495_2;
    wire c13495;
    assign in13495_1 = {s12159[0]};
    assign in13495_2 = {s12160[0]};
    Full_Adder FA_13495(s13495, c13495, in13495_1, in13495_2, c12158);
    wire[0:0] s13496, in13496_1, in13496_2;
    wire c13496;
    assign in13496_1 = {s12162[0]};
    assign in13496_2 = {s12163[0]};
    Full_Adder FA_13496(s13496, c13496, in13496_1, in13496_2, s12161[0]);
    wire[0:0] s13497, in13497_1, in13497_2;
    wire c13497;
    assign in13497_1 = {s12165[0]};
    assign in13497_2 = {s12166[0]};
    Full_Adder FA_13497(s13497, c13497, in13497_1, in13497_2, s12164[0]);
    wire[0:0] s13498, in13498_1, in13498_2;
    wire c13498;
    assign in13498_1 = {s10506[0]};
    assign in13498_2 = {c12159};
    Full_Adder FA_13498(s13498, c13498, in13498_1, in13498_2, c10505);
    wire[0:0] s13499, in13499_1, in13499_2;
    wire c13499;
    assign in13499_1 = {c12161};
    assign in13499_2 = {c12162};
    Full_Adder FA_13499(s13499, c13499, in13499_1, in13499_2, c12160);
    wire[0:0] s13500, in13500_1, in13500_2;
    wire c13500;
    assign in13500_1 = {c12164};
    assign in13500_2 = {c12165};
    Full_Adder FA_13500(s13500, c13500, in13500_1, in13500_2, c12163);
    wire[0:0] s13501, in13501_1, in13501_2;
    wire c13501;
    assign in13501_1 = {s12167[0]};
    assign in13501_2 = {s12168[0]};
    Full_Adder FA_13501(s13501, c13501, in13501_1, in13501_2, c12166);
    wire[0:0] s13502, in13502_1, in13502_2;
    wire c13502;
    assign in13502_1 = {s12170[0]};
    assign in13502_2 = {s12171[0]};
    Full_Adder FA_13502(s13502, c13502, in13502_1, in13502_2, s12169[0]);
    wire[0:0] s13503, in13503_1, in13503_2;
    wire c13503;
    assign in13503_1 = {s12173[0]};
    assign in13503_2 = {s12174[0]};
    Full_Adder FA_13503(s13503, c13503, in13503_1, in13503_2, s12172[0]);
    wire[0:0] s13504, in13504_1, in13504_2;
    wire c13504;
    assign in13504_1 = {c10506};
    assign in13504_2 = {c12167};
    Full_Adder FA_13504(s13504, c13504, in13504_1, in13504_2, pp127[103]);
    wire[0:0] s13505, in13505_1, in13505_2;
    wire c13505;
    assign in13505_1 = {c12169};
    assign in13505_2 = {c12170};
    Full_Adder FA_13505(s13505, c13505, in13505_1, in13505_2, c12168);
    wire[0:0] s13506, in13506_1, in13506_2;
    wire c13506;
    assign in13506_1 = {c12172};
    assign in13506_2 = {c12173};
    Full_Adder FA_13506(s13506, c13506, in13506_1, in13506_2, c12171);
    wire[0:0] s13507, in13507_1, in13507_2;
    wire c13507;
    assign in13507_1 = {s12175[0]};
    assign in13507_2 = {s12176[0]};
    Full_Adder FA_13507(s13507, c13507, in13507_1, in13507_2, c12174);
    wire[0:0] s13508, in13508_1, in13508_2;
    wire c13508;
    assign in13508_1 = {s12178[0]};
    assign in13508_2 = {s12179[0]};
    Full_Adder FA_13508(s13508, c13508, in13508_1, in13508_2, s12177[0]);
    wire[0:0] s13509, in13509_1, in13509_2;
    wire c13509;
    assign in13509_1 = {s12181[0]};
    assign in13509_2 = {s12182[0]};
    Full_Adder FA_13509(s13509, c13509, in13509_1, in13509_2, s12180[0]);
    wire[0:0] s13510, in13510_1, in13510_2;
    wire c13510;
    assign in13510_1 = {pp126[105]};
    assign in13510_2 = {pp127[104]};
    Full_Adder FA_13510(s13510, c13510, in13510_1, in13510_2, pp125[106]);
    wire[0:0] s13511, in13511_1, in13511_2;
    wire c13511;
    assign in13511_1 = {c12176};
    assign in13511_2 = {c12177};
    Full_Adder FA_13511(s13511, c13511, in13511_1, in13511_2, c12175);
    wire[0:0] s13512, in13512_1, in13512_2;
    wire c13512;
    assign in13512_1 = {c12179};
    assign in13512_2 = {c12180};
    Full_Adder FA_13512(s13512, c13512, in13512_1, in13512_2, c12178);
    wire[0:0] s13513, in13513_1, in13513_2;
    wire c13513;
    assign in13513_1 = {c12182};
    assign in13513_2 = {s12183[0]};
    Full_Adder FA_13513(s13513, c13513, in13513_1, in13513_2, c12181);
    wire[0:0] s13514, in13514_1, in13514_2;
    wire c13514;
    assign in13514_1 = {s12185[0]};
    assign in13514_2 = {s12186[0]};
    Full_Adder FA_13514(s13514, c13514, in13514_1, in13514_2, s12184[0]);
    wire[0:0] s13515, in13515_1, in13515_2;
    wire c13515;
    assign in13515_1 = {s12188[0]};
    assign in13515_2 = {s12189[0]};
    Full_Adder FA_13515(s13515, c13515, in13515_1, in13515_2, s12187[0]);
    wire[0:0] s13516, in13516_1, in13516_2;
    wire c13516;
    assign in13516_1 = {pp124[108]};
    assign in13516_2 = {pp125[107]};
    Full_Adder FA_13516(s13516, c13516, in13516_1, in13516_2, pp123[109]);
    wire[0:0] s13517, in13517_1, in13517_2;
    wire c13517;
    assign in13517_1 = {pp127[105]};
    assign in13517_2 = {c12183};
    Full_Adder FA_13517(s13517, c13517, in13517_1, in13517_2, pp126[106]);
    wire[0:0] s13518, in13518_1, in13518_2;
    wire c13518;
    assign in13518_1 = {c12185};
    assign in13518_2 = {c12186};
    Full_Adder FA_13518(s13518, c13518, in13518_1, in13518_2, c12184);
    wire[0:0] s13519, in13519_1, in13519_2;
    wire c13519;
    assign in13519_1 = {c12188};
    assign in13519_2 = {c12189};
    Full_Adder FA_13519(s13519, c13519, in13519_1, in13519_2, c12187);
    wire[0:0] s13520, in13520_1, in13520_2;
    wire c13520;
    assign in13520_1 = {s12191[0]};
    assign in13520_2 = {s12192[0]};
    Full_Adder FA_13520(s13520, c13520, in13520_1, in13520_2, s12190[0]);
    wire[0:0] s13521, in13521_1, in13521_2;
    wire c13521;
    assign in13521_1 = {s12194[0]};
    assign in13521_2 = {s12195[0]};
    Full_Adder FA_13521(s13521, c13521, in13521_1, in13521_2, s12193[0]);
    wire[0:0] s13522, in13522_1, in13522_2;
    wire c13522;
    assign in13522_1 = {pp122[111]};
    assign in13522_2 = {pp123[110]};
    Full_Adder FA_13522(s13522, c13522, in13522_1, in13522_2, pp121[112]);
    wire[0:0] s13523, in13523_1, in13523_2;
    wire c13523;
    assign in13523_1 = {pp125[108]};
    assign in13523_2 = {pp126[107]};
    Full_Adder FA_13523(s13523, c13523, in13523_1, in13523_2, pp124[109]);
    wire[0:0] s13524, in13524_1, in13524_2;
    wire c13524;
    assign in13524_1 = {c12190};
    assign in13524_2 = {c12191};
    Full_Adder FA_13524(s13524, c13524, in13524_1, in13524_2, pp127[106]);
    wire[0:0] s13525, in13525_1, in13525_2;
    wire c13525;
    assign in13525_1 = {c12193};
    assign in13525_2 = {c12194};
    Full_Adder FA_13525(s13525, c13525, in13525_1, in13525_2, c12192);
    wire[0:0] s13526, in13526_1, in13526_2;
    wire c13526;
    assign in13526_1 = {s12196[0]};
    assign in13526_2 = {s12197[0]};
    Full_Adder FA_13526(s13526, c13526, in13526_1, in13526_2, c12195);
    wire[0:0] s13527, in13527_1, in13527_2;
    wire c13527;
    assign in13527_1 = {s12199[0]};
    assign in13527_2 = {s12200[0]};
    Full_Adder FA_13527(s13527, c13527, in13527_1, in13527_2, s12198[0]);
    wire[0:0] s13528, in13528_1, in13528_2;
    wire c13528;
    assign in13528_1 = {pp120[114]};
    assign in13528_2 = {pp121[113]};
    Full_Adder FA_13528(s13528, c13528, in13528_1, in13528_2, pp119[115]);
    wire[0:0] s13529, in13529_1, in13529_2;
    wire c13529;
    assign in13529_1 = {pp123[111]};
    assign in13529_2 = {pp124[110]};
    Full_Adder FA_13529(s13529, c13529, in13529_1, in13529_2, pp122[112]);
    wire[0:0] s13530, in13530_1, in13530_2;
    wire c13530;
    assign in13530_1 = {pp126[108]};
    assign in13530_2 = {pp127[107]};
    Full_Adder FA_13530(s13530, c13530, in13530_1, in13530_2, pp125[109]);
    wire[0:0] s13531, in13531_1, in13531_2;
    wire c13531;
    assign in13531_1 = {c12197};
    assign in13531_2 = {c12198};
    Full_Adder FA_13531(s13531, c13531, in13531_1, in13531_2, c12196);
    wire[0:0] s13532, in13532_1, in13532_2;
    wire c13532;
    assign in13532_1 = {c12200};
    assign in13532_2 = {s12201[0]};
    Full_Adder FA_13532(s13532, c13532, in13532_1, in13532_2, c12199);
    wire[0:0] s13533, in13533_1, in13533_2;
    wire c13533;
    assign in13533_1 = {s12203[0]};
    assign in13533_2 = {s12204[0]};
    Full_Adder FA_13533(s13533, c13533, in13533_1, in13533_2, s12202[0]);
    wire[0:0] s13534, in13534_1, in13534_2;
    wire c13534;
    assign in13534_1 = {pp118[117]};
    assign in13534_2 = {pp119[116]};
    Full_Adder FA_13534(s13534, c13534, in13534_1, in13534_2, pp117[118]);
    wire[0:0] s13535, in13535_1, in13535_2;
    wire c13535;
    assign in13535_1 = {pp121[114]};
    assign in13535_2 = {pp122[113]};
    Full_Adder FA_13535(s13535, c13535, in13535_1, in13535_2, pp120[115]);
    wire[0:0] s13536, in13536_1, in13536_2;
    wire c13536;
    assign in13536_1 = {pp124[111]};
    assign in13536_2 = {pp125[110]};
    Full_Adder FA_13536(s13536, c13536, in13536_1, in13536_2, pp123[112]);
    wire[0:0] s13537, in13537_1, in13537_2;
    wire c13537;
    assign in13537_1 = {pp127[108]};
    assign in13537_2 = {c12201};
    Full_Adder FA_13537(s13537, c13537, in13537_1, in13537_2, pp126[109]);
    wire[0:0] s13538, in13538_1, in13538_2;
    wire c13538;
    assign in13538_1 = {c12203};
    assign in13538_2 = {c12204};
    Full_Adder FA_13538(s13538, c13538, in13538_1, in13538_2, c12202);
    wire[0:0] s13539, in13539_1, in13539_2;
    wire c13539;
    assign in13539_1 = {s12206[0]};
    assign in13539_2 = {s12207[0]};
    Full_Adder FA_13539(s13539, c13539, in13539_1, in13539_2, s12205[0]);
    wire[0:0] s13540, in13540_1, in13540_2;
    wire c13540;
    assign in13540_1 = {pp116[120]};
    assign in13540_2 = {pp117[119]};
    Full_Adder FA_13540(s13540, c13540, in13540_1, in13540_2, pp115[121]);
    wire[0:0] s13541, in13541_1, in13541_2;
    wire c13541;
    assign in13541_1 = {pp119[117]};
    assign in13541_2 = {pp120[116]};
    Full_Adder FA_13541(s13541, c13541, in13541_1, in13541_2, pp118[118]);
    wire[0:0] s13542, in13542_1, in13542_2;
    wire c13542;
    assign in13542_1 = {pp122[114]};
    assign in13542_2 = {pp123[113]};
    Full_Adder FA_13542(s13542, c13542, in13542_1, in13542_2, pp121[115]);
    wire[0:0] s13543, in13543_1, in13543_2;
    wire c13543;
    assign in13543_1 = {pp125[111]};
    assign in13543_2 = {pp126[110]};
    Full_Adder FA_13543(s13543, c13543, in13543_1, in13543_2, pp124[112]);
    wire[0:0] s13544, in13544_1, in13544_2;
    wire c13544;
    assign in13544_1 = {c12205};
    assign in13544_2 = {c12206};
    Full_Adder FA_13544(s13544, c13544, in13544_1, in13544_2, pp127[109]);
    wire[0:0] s13545, in13545_1, in13545_2;
    wire c13545;
    assign in13545_1 = {s12208[0]};
    assign in13545_2 = {s12209[0]};
    Full_Adder FA_13545(s13545, c13545, in13545_1, in13545_2, c12207);
    wire[0:0] s13546, in13546_1, in13546_2;
    wire c13546;
    assign in13546_1 = {pp114[123]};
    assign in13546_2 = {pp115[122]};
    Full_Adder FA_13546(s13546, c13546, in13546_1, in13546_2, pp113[124]);
    wire[0:0] s13547, in13547_1, in13547_2;
    wire c13547;
    assign in13547_1 = {pp117[120]};
    assign in13547_2 = {pp118[119]};
    Full_Adder FA_13547(s13547, c13547, in13547_1, in13547_2, pp116[121]);
    wire[0:0] s13548, in13548_1, in13548_2;
    wire c13548;
    assign in13548_1 = {pp120[117]};
    assign in13548_2 = {pp121[116]};
    Full_Adder FA_13548(s13548, c13548, in13548_1, in13548_2, pp119[118]);
    wire[0:0] s13549, in13549_1, in13549_2;
    wire c13549;
    assign in13549_1 = {pp123[114]};
    assign in13549_2 = {pp124[113]};
    Full_Adder FA_13549(s13549, c13549, in13549_1, in13549_2, pp122[115]);
    wire[0:0] s13550, in13550_1, in13550_2;
    wire c13550;
    assign in13550_1 = {pp126[111]};
    assign in13550_2 = {pp127[110]};
    Full_Adder FA_13550(s13550, c13550, in13550_1, in13550_2, pp125[112]);
    wire[0:0] s13551, in13551_1, in13551_2;
    wire c13551;
    assign in13551_1 = {c12209};
    assign in13551_2 = {s12210[0]};
    Full_Adder FA_13551(s13551, c13551, in13551_1, in13551_2, c12208);
    wire[0:0] s13552, in13552_1, in13552_2;
    wire c13552;
    assign in13552_1 = {pp112[126]};
    assign in13552_2 = {pp113[125]};
    Full_Adder FA_13552(s13552, c13552, in13552_1, in13552_2, pp111[127]);
    wire[0:0] s13553, in13553_1, in13553_2;
    wire c13553;
    assign in13553_1 = {pp115[123]};
    assign in13553_2 = {pp116[122]};
    Full_Adder FA_13553(s13553, c13553, in13553_1, in13553_2, pp114[124]);
    wire[0:0] s13554, in13554_1, in13554_2;
    wire c13554;
    assign in13554_1 = {pp118[120]};
    assign in13554_2 = {pp119[119]};
    Full_Adder FA_13554(s13554, c13554, in13554_1, in13554_2, pp117[121]);
    wire[0:0] s13555, in13555_1, in13555_2;
    wire c13555;
    assign in13555_1 = {pp121[117]};
    assign in13555_2 = {pp122[116]};
    Full_Adder FA_13555(s13555, c13555, in13555_1, in13555_2, pp120[118]);
    wire[0:0] s13556, in13556_1, in13556_2;
    wire c13556;
    assign in13556_1 = {pp124[114]};
    assign in13556_2 = {pp125[113]};
    Full_Adder FA_13556(s13556, c13556, in13556_1, in13556_2, pp123[115]);
    wire[0:0] s13557, in13557_1, in13557_2;
    wire c13557;
    assign in13557_1 = {pp127[111]};
    assign in13557_2 = {c12210};
    Full_Adder FA_13557(s13557, c13557, in13557_1, in13557_2, pp126[112]);
    wire[0:0] s13558, in13558_1, in13558_2;
    wire c13558;
    assign in13558_1 = {pp113[126]};
    assign in13558_2 = {pp114[125]};
    Full_Adder FA_13558(s13558, c13558, in13558_1, in13558_2, pp112[127]);
    wire[0:0] s13559, in13559_1, in13559_2;
    wire c13559;
    assign in13559_1 = {pp116[123]};
    assign in13559_2 = {pp117[122]};
    Full_Adder FA_13559(s13559, c13559, in13559_1, in13559_2, pp115[124]);
    wire[0:0] s13560, in13560_1, in13560_2;
    wire c13560;
    assign in13560_1 = {pp119[120]};
    assign in13560_2 = {pp120[119]};
    Full_Adder FA_13560(s13560, c13560, in13560_1, in13560_2, pp118[121]);
    wire[0:0] s13561, in13561_1, in13561_2;
    wire c13561;
    assign in13561_1 = {pp122[117]};
    assign in13561_2 = {pp123[116]};
    Full_Adder FA_13561(s13561, c13561, in13561_1, in13561_2, pp121[118]);
    wire[0:0] s13562, in13562_1, in13562_2;
    wire c13562;
    assign in13562_1 = {pp125[114]};
    assign in13562_2 = {pp126[113]};
    Full_Adder FA_13562(s13562, c13562, in13562_1, in13562_2, pp124[115]);
    wire[0:0] s13563, in13563_1, in13563_2;
    wire c13563;
    assign in13563_1 = {pp114[126]};
    assign in13563_2 = {pp115[125]};
    Full_Adder FA_13563(s13563, c13563, in13563_1, in13563_2, pp113[127]);
    wire[0:0] s13564, in13564_1, in13564_2;
    wire c13564;
    assign in13564_1 = {pp117[123]};
    assign in13564_2 = {pp118[122]};
    Full_Adder FA_13564(s13564, c13564, in13564_1, in13564_2, pp116[124]);
    wire[0:0] s13565, in13565_1, in13565_2;
    wire c13565;
    assign in13565_1 = {pp120[120]};
    assign in13565_2 = {pp121[119]};
    Full_Adder FA_13565(s13565, c13565, in13565_1, in13565_2, pp119[121]);
    wire[0:0] s13566, in13566_1, in13566_2;
    wire c13566;
    assign in13566_1 = {pp123[117]};
    assign in13566_2 = {pp124[116]};
    Full_Adder FA_13566(s13566, c13566, in13566_1, in13566_2, pp122[118]);
    wire[0:0] s13567, in13567_1, in13567_2;
    wire c13567;
    assign in13567_1 = {pp115[126]};
    assign in13567_2 = {pp116[125]};
    Full_Adder FA_13567(s13567, c13567, in13567_1, in13567_2, pp114[127]);
    wire[0:0] s13568, in13568_1, in13568_2;
    wire c13568;
    assign in13568_1 = {pp118[123]};
    assign in13568_2 = {pp119[122]};
    Full_Adder FA_13568(s13568, c13568, in13568_1, in13568_2, pp117[124]);
    wire[0:0] s13569, in13569_1, in13569_2;
    wire c13569;
    assign in13569_1 = {pp121[120]};
    assign in13569_2 = {pp122[119]};
    Full_Adder FA_13569(s13569, c13569, in13569_1, in13569_2, pp120[121]);
    wire[0:0] s13570, in13570_1, in13570_2;
    wire c13570;
    assign in13570_1 = {pp116[126]};
    assign in13570_2 = {pp117[125]};
    Full_Adder FA_13570(s13570, c13570, in13570_1, in13570_2, pp115[127]);
    wire[0:0] s13571, in13571_1, in13571_2;
    wire c13571;
    assign in13571_1 = {pp119[123]};
    assign in13571_2 = {pp120[122]};
    Full_Adder FA_13571(s13571, c13571, in13571_1, in13571_2, pp118[124]);
    wire[0:0] s13572, in13572_1, in13572_2;
    wire c13572;
    assign in13572_1 = {pp117[126]};
    assign in13572_2 = {pp118[125]};
    Full_Adder FA_13572(s13572, c13572, in13572_1, in13572_2, pp116[127]);

    /*Stage 7*/
    wire[0:0] s13573, in13573_1, in13573_2;
    wire c13573;
    assign in13573_1 = {pp0[8]};
    assign in13573_2 = {pp1[7]};
    Half_Adder HA_13573(s13573, c13573, in13573_1, in13573_2);
    wire[0:0] s13574, in13574_1, in13574_2;
    wire c13574;
    assign in13574_1 = {pp1[8]};
    assign in13574_2 = {pp2[7]};
    Full_Adder FA_13574(s13574, c13574, in13574_1, in13574_2, pp0[9]);
    wire[0:0] s13575, in13575_1, in13575_2;
    wire c13575;
    assign in13575_1 = {pp3[6]};
    assign in13575_2 = {pp4[5]};
    Half_Adder HA_13575(s13575, c13575, in13575_1, in13575_2);
    wire[0:0] s13576, in13576_1, in13576_2;
    wire c13576;
    assign in13576_1 = {pp1[9]};
    assign in13576_2 = {pp2[8]};
    Full_Adder FA_13576(s13576, c13576, in13576_1, in13576_2, pp0[10]);
    wire[0:0] s13577, in13577_1, in13577_2;
    wire c13577;
    assign in13577_1 = {pp4[6]};
    assign in13577_2 = {pp5[5]};
    Full_Adder FA_13577(s13577, c13577, in13577_1, in13577_2, pp3[7]);
    wire[0:0] s13578, in13578_1, in13578_2;
    wire c13578;
    assign in13578_1 = {pp6[4]};
    assign in13578_2 = {pp7[3]};
    Half_Adder HA_13578(s13578, c13578, in13578_1, in13578_2);
    wire[0:0] s13579, in13579_1, in13579_2;
    wire c13579;
    assign in13579_1 = {pp1[10]};
    assign in13579_2 = {pp2[9]};
    Full_Adder FA_13579(s13579, c13579, in13579_1, in13579_2, pp0[11]);
    wire[0:0] s13580, in13580_1, in13580_2;
    wire c13580;
    assign in13580_1 = {pp4[7]};
    assign in13580_2 = {pp5[6]};
    Full_Adder FA_13580(s13580, c13580, in13580_1, in13580_2, pp3[8]);
    wire[0:0] s13581, in13581_1, in13581_2;
    wire c13581;
    assign in13581_1 = {pp7[4]};
    assign in13581_2 = {pp8[3]};
    Full_Adder FA_13581(s13581, c13581, in13581_1, in13581_2, pp6[5]);
    wire[0:0] s13582, in13582_1, in13582_2;
    wire c13582;
    assign in13582_1 = {pp9[2]};
    assign in13582_2 = {pp10[1]};
    Half_Adder HA_13582(s13582, c13582, in13582_1, in13582_2);
    wire[0:0] s13583, in13583_1, in13583_2;
    wire c13583;
    assign in13583_1 = {pp3[9]};
    assign in13583_2 = {pp4[8]};
    Full_Adder FA_13583(s13583, c13583, in13583_1, in13583_2, pp2[10]);
    wire[0:0] s13584, in13584_1, in13584_2;
    wire c13584;
    assign in13584_1 = {pp6[6]};
    assign in13584_2 = {pp7[5]};
    Full_Adder FA_13584(s13584, c13584, in13584_1, in13584_2, pp5[7]);
    wire[0:0] s13585, in13585_1, in13585_2;
    wire c13585;
    assign in13585_1 = {pp9[3]};
    assign in13585_2 = {pp10[2]};
    Full_Adder FA_13585(s13585, c13585, in13585_1, in13585_2, pp8[4]);
    wire[0:0] s13586, in13586_1, in13586_2;
    wire c13586;
    assign in13586_1 = {pp12[0]};
    assign in13586_2 = {s12211[0]};
    Full_Adder FA_13586(s13586, c13586, in13586_1, in13586_2, pp11[1]);
    wire[0:0] s13587, in13587_1, in13587_2;
    wire c13587;
    assign in13587_1 = {pp6[7]};
    assign in13587_2 = {pp7[6]};
    Full_Adder FA_13587(s13587, c13587, in13587_1, in13587_2, pp5[8]);
    wire[0:0] s13588, in13588_1, in13588_2;
    wire c13588;
    assign in13588_1 = {pp9[4]};
    assign in13588_2 = {pp10[3]};
    Full_Adder FA_13588(s13588, c13588, in13588_1, in13588_2, pp8[5]);
    wire[0:0] s13589, in13589_1, in13589_2;
    wire c13589;
    assign in13589_1 = {pp12[1]};
    assign in13589_2 = {pp13[0]};
    Full_Adder FA_13589(s13589, c13589, in13589_1, in13589_2, pp11[2]);
    wire[0:0] s13590, in13590_1, in13590_2;
    wire c13590;
    assign in13590_1 = {s12212[0]};
    assign in13590_2 = {s12213[0]};
    Full_Adder FA_13590(s13590, c13590, in13590_1, in13590_2, c12211);
    wire[0:0] s13591, in13591_1, in13591_2;
    wire c13591;
    assign in13591_1 = {pp9[5]};
    assign in13591_2 = {pp10[4]};
    Full_Adder FA_13591(s13591, c13591, in13591_1, in13591_2, pp8[6]);
    wire[0:0] s13592, in13592_1, in13592_2;
    wire c13592;
    assign in13592_1 = {pp12[2]};
    assign in13592_2 = {pp13[1]};
    Full_Adder FA_13592(s13592, c13592, in13592_1, in13592_2, pp11[3]);
    wire[0:0] s13593, in13593_1, in13593_2;
    wire c13593;
    assign in13593_1 = {c12212};
    assign in13593_2 = {c12213};
    Full_Adder FA_13593(s13593, c13593, in13593_1, in13593_2, pp14[0]);
    wire[0:0] s13594, in13594_1, in13594_2;
    wire c13594;
    assign in13594_1 = {s12215[0]};
    assign in13594_2 = {s12216[0]};
    Full_Adder FA_13594(s13594, c13594, in13594_1, in13594_2, s12214[0]);
    wire[0:0] s13595, in13595_1, in13595_2;
    wire c13595;
    assign in13595_1 = {pp12[3]};
    assign in13595_2 = {pp13[2]};
    Full_Adder FA_13595(s13595, c13595, in13595_1, in13595_2, pp11[4]);
    wire[0:0] s13596, in13596_1, in13596_2;
    wire c13596;
    assign in13596_1 = {pp15[0]};
    assign in13596_2 = {c12214};
    Full_Adder FA_13596(s13596, c13596, in13596_1, in13596_2, pp14[1]);
    wire[0:0] s13597, in13597_1, in13597_2;
    wire c13597;
    assign in13597_1 = {c12216};
    assign in13597_2 = {s12217[0]};
    Full_Adder FA_13597(s13597, c13597, in13597_1, in13597_2, c12215);
    wire[0:0] s13598, in13598_1, in13598_2;
    wire c13598;
    assign in13598_1 = {s12219[0]};
    assign in13598_2 = {s12220[0]};
    Full_Adder FA_13598(s13598, c13598, in13598_1, in13598_2, s12218[0]);
    wire[0:0] s13599, in13599_1, in13599_2;
    wire c13599;
    assign in13599_1 = {pp15[1]};
    assign in13599_2 = {pp16[0]};
    Full_Adder FA_13599(s13599, c13599, in13599_1, in13599_2, pp14[2]);
    wire[0:0] s13600, in13600_1, in13600_2;
    wire c13600;
    assign in13600_1 = {c12218};
    assign in13600_2 = {c12219};
    Full_Adder FA_13600(s13600, c13600, in13600_1, in13600_2, c12217);
    wire[0:0] s13601, in13601_1, in13601_2;
    wire c13601;
    assign in13601_1 = {s12221[0]};
    assign in13601_2 = {s12222[0]};
    Full_Adder FA_13601(s13601, c13601, in13601_1, in13601_2, c12220);
    wire[0:0] s13602, in13602_1, in13602_2;
    wire c13602;
    assign in13602_1 = {s12224[0]};
    assign in13602_2 = {s12225[0]};
    Full_Adder FA_13602(s13602, c13602, in13602_1, in13602_2, s12223[0]);
    wire[0:0] s13603, in13603_1, in13603_2;
    wire c13603;
    assign in13603_1 = {c12221};
    assign in13603_2 = {c12222};
    Full_Adder FA_13603(s13603, c13603, in13603_1, in13603_2, pp17[0]);
    wire[0:0] s13604, in13604_1, in13604_2;
    wire c13604;
    assign in13604_1 = {c12224};
    assign in13604_2 = {c12225};
    Full_Adder FA_13604(s13604, c13604, in13604_1, in13604_2, c12223);
    wire[0:0] s13605, in13605_1, in13605_2;
    wire c13605;
    assign in13605_1 = {s12227[0]};
    assign in13605_2 = {s12228[0]};
    Full_Adder FA_13605(s13605, c13605, in13605_1, in13605_2, s12226[0]);
    wire[0:0] s13606, in13606_1, in13606_2;
    wire c13606;
    assign in13606_1 = {s12230[0]};
    assign in13606_2 = {s12231[0]};
    Full_Adder FA_13606(s13606, c13606, in13606_1, in13606_2, s12229[0]);
    wire[0:0] s13607, in13607_1, in13607_2;
    wire c13607;
    assign in13607_1 = {c12227};
    assign in13607_2 = {c12228};
    Full_Adder FA_13607(s13607, c13607, in13607_1, in13607_2, c12226);
    wire[0:0] s13608, in13608_1, in13608_2;
    wire c13608;
    assign in13608_1 = {c12230};
    assign in13608_2 = {c12231};
    Full_Adder FA_13608(s13608, c13608, in13608_1, in13608_2, c12229);
    wire[0:0] s13609, in13609_1, in13609_2;
    wire c13609;
    assign in13609_1 = {s12233[0]};
    assign in13609_2 = {s12234[0]};
    Full_Adder FA_13609(s13609, c13609, in13609_1, in13609_2, s12232[0]);
    wire[0:0] s13610, in13610_1, in13610_2;
    wire c13610;
    assign in13610_1 = {s12236[0]};
    assign in13610_2 = {s12237[0]};
    Full_Adder FA_13610(s13610, c13610, in13610_1, in13610_2, s12235[0]);
    wire[0:0] s13611, in13611_1, in13611_2;
    wire c13611;
    assign in13611_1 = {c12233};
    assign in13611_2 = {c12234};
    Full_Adder FA_13611(s13611, c13611, in13611_1, in13611_2, c12232);
    wire[0:0] s13612, in13612_1, in13612_2;
    wire c13612;
    assign in13612_1 = {c12236};
    assign in13612_2 = {c12237};
    Full_Adder FA_13612(s13612, c13612, in13612_1, in13612_2, c12235);
    wire[0:0] s13613, in13613_1, in13613_2;
    wire c13613;
    assign in13613_1 = {s12239[0]};
    assign in13613_2 = {s12240[0]};
    Full_Adder FA_13613(s13613, c13613, in13613_1, in13613_2, s12238[0]);
    wire[0:0] s13614, in13614_1, in13614_2;
    wire c13614;
    assign in13614_1 = {s12242[0]};
    assign in13614_2 = {s12243[0]};
    Full_Adder FA_13614(s13614, c13614, in13614_1, in13614_2, s12241[0]);
    wire[0:0] s13615, in13615_1, in13615_2;
    wire c13615;
    assign in13615_1 = {c12239};
    assign in13615_2 = {c12240};
    Full_Adder FA_13615(s13615, c13615, in13615_1, in13615_2, c12238);
    wire[0:0] s13616, in13616_1, in13616_2;
    wire c13616;
    assign in13616_1 = {c12242};
    assign in13616_2 = {c12243};
    Full_Adder FA_13616(s13616, c13616, in13616_1, in13616_2, c12241);
    wire[0:0] s13617, in13617_1, in13617_2;
    wire c13617;
    assign in13617_1 = {s12245[0]};
    assign in13617_2 = {s12246[0]};
    Full_Adder FA_13617(s13617, c13617, in13617_1, in13617_2, s12244[0]);
    wire[0:0] s13618, in13618_1, in13618_2;
    wire c13618;
    assign in13618_1 = {s12248[0]};
    assign in13618_2 = {s12249[0]};
    Full_Adder FA_13618(s13618, c13618, in13618_1, in13618_2, s12247[0]);
    wire[0:0] s13619, in13619_1, in13619_2;
    wire c13619;
    assign in13619_1 = {c12245};
    assign in13619_2 = {c12246};
    Full_Adder FA_13619(s13619, c13619, in13619_1, in13619_2, c12244);
    wire[0:0] s13620, in13620_1, in13620_2;
    wire c13620;
    assign in13620_1 = {c12248};
    assign in13620_2 = {c12249};
    Full_Adder FA_13620(s13620, c13620, in13620_1, in13620_2, c12247);
    wire[0:0] s13621, in13621_1, in13621_2;
    wire c13621;
    assign in13621_1 = {s12251[0]};
    assign in13621_2 = {s12252[0]};
    Full_Adder FA_13621(s13621, c13621, in13621_1, in13621_2, s12250[0]);
    wire[0:0] s13622, in13622_1, in13622_2;
    wire c13622;
    assign in13622_1 = {s12254[0]};
    assign in13622_2 = {s12255[0]};
    Full_Adder FA_13622(s13622, c13622, in13622_1, in13622_2, s12253[0]);
    wire[0:0] s13623, in13623_1, in13623_2;
    wire c13623;
    assign in13623_1 = {c12251};
    assign in13623_2 = {c12252};
    Full_Adder FA_13623(s13623, c13623, in13623_1, in13623_2, c12250);
    wire[0:0] s13624, in13624_1, in13624_2;
    wire c13624;
    assign in13624_1 = {c12254};
    assign in13624_2 = {c12255};
    Full_Adder FA_13624(s13624, c13624, in13624_1, in13624_2, c12253);
    wire[0:0] s13625, in13625_1, in13625_2;
    wire c13625;
    assign in13625_1 = {s12257[0]};
    assign in13625_2 = {s12258[0]};
    Full_Adder FA_13625(s13625, c13625, in13625_1, in13625_2, s12256[0]);
    wire[0:0] s13626, in13626_1, in13626_2;
    wire c13626;
    assign in13626_1 = {s12260[0]};
    assign in13626_2 = {s12261[0]};
    Full_Adder FA_13626(s13626, c13626, in13626_1, in13626_2, s12259[0]);
    wire[0:0] s13627, in13627_1, in13627_2;
    wire c13627;
    assign in13627_1 = {c12257};
    assign in13627_2 = {c12258};
    Full_Adder FA_13627(s13627, c13627, in13627_1, in13627_2, c12256);
    wire[0:0] s13628, in13628_1, in13628_2;
    wire c13628;
    assign in13628_1 = {c12260};
    assign in13628_2 = {c12261};
    Full_Adder FA_13628(s13628, c13628, in13628_1, in13628_2, c12259);
    wire[0:0] s13629, in13629_1, in13629_2;
    wire c13629;
    assign in13629_1 = {s12263[0]};
    assign in13629_2 = {s12264[0]};
    Full_Adder FA_13629(s13629, c13629, in13629_1, in13629_2, s12262[0]);
    wire[0:0] s13630, in13630_1, in13630_2;
    wire c13630;
    assign in13630_1 = {s12266[0]};
    assign in13630_2 = {s12267[0]};
    Full_Adder FA_13630(s13630, c13630, in13630_1, in13630_2, s12265[0]);
    wire[0:0] s13631, in13631_1, in13631_2;
    wire c13631;
    assign in13631_1 = {c12263};
    assign in13631_2 = {c12264};
    Full_Adder FA_13631(s13631, c13631, in13631_1, in13631_2, c12262);
    wire[0:0] s13632, in13632_1, in13632_2;
    wire c13632;
    assign in13632_1 = {c12266};
    assign in13632_2 = {c12267};
    Full_Adder FA_13632(s13632, c13632, in13632_1, in13632_2, c12265);
    wire[0:0] s13633, in13633_1, in13633_2;
    wire c13633;
    assign in13633_1 = {s12269[0]};
    assign in13633_2 = {s12270[0]};
    Full_Adder FA_13633(s13633, c13633, in13633_1, in13633_2, s12268[0]);
    wire[0:0] s13634, in13634_1, in13634_2;
    wire c13634;
    assign in13634_1 = {s12272[0]};
    assign in13634_2 = {s12273[0]};
    Full_Adder FA_13634(s13634, c13634, in13634_1, in13634_2, s12271[0]);
    wire[0:0] s13635, in13635_1, in13635_2;
    wire c13635;
    assign in13635_1 = {c12269};
    assign in13635_2 = {c12270};
    Full_Adder FA_13635(s13635, c13635, in13635_1, in13635_2, c12268);
    wire[0:0] s13636, in13636_1, in13636_2;
    wire c13636;
    assign in13636_1 = {c12272};
    assign in13636_2 = {c12273};
    Full_Adder FA_13636(s13636, c13636, in13636_1, in13636_2, c12271);
    wire[0:0] s13637, in13637_1, in13637_2;
    wire c13637;
    assign in13637_1 = {s12275[0]};
    assign in13637_2 = {s12276[0]};
    Full_Adder FA_13637(s13637, c13637, in13637_1, in13637_2, s12274[0]);
    wire[0:0] s13638, in13638_1, in13638_2;
    wire c13638;
    assign in13638_1 = {s12278[0]};
    assign in13638_2 = {s12279[0]};
    Full_Adder FA_13638(s13638, c13638, in13638_1, in13638_2, s12277[0]);
    wire[0:0] s13639, in13639_1, in13639_2;
    wire c13639;
    assign in13639_1 = {c12275};
    assign in13639_2 = {c12276};
    Full_Adder FA_13639(s13639, c13639, in13639_1, in13639_2, c12274);
    wire[0:0] s13640, in13640_1, in13640_2;
    wire c13640;
    assign in13640_1 = {c12278};
    assign in13640_2 = {c12279};
    Full_Adder FA_13640(s13640, c13640, in13640_1, in13640_2, c12277);
    wire[0:0] s13641, in13641_1, in13641_2;
    wire c13641;
    assign in13641_1 = {s12281[0]};
    assign in13641_2 = {s12282[0]};
    Full_Adder FA_13641(s13641, c13641, in13641_1, in13641_2, s12280[0]);
    wire[0:0] s13642, in13642_1, in13642_2;
    wire c13642;
    assign in13642_1 = {s12284[0]};
    assign in13642_2 = {s12285[0]};
    Full_Adder FA_13642(s13642, c13642, in13642_1, in13642_2, s12283[0]);
    wire[0:0] s13643, in13643_1, in13643_2;
    wire c13643;
    assign in13643_1 = {c12281};
    assign in13643_2 = {c12282};
    Full_Adder FA_13643(s13643, c13643, in13643_1, in13643_2, c12280);
    wire[0:0] s13644, in13644_1, in13644_2;
    wire c13644;
    assign in13644_1 = {c12284};
    assign in13644_2 = {c12285};
    Full_Adder FA_13644(s13644, c13644, in13644_1, in13644_2, c12283);
    wire[0:0] s13645, in13645_1, in13645_2;
    wire c13645;
    assign in13645_1 = {s12287[0]};
    assign in13645_2 = {s12288[0]};
    Full_Adder FA_13645(s13645, c13645, in13645_1, in13645_2, s12286[0]);
    wire[0:0] s13646, in13646_1, in13646_2;
    wire c13646;
    assign in13646_1 = {s12290[0]};
    assign in13646_2 = {s12291[0]};
    Full_Adder FA_13646(s13646, c13646, in13646_1, in13646_2, s12289[0]);
    wire[0:0] s13647, in13647_1, in13647_2;
    wire c13647;
    assign in13647_1 = {c12287};
    assign in13647_2 = {c12288};
    Full_Adder FA_13647(s13647, c13647, in13647_1, in13647_2, c12286);
    wire[0:0] s13648, in13648_1, in13648_2;
    wire c13648;
    assign in13648_1 = {c12290};
    assign in13648_2 = {c12291};
    Full_Adder FA_13648(s13648, c13648, in13648_1, in13648_2, c12289);
    wire[0:0] s13649, in13649_1, in13649_2;
    wire c13649;
    assign in13649_1 = {s12293[0]};
    assign in13649_2 = {s12294[0]};
    Full_Adder FA_13649(s13649, c13649, in13649_1, in13649_2, s12292[0]);
    wire[0:0] s13650, in13650_1, in13650_2;
    wire c13650;
    assign in13650_1 = {s12296[0]};
    assign in13650_2 = {s12297[0]};
    Full_Adder FA_13650(s13650, c13650, in13650_1, in13650_2, s12295[0]);
    wire[0:0] s13651, in13651_1, in13651_2;
    wire c13651;
    assign in13651_1 = {c12293};
    assign in13651_2 = {c12294};
    Full_Adder FA_13651(s13651, c13651, in13651_1, in13651_2, c12292);
    wire[0:0] s13652, in13652_1, in13652_2;
    wire c13652;
    assign in13652_1 = {c12296};
    assign in13652_2 = {c12297};
    Full_Adder FA_13652(s13652, c13652, in13652_1, in13652_2, c12295);
    wire[0:0] s13653, in13653_1, in13653_2;
    wire c13653;
    assign in13653_1 = {s12299[0]};
    assign in13653_2 = {s12300[0]};
    Full_Adder FA_13653(s13653, c13653, in13653_1, in13653_2, s12298[0]);
    wire[0:0] s13654, in13654_1, in13654_2;
    wire c13654;
    assign in13654_1 = {s12302[0]};
    assign in13654_2 = {s12303[0]};
    Full_Adder FA_13654(s13654, c13654, in13654_1, in13654_2, s12301[0]);
    wire[0:0] s13655, in13655_1, in13655_2;
    wire c13655;
    assign in13655_1 = {c12299};
    assign in13655_2 = {c12300};
    Full_Adder FA_13655(s13655, c13655, in13655_1, in13655_2, c12298);
    wire[0:0] s13656, in13656_1, in13656_2;
    wire c13656;
    assign in13656_1 = {c12302};
    assign in13656_2 = {c12303};
    Full_Adder FA_13656(s13656, c13656, in13656_1, in13656_2, c12301);
    wire[0:0] s13657, in13657_1, in13657_2;
    wire c13657;
    assign in13657_1 = {s12305[0]};
    assign in13657_2 = {s12306[0]};
    Full_Adder FA_13657(s13657, c13657, in13657_1, in13657_2, s12304[0]);
    wire[0:0] s13658, in13658_1, in13658_2;
    wire c13658;
    assign in13658_1 = {s12308[0]};
    assign in13658_2 = {s12309[0]};
    Full_Adder FA_13658(s13658, c13658, in13658_1, in13658_2, s12307[0]);
    wire[0:0] s13659, in13659_1, in13659_2;
    wire c13659;
    assign in13659_1 = {c12305};
    assign in13659_2 = {c12306};
    Full_Adder FA_13659(s13659, c13659, in13659_1, in13659_2, c12304);
    wire[0:0] s13660, in13660_1, in13660_2;
    wire c13660;
    assign in13660_1 = {c12308};
    assign in13660_2 = {c12309};
    Full_Adder FA_13660(s13660, c13660, in13660_1, in13660_2, c12307);
    wire[0:0] s13661, in13661_1, in13661_2;
    wire c13661;
    assign in13661_1 = {s12311[0]};
    assign in13661_2 = {s12312[0]};
    Full_Adder FA_13661(s13661, c13661, in13661_1, in13661_2, s12310[0]);
    wire[0:0] s13662, in13662_1, in13662_2;
    wire c13662;
    assign in13662_1 = {s12314[0]};
    assign in13662_2 = {s12315[0]};
    Full_Adder FA_13662(s13662, c13662, in13662_1, in13662_2, s12313[0]);
    wire[0:0] s13663, in13663_1, in13663_2;
    wire c13663;
    assign in13663_1 = {c12311};
    assign in13663_2 = {c12312};
    Full_Adder FA_13663(s13663, c13663, in13663_1, in13663_2, c12310);
    wire[0:0] s13664, in13664_1, in13664_2;
    wire c13664;
    assign in13664_1 = {c12314};
    assign in13664_2 = {c12315};
    Full_Adder FA_13664(s13664, c13664, in13664_1, in13664_2, c12313);
    wire[0:0] s13665, in13665_1, in13665_2;
    wire c13665;
    assign in13665_1 = {s12317[0]};
    assign in13665_2 = {s12318[0]};
    Full_Adder FA_13665(s13665, c13665, in13665_1, in13665_2, s12316[0]);
    wire[0:0] s13666, in13666_1, in13666_2;
    wire c13666;
    assign in13666_1 = {s12320[0]};
    assign in13666_2 = {s12321[0]};
    Full_Adder FA_13666(s13666, c13666, in13666_1, in13666_2, s12319[0]);
    wire[0:0] s13667, in13667_1, in13667_2;
    wire c13667;
    assign in13667_1 = {c12317};
    assign in13667_2 = {c12318};
    Full_Adder FA_13667(s13667, c13667, in13667_1, in13667_2, c12316);
    wire[0:0] s13668, in13668_1, in13668_2;
    wire c13668;
    assign in13668_1 = {c12320};
    assign in13668_2 = {c12321};
    Full_Adder FA_13668(s13668, c13668, in13668_1, in13668_2, c12319);
    wire[0:0] s13669, in13669_1, in13669_2;
    wire c13669;
    assign in13669_1 = {s12323[0]};
    assign in13669_2 = {s12324[0]};
    Full_Adder FA_13669(s13669, c13669, in13669_1, in13669_2, s12322[0]);
    wire[0:0] s13670, in13670_1, in13670_2;
    wire c13670;
    assign in13670_1 = {s12326[0]};
    assign in13670_2 = {s12327[0]};
    Full_Adder FA_13670(s13670, c13670, in13670_1, in13670_2, s12325[0]);
    wire[0:0] s13671, in13671_1, in13671_2;
    wire c13671;
    assign in13671_1 = {c12323};
    assign in13671_2 = {c12324};
    Full_Adder FA_13671(s13671, c13671, in13671_1, in13671_2, c12322);
    wire[0:0] s13672, in13672_1, in13672_2;
    wire c13672;
    assign in13672_1 = {c12326};
    assign in13672_2 = {c12327};
    Full_Adder FA_13672(s13672, c13672, in13672_1, in13672_2, c12325);
    wire[0:0] s13673, in13673_1, in13673_2;
    wire c13673;
    assign in13673_1 = {s12329[0]};
    assign in13673_2 = {s12330[0]};
    Full_Adder FA_13673(s13673, c13673, in13673_1, in13673_2, s12328[0]);
    wire[0:0] s13674, in13674_1, in13674_2;
    wire c13674;
    assign in13674_1 = {s12332[0]};
    assign in13674_2 = {s12333[0]};
    Full_Adder FA_13674(s13674, c13674, in13674_1, in13674_2, s12331[0]);
    wire[0:0] s13675, in13675_1, in13675_2;
    wire c13675;
    assign in13675_1 = {c12329};
    assign in13675_2 = {c12330};
    Full_Adder FA_13675(s13675, c13675, in13675_1, in13675_2, c12328);
    wire[0:0] s13676, in13676_1, in13676_2;
    wire c13676;
    assign in13676_1 = {c12332};
    assign in13676_2 = {c12333};
    Full_Adder FA_13676(s13676, c13676, in13676_1, in13676_2, c12331);
    wire[0:0] s13677, in13677_1, in13677_2;
    wire c13677;
    assign in13677_1 = {s12335[0]};
    assign in13677_2 = {s12336[0]};
    Full_Adder FA_13677(s13677, c13677, in13677_1, in13677_2, s12334[0]);
    wire[0:0] s13678, in13678_1, in13678_2;
    wire c13678;
    assign in13678_1 = {s12338[0]};
    assign in13678_2 = {s12339[0]};
    Full_Adder FA_13678(s13678, c13678, in13678_1, in13678_2, s12337[0]);
    wire[0:0] s13679, in13679_1, in13679_2;
    wire c13679;
    assign in13679_1 = {c12335};
    assign in13679_2 = {c12336};
    Full_Adder FA_13679(s13679, c13679, in13679_1, in13679_2, c12334);
    wire[0:0] s13680, in13680_1, in13680_2;
    wire c13680;
    assign in13680_1 = {c12338};
    assign in13680_2 = {c12339};
    Full_Adder FA_13680(s13680, c13680, in13680_1, in13680_2, c12337);
    wire[0:0] s13681, in13681_1, in13681_2;
    wire c13681;
    assign in13681_1 = {s12341[0]};
    assign in13681_2 = {s12342[0]};
    Full_Adder FA_13681(s13681, c13681, in13681_1, in13681_2, s12340[0]);
    wire[0:0] s13682, in13682_1, in13682_2;
    wire c13682;
    assign in13682_1 = {s12344[0]};
    assign in13682_2 = {s12345[0]};
    Full_Adder FA_13682(s13682, c13682, in13682_1, in13682_2, s12343[0]);
    wire[0:0] s13683, in13683_1, in13683_2;
    wire c13683;
    assign in13683_1 = {c12341};
    assign in13683_2 = {c12342};
    Full_Adder FA_13683(s13683, c13683, in13683_1, in13683_2, c12340);
    wire[0:0] s13684, in13684_1, in13684_2;
    wire c13684;
    assign in13684_1 = {c12344};
    assign in13684_2 = {c12345};
    Full_Adder FA_13684(s13684, c13684, in13684_1, in13684_2, c12343);
    wire[0:0] s13685, in13685_1, in13685_2;
    wire c13685;
    assign in13685_1 = {s12347[0]};
    assign in13685_2 = {s12348[0]};
    Full_Adder FA_13685(s13685, c13685, in13685_1, in13685_2, s12346[0]);
    wire[0:0] s13686, in13686_1, in13686_2;
    wire c13686;
    assign in13686_1 = {s12350[0]};
    assign in13686_2 = {s12351[0]};
    Full_Adder FA_13686(s13686, c13686, in13686_1, in13686_2, s12349[0]);
    wire[0:0] s13687, in13687_1, in13687_2;
    wire c13687;
    assign in13687_1 = {c12347};
    assign in13687_2 = {c12348};
    Full_Adder FA_13687(s13687, c13687, in13687_1, in13687_2, c12346);
    wire[0:0] s13688, in13688_1, in13688_2;
    wire c13688;
    assign in13688_1 = {c12350};
    assign in13688_2 = {c12351};
    Full_Adder FA_13688(s13688, c13688, in13688_1, in13688_2, c12349);
    wire[0:0] s13689, in13689_1, in13689_2;
    wire c13689;
    assign in13689_1 = {s12353[0]};
    assign in13689_2 = {s12354[0]};
    Full_Adder FA_13689(s13689, c13689, in13689_1, in13689_2, s12352[0]);
    wire[0:0] s13690, in13690_1, in13690_2;
    wire c13690;
    assign in13690_1 = {s12356[0]};
    assign in13690_2 = {s12357[0]};
    Full_Adder FA_13690(s13690, c13690, in13690_1, in13690_2, s12355[0]);
    wire[0:0] s13691, in13691_1, in13691_2;
    wire c13691;
    assign in13691_1 = {c12353};
    assign in13691_2 = {c12354};
    Full_Adder FA_13691(s13691, c13691, in13691_1, in13691_2, c12352);
    wire[0:0] s13692, in13692_1, in13692_2;
    wire c13692;
    assign in13692_1 = {c12356};
    assign in13692_2 = {c12357};
    Full_Adder FA_13692(s13692, c13692, in13692_1, in13692_2, c12355);
    wire[0:0] s13693, in13693_1, in13693_2;
    wire c13693;
    assign in13693_1 = {s12359[0]};
    assign in13693_2 = {s12360[0]};
    Full_Adder FA_13693(s13693, c13693, in13693_1, in13693_2, s12358[0]);
    wire[0:0] s13694, in13694_1, in13694_2;
    wire c13694;
    assign in13694_1 = {s12362[0]};
    assign in13694_2 = {s12363[0]};
    Full_Adder FA_13694(s13694, c13694, in13694_1, in13694_2, s12361[0]);
    wire[0:0] s13695, in13695_1, in13695_2;
    wire c13695;
    assign in13695_1 = {c12359};
    assign in13695_2 = {c12360};
    Full_Adder FA_13695(s13695, c13695, in13695_1, in13695_2, c12358);
    wire[0:0] s13696, in13696_1, in13696_2;
    wire c13696;
    assign in13696_1 = {c12362};
    assign in13696_2 = {c12363};
    Full_Adder FA_13696(s13696, c13696, in13696_1, in13696_2, c12361);
    wire[0:0] s13697, in13697_1, in13697_2;
    wire c13697;
    assign in13697_1 = {s12365[0]};
    assign in13697_2 = {s12366[0]};
    Full_Adder FA_13697(s13697, c13697, in13697_1, in13697_2, s12364[0]);
    wire[0:0] s13698, in13698_1, in13698_2;
    wire c13698;
    assign in13698_1 = {s12368[0]};
    assign in13698_2 = {s12369[0]};
    Full_Adder FA_13698(s13698, c13698, in13698_1, in13698_2, s12367[0]);
    wire[0:0] s13699, in13699_1, in13699_2;
    wire c13699;
    assign in13699_1 = {c12365};
    assign in13699_2 = {c12366};
    Full_Adder FA_13699(s13699, c13699, in13699_1, in13699_2, c12364);
    wire[0:0] s13700, in13700_1, in13700_2;
    wire c13700;
    assign in13700_1 = {c12368};
    assign in13700_2 = {c12369};
    Full_Adder FA_13700(s13700, c13700, in13700_1, in13700_2, c12367);
    wire[0:0] s13701, in13701_1, in13701_2;
    wire c13701;
    assign in13701_1 = {s12371[0]};
    assign in13701_2 = {s12372[0]};
    Full_Adder FA_13701(s13701, c13701, in13701_1, in13701_2, s12370[0]);
    wire[0:0] s13702, in13702_1, in13702_2;
    wire c13702;
    assign in13702_1 = {s12374[0]};
    assign in13702_2 = {s12375[0]};
    Full_Adder FA_13702(s13702, c13702, in13702_1, in13702_2, s12373[0]);
    wire[0:0] s13703, in13703_1, in13703_2;
    wire c13703;
    assign in13703_1 = {c12371};
    assign in13703_2 = {c12372};
    Full_Adder FA_13703(s13703, c13703, in13703_1, in13703_2, c12370);
    wire[0:0] s13704, in13704_1, in13704_2;
    wire c13704;
    assign in13704_1 = {c12374};
    assign in13704_2 = {c12375};
    Full_Adder FA_13704(s13704, c13704, in13704_1, in13704_2, c12373);
    wire[0:0] s13705, in13705_1, in13705_2;
    wire c13705;
    assign in13705_1 = {s12377[0]};
    assign in13705_2 = {s12378[0]};
    Full_Adder FA_13705(s13705, c13705, in13705_1, in13705_2, s12376[0]);
    wire[0:0] s13706, in13706_1, in13706_2;
    wire c13706;
    assign in13706_1 = {s12380[0]};
    assign in13706_2 = {s12381[0]};
    Full_Adder FA_13706(s13706, c13706, in13706_1, in13706_2, s12379[0]);
    wire[0:0] s13707, in13707_1, in13707_2;
    wire c13707;
    assign in13707_1 = {c12377};
    assign in13707_2 = {c12378};
    Full_Adder FA_13707(s13707, c13707, in13707_1, in13707_2, c12376);
    wire[0:0] s13708, in13708_1, in13708_2;
    wire c13708;
    assign in13708_1 = {c12380};
    assign in13708_2 = {c12381};
    Full_Adder FA_13708(s13708, c13708, in13708_1, in13708_2, c12379);
    wire[0:0] s13709, in13709_1, in13709_2;
    wire c13709;
    assign in13709_1 = {s12383[0]};
    assign in13709_2 = {s12384[0]};
    Full_Adder FA_13709(s13709, c13709, in13709_1, in13709_2, s12382[0]);
    wire[0:0] s13710, in13710_1, in13710_2;
    wire c13710;
    assign in13710_1 = {s12386[0]};
    assign in13710_2 = {s12387[0]};
    Full_Adder FA_13710(s13710, c13710, in13710_1, in13710_2, s12385[0]);
    wire[0:0] s13711, in13711_1, in13711_2;
    wire c13711;
    assign in13711_1 = {c12383};
    assign in13711_2 = {c12384};
    Full_Adder FA_13711(s13711, c13711, in13711_1, in13711_2, c12382);
    wire[0:0] s13712, in13712_1, in13712_2;
    wire c13712;
    assign in13712_1 = {c12386};
    assign in13712_2 = {c12387};
    Full_Adder FA_13712(s13712, c13712, in13712_1, in13712_2, c12385);
    wire[0:0] s13713, in13713_1, in13713_2;
    wire c13713;
    assign in13713_1 = {s12389[0]};
    assign in13713_2 = {s12390[0]};
    Full_Adder FA_13713(s13713, c13713, in13713_1, in13713_2, s12388[0]);
    wire[0:0] s13714, in13714_1, in13714_2;
    wire c13714;
    assign in13714_1 = {s12392[0]};
    assign in13714_2 = {s12393[0]};
    Full_Adder FA_13714(s13714, c13714, in13714_1, in13714_2, s12391[0]);
    wire[0:0] s13715, in13715_1, in13715_2;
    wire c13715;
    assign in13715_1 = {c12389};
    assign in13715_2 = {c12390};
    Full_Adder FA_13715(s13715, c13715, in13715_1, in13715_2, c12388);
    wire[0:0] s13716, in13716_1, in13716_2;
    wire c13716;
    assign in13716_1 = {c12392};
    assign in13716_2 = {c12393};
    Full_Adder FA_13716(s13716, c13716, in13716_1, in13716_2, c12391);
    wire[0:0] s13717, in13717_1, in13717_2;
    wire c13717;
    assign in13717_1 = {s12395[0]};
    assign in13717_2 = {s12396[0]};
    Full_Adder FA_13717(s13717, c13717, in13717_1, in13717_2, s12394[0]);
    wire[0:0] s13718, in13718_1, in13718_2;
    wire c13718;
    assign in13718_1 = {s12398[0]};
    assign in13718_2 = {s12399[0]};
    Full_Adder FA_13718(s13718, c13718, in13718_1, in13718_2, s12397[0]);
    wire[0:0] s13719, in13719_1, in13719_2;
    wire c13719;
    assign in13719_1 = {c12395};
    assign in13719_2 = {c12396};
    Full_Adder FA_13719(s13719, c13719, in13719_1, in13719_2, c12394);
    wire[0:0] s13720, in13720_1, in13720_2;
    wire c13720;
    assign in13720_1 = {c12398};
    assign in13720_2 = {c12399};
    Full_Adder FA_13720(s13720, c13720, in13720_1, in13720_2, c12397);
    wire[0:0] s13721, in13721_1, in13721_2;
    wire c13721;
    assign in13721_1 = {s12401[0]};
    assign in13721_2 = {s12402[0]};
    Full_Adder FA_13721(s13721, c13721, in13721_1, in13721_2, s12400[0]);
    wire[0:0] s13722, in13722_1, in13722_2;
    wire c13722;
    assign in13722_1 = {s12404[0]};
    assign in13722_2 = {s12405[0]};
    Full_Adder FA_13722(s13722, c13722, in13722_1, in13722_2, s12403[0]);
    wire[0:0] s13723, in13723_1, in13723_2;
    wire c13723;
    assign in13723_1 = {c12401};
    assign in13723_2 = {c12402};
    Full_Adder FA_13723(s13723, c13723, in13723_1, in13723_2, c12400);
    wire[0:0] s13724, in13724_1, in13724_2;
    wire c13724;
    assign in13724_1 = {c12404};
    assign in13724_2 = {c12405};
    Full_Adder FA_13724(s13724, c13724, in13724_1, in13724_2, c12403);
    wire[0:0] s13725, in13725_1, in13725_2;
    wire c13725;
    assign in13725_1 = {s12407[0]};
    assign in13725_2 = {s12408[0]};
    Full_Adder FA_13725(s13725, c13725, in13725_1, in13725_2, s12406[0]);
    wire[0:0] s13726, in13726_1, in13726_2;
    wire c13726;
    assign in13726_1 = {s12410[0]};
    assign in13726_2 = {s12411[0]};
    Full_Adder FA_13726(s13726, c13726, in13726_1, in13726_2, s12409[0]);
    wire[0:0] s13727, in13727_1, in13727_2;
    wire c13727;
    assign in13727_1 = {c12407};
    assign in13727_2 = {c12408};
    Full_Adder FA_13727(s13727, c13727, in13727_1, in13727_2, c12406);
    wire[0:0] s13728, in13728_1, in13728_2;
    wire c13728;
    assign in13728_1 = {c12410};
    assign in13728_2 = {c12411};
    Full_Adder FA_13728(s13728, c13728, in13728_1, in13728_2, c12409);
    wire[0:0] s13729, in13729_1, in13729_2;
    wire c13729;
    assign in13729_1 = {s12413[0]};
    assign in13729_2 = {s12414[0]};
    Full_Adder FA_13729(s13729, c13729, in13729_1, in13729_2, s12412[0]);
    wire[0:0] s13730, in13730_1, in13730_2;
    wire c13730;
    assign in13730_1 = {s12416[0]};
    assign in13730_2 = {s12417[0]};
    Full_Adder FA_13730(s13730, c13730, in13730_1, in13730_2, s12415[0]);
    wire[0:0] s13731, in13731_1, in13731_2;
    wire c13731;
    assign in13731_1 = {c12413};
    assign in13731_2 = {c12414};
    Full_Adder FA_13731(s13731, c13731, in13731_1, in13731_2, c12412);
    wire[0:0] s13732, in13732_1, in13732_2;
    wire c13732;
    assign in13732_1 = {c12416};
    assign in13732_2 = {c12417};
    Full_Adder FA_13732(s13732, c13732, in13732_1, in13732_2, c12415);
    wire[0:0] s13733, in13733_1, in13733_2;
    wire c13733;
    assign in13733_1 = {s12419[0]};
    assign in13733_2 = {s12420[0]};
    Full_Adder FA_13733(s13733, c13733, in13733_1, in13733_2, s12418[0]);
    wire[0:0] s13734, in13734_1, in13734_2;
    wire c13734;
    assign in13734_1 = {s12422[0]};
    assign in13734_2 = {s12423[0]};
    Full_Adder FA_13734(s13734, c13734, in13734_1, in13734_2, s12421[0]);
    wire[0:0] s13735, in13735_1, in13735_2;
    wire c13735;
    assign in13735_1 = {c12419};
    assign in13735_2 = {c12420};
    Full_Adder FA_13735(s13735, c13735, in13735_1, in13735_2, c12418);
    wire[0:0] s13736, in13736_1, in13736_2;
    wire c13736;
    assign in13736_1 = {c12422};
    assign in13736_2 = {c12423};
    Full_Adder FA_13736(s13736, c13736, in13736_1, in13736_2, c12421);
    wire[0:0] s13737, in13737_1, in13737_2;
    wire c13737;
    assign in13737_1 = {s12425[0]};
    assign in13737_2 = {s12426[0]};
    Full_Adder FA_13737(s13737, c13737, in13737_1, in13737_2, s12424[0]);
    wire[0:0] s13738, in13738_1, in13738_2;
    wire c13738;
    assign in13738_1 = {s12428[0]};
    assign in13738_2 = {s12429[0]};
    Full_Adder FA_13738(s13738, c13738, in13738_1, in13738_2, s12427[0]);
    wire[0:0] s13739, in13739_1, in13739_2;
    wire c13739;
    assign in13739_1 = {c12425};
    assign in13739_2 = {c12426};
    Full_Adder FA_13739(s13739, c13739, in13739_1, in13739_2, c12424);
    wire[0:0] s13740, in13740_1, in13740_2;
    wire c13740;
    assign in13740_1 = {c12428};
    assign in13740_2 = {c12429};
    Full_Adder FA_13740(s13740, c13740, in13740_1, in13740_2, c12427);
    wire[0:0] s13741, in13741_1, in13741_2;
    wire c13741;
    assign in13741_1 = {s12431[0]};
    assign in13741_2 = {s12432[0]};
    Full_Adder FA_13741(s13741, c13741, in13741_1, in13741_2, s12430[0]);
    wire[0:0] s13742, in13742_1, in13742_2;
    wire c13742;
    assign in13742_1 = {s12434[0]};
    assign in13742_2 = {s12435[0]};
    Full_Adder FA_13742(s13742, c13742, in13742_1, in13742_2, s12433[0]);
    wire[0:0] s13743, in13743_1, in13743_2;
    wire c13743;
    assign in13743_1 = {c12431};
    assign in13743_2 = {c12432};
    Full_Adder FA_13743(s13743, c13743, in13743_1, in13743_2, c12430);
    wire[0:0] s13744, in13744_1, in13744_2;
    wire c13744;
    assign in13744_1 = {c12434};
    assign in13744_2 = {c12435};
    Full_Adder FA_13744(s13744, c13744, in13744_1, in13744_2, c12433);
    wire[0:0] s13745, in13745_1, in13745_2;
    wire c13745;
    assign in13745_1 = {s12437[0]};
    assign in13745_2 = {s12438[0]};
    Full_Adder FA_13745(s13745, c13745, in13745_1, in13745_2, s12436[0]);
    wire[0:0] s13746, in13746_1, in13746_2;
    wire c13746;
    assign in13746_1 = {s12440[0]};
    assign in13746_2 = {s12441[0]};
    Full_Adder FA_13746(s13746, c13746, in13746_1, in13746_2, s12439[0]);
    wire[0:0] s13747, in13747_1, in13747_2;
    wire c13747;
    assign in13747_1 = {c12437};
    assign in13747_2 = {c12438};
    Full_Adder FA_13747(s13747, c13747, in13747_1, in13747_2, c12436);
    wire[0:0] s13748, in13748_1, in13748_2;
    wire c13748;
    assign in13748_1 = {c12440};
    assign in13748_2 = {c12441};
    Full_Adder FA_13748(s13748, c13748, in13748_1, in13748_2, c12439);
    wire[0:0] s13749, in13749_1, in13749_2;
    wire c13749;
    assign in13749_1 = {s12443[0]};
    assign in13749_2 = {s12444[0]};
    Full_Adder FA_13749(s13749, c13749, in13749_1, in13749_2, s12442[0]);
    wire[0:0] s13750, in13750_1, in13750_2;
    wire c13750;
    assign in13750_1 = {s12446[0]};
    assign in13750_2 = {s12447[0]};
    Full_Adder FA_13750(s13750, c13750, in13750_1, in13750_2, s12445[0]);
    wire[0:0] s13751, in13751_1, in13751_2;
    wire c13751;
    assign in13751_1 = {c12443};
    assign in13751_2 = {c12444};
    Full_Adder FA_13751(s13751, c13751, in13751_1, in13751_2, c12442);
    wire[0:0] s13752, in13752_1, in13752_2;
    wire c13752;
    assign in13752_1 = {c12446};
    assign in13752_2 = {c12447};
    Full_Adder FA_13752(s13752, c13752, in13752_1, in13752_2, c12445);
    wire[0:0] s13753, in13753_1, in13753_2;
    wire c13753;
    assign in13753_1 = {s12449[0]};
    assign in13753_2 = {s12450[0]};
    Full_Adder FA_13753(s13753, c13753, in13753_1, in13753_2, s12448[0]);
    wire[0:0] s13754, in13754_1, in13754_2;
    wire c13754;
    assign in13754_1 = {s12452[0]};
    assign in13754_2 = {s12453[0]};
    Full_Adder FA_13754(s13754, c13754, in13754_1, in13754_2, s12451[0]);
    wire[0:0] s13755, in13755_1, in13755_2;
    wire c13755;
    assign in13755_1 = {c12449};
    assign in13755_2 = {c12450};
    Full_Adder FA_13755(s13755, c13755, in13755_1, in13755_2, c12448);
    wire[0:0] s13756, in13756_1, in13756_2;
    wire c13756;
    assign in13756_1 = {c12452};
    assign in13756_2 = {c12453};
    Full_Adder FA_13756(s13756, c13756, in13756_1, in13756_2, c12451);
    wire[0:0] s13757, in13757_1, in13757_2;
    wire c13757;
    assign in13757_1 = {s12455[0]};
    assign in13757_2 = {s12456[0]};
    Full_Adder FA_13757(s13757, c13757, in13757_1, in13757_2, s12454[0]);
    wire[0:0] s13758, in13758_1, in13758_2;
    wire c13758;
    assign in13758_1 = {s12458[0]};
    assign in13758_2 = {s12459[0]};
    Full_Adder FA_13758(s13758, c13758, in13758_1, in13758_2, s12457[0]);
    wire[0:0] s13759, in13759_1, in13759_2;
    wire c13759;
    assign in13759_1 = {c12455};
    assign in13759_2 = {c12456};
    Full_Adder FA_13759(s13759, c13759, in13759_1, in13759_2, c12454);
    wire[0:0] s13760, in13760_1, in13760_2;
    wire c13760;
    assign in13760_1 = {c12458};
    assign in13760_2 = {c12459};
    Full_Adder FA_13760(s13760, c13760, in13760_1, in13760_2, c12457);
    wire[0:0] s13761, in13761_1, in13761_2;
    wire c13761;
    assign in13761_1 = {s12461[0]};
    assign in13761_2 = {s12462[0]};
    Full_Adder FA_13761(s13761, c13761, in13761_1, in13761_2, s12460[0]);
    wire[0:0] s13762, in13762_1, in13762_2;
    wire c13762;
    assign in13762_1 = {s12464[0]};
    assign in13762_2 = {s12465[0]};
    Full_Adder FA_13762(s13762, c13762, in13762_1, in13762_2, s12463[0]);
    wire[0:0] s13763, in13763_1, in13763_2;
    wire c13763;
    assign in13763_1 = {c12461};
    assign in13763_2 = {c12462};
    Full_Adder FA_13763(s13763, c13763, in13763_1, in13763_2, c12460);
    wire[0:0] s13764, in13764_1, in13764_2;
    wire c13764;
    assign in13764_1 = {c12464};
    assign in13764_2 = {c12465};
    Full_Adder FA_13764(s13764, c13764, in13764_1, in13764_2, c12463);
    wire[0:0] s13765, in13765_1, in13765_2;
    wire c13765;
    assign in13765_1 = {s12467[0]};
    assign in13765_2 = {s12468[0]};
    Full_Adder FA_13765(s13765, c13765, in13765_1, in13765_2, s12466[0]);
    wire[0:0] s13766, in13766_1, in13766_2;
    wire c13766;
    assign in13766_1 = {s12470[0]};
    assign in13766_2 = {s12471[0]};
    Full_Adder FA_13766(s13766, c13766, in13766_1, in13766_2, s12469[0]);
    wire[0:0] s13767, in13767_1, in13767_2;
    wire c13767;
    assign in13767_1 = {c12467};
    assign in13767_2 = {c12468};
    Full_Adder FA_13767(s13767, c13767, in13767_1, in13767_2, c12466);
    wire[0:0] s13768, in13768_1, in13768_2;
    wire c13768;
    assign in13768_1 = {c12470};
    assign in13768_2 = {c12471};
    Full_Adder FA_13768(s13768, c13768, in13768_1, in13768_2, c12469);
    wire[0:0] s13769, in13769_1, in13769_2;
    wire c13769;
    assign in13769_1 = {s12473[0]};
    assign in13769_2 = {s12474[0]};
    Full_Adder FA_13769(s13769, c13769, in13769_1, in13769_2, s12472[0]);
    wire[0:0] s13770, in13770_1, in13770_2;
    wire c13770;
    assign in13770_1 = {s12476[0]};
    assign in13770_2 = {s12477[0]};
    Full_Adder FA_13770(s13770, c13770, in13770_1, in13770_2, s12475[0]);
    wire[0:0] s13771, in13771_1, in13771_2;
    wire c13771;
    assign in13771_1 = {c12473};
    assign in13771_2 = {c12474};
    Full_Adder FA_13771(s13771, c13771, in13771_1, in13771_2, c12472);
    wire[0:0] s13772, in13772_1, in13772_2;
    wire c13772;
    assign in13772_1 = {c12476};
    assign in13772_2 = {c12477};
    Full_Adder FA_13772(s13772, c13772, in13772_1, in13772_2, c12475);
    wire[0:0] s13773, in13773_1, in13773_2;
    wire c13773;
    assign in13773_1 = {s12479[0]};
    assign in13773_2 = {s12480[0]};
    Full_Adder FA_13773(s13773, c13773, in13773_1, in13773_2, s12478[0]);
    wire[0:0] s13774, in13774_1, in13774_2;
    wire c13774;
    assign in13774_1 = {s12482[0]};
    assign in13774_2 = {s12483[0]};
    Full_Adder FA_13774(s13774, c13774, in13774_1, in13774_2, s12481[0]);
    wire[0:0] s13775, in13775_1, in13775_2;
    wire c13775;
    assign in13775_1 = {c12479};
    assign in13775_2 = {c12480};
    Full_Adder FA_13775(s13775, c13775, in13775_1, in13775_2, c12478);
    wire[0:0] s13776, in13776_1, in13776_2;
    wire c13776;
    assign in13776_1 = {c12482};
    assign in13776_2 = {c12483};
    Full_Adder FA_13776(s13776, c13776, in13776_1, in13776_2, c12481);
    wire[0:0] s13777, in13777_1, in13777_2;
    wire c13777;
    assign in13777_1 = {s12485[0]};
    assign in13777_2 = {s12486[0]};
    Full_Adder FA_13777(s13777, c13777, in13777_1, in13777_2, s12484[0]);
    wire[0:0] s13778, in13778_1, in13778_2;
    wire c13778;
    assign in13778_1 = {s12488[0]};
    assign in13778_2 = {s12489[0]};
    Full_Adder FA_13778(s13778, c13778, in13778_1, in13778_2, s12487[0]);
    wire[0:0] s13779, in13779_1, in13779_2;
    wire c13779;
    assign in13779_1 = {c12485};
    assign in13779_2 = {c12486};
    Full_Adder FA_13779(s13779, c13779, in13779_1, in13779_2, c12484);
    wire[0:0] s13780, in13780_1, in13780_2;
    wire c13780;
    assign in13780_1 = {c12488};
    assign in13780_2 = {c12489};
    Full_Adder FA_13780(s13780, c13780, in13780_1, in13780_2, c12487);
    wire[0:0] s13781, in13781_1, in13781_2;
    wire c13781;
    assign in13781_1 = {s12491[0]};
    assign in13781_2 = {s12492[0]};
    Full_Adder FA_13781(s13781, c13781, in13781_1, in13781_2, s12490[0]);
    wire[0:0] s13782, in13782_1, in13782_2;
    wire c13782;
    assign in13782_1 = {s12494[0]};
    assign in13782_2 = {s12495[0]};
    Full_Adder FA_13782(s13782, c13782, in13782_1, in13782_2, s12493[0]);
    wire[0:0] s13783, in13783_1, in13783_2;
    wire c13783;
    assign in13783_1 = {c12491};
    assign in13783_2 = {c12492};
    Full_Adder FA_13783(s13783, c13783, in13783_1, in13783_2, c12490);
    wire[0:0] s13784, in13784_1, in13784_2;
    wire c13784;
    assign in13784_1 = {c12494};
    assign in13784_2 = {c12495};
    Full_Adder FA_13784(s13784, c13784, in13784_1, in13784_2, c12493);
    wire[0:0] s13785, in13785_1, in13785_2;
    wire c13785;
    assign in13785_1 = {s12497[0]};
    assign in13785_2 = {s12498[0]};
    Full_Adder FA_13785(s13785, c13785, in13785_1, in13785_2, s12496[0]);
    wire[0:0] s13786, in13786_1, in13786_2;
    wire c13786;
    assign in13786_1 = {s12500[0]};
    assign in13786_2 = {s12501[0]};
    Full_Adder FA_13786(s13786, c13786, in13786_1, in13786_2, s12499[0]);
    wire[0:0] s13787, in13787_1, in13787_2;
    wire c13787;
    assign in13787_1 = {c12497};
    assign in13787_2 = {c12498};
    Full_Adder FA_13787(s13787, c13787, in13787_1, in13787_2, c12496);
    wire[0:0] s13788, in13788_1, in13788_2;
    wire c13788;
    assign in13788_1 = {c12500};
    assign in13788_2 = {c12501};
    Full_Adder FA_13788(s13788, c13788, in13788_1, in13788_2, c12499);
    wire[0:0] s13789, in13789_1, in13789_2;
    wire c13789;
    assign in13789_1 = {s12503[0]};
    assign in13789_2 = {s12504[0]};
    Full_Adder FA_13789(s13789, c13789, in13789_1, in13789_2, s12502[0]);
    wire[0:0] s13790, in13790_1, in13790_2;
    wire c13790;
    assign in13790_1 = {s12506[0]};
    assign in13790_2 = {s12507[0]};
    Full_Adder FA_13790(s13790, c13790, in13790_1, in13790_2, s12505[0]);
    wire[0:0] s13791, in13791_1, in13791_2;
    wire c13791;
    assign in13791_1 = {c12503};
    assign in13791_2 = {c12504};
    Full_Adder FA_13791(s13791, c13791, in13791_1, in13791_2, c12502);
    wire[0:0] s13792, in13792_1, in13792_2;
    wire c13792;
    assign in13792_1 = {c12506};
    assign in13792_2 = {c12507};
    Full_Adder FA_13792(s13792, c13792, in13792_1, in13792_2, c12505);
    wire[0:0] s13793, in13793_1, in13793_2;
    wire c13793;
    assign in13793_1 = {s12509[0]};
    assign in13793_2 = {s12510[0]};
    Full_Adder FA_13793(s13793, c13793, in13793_1, in13793_2, s12508[0]);
    wire[0:0] s13794, in13794_1, in13794_2;
    wire c13794;
    assign in13794_1 = {s12512[0]};
    assign in13794_2 = {s12513[0]};
    Full_Adder FA_13794(s13794, c13794, in13794_1, in13794_2, s12511[0]);
    wire[0:0] s13795, in13795_1, in13795_2;
    wire c13795;
    assign in13795_1 = {c12509};
    assign in13795_2 = {c12510};
    Full_Adder FA_13795(s13795, c13795, in13795_1, in13795_2, c12508);
    wire[0:0] s13796, in13796_1, in13796_2;
    wire c13796;
    assign in13796_1 = {c12512};
    assign in13796_2 = {c12513};
    Full_Adder FA_13796(s13796, c13796, in13796_1, in13796_2, c12511);
    wire[0:0] s13797, in13797_1, in13797_2;
    wire c13797;
    assign in13797_1 = {s12515[0]};
    assign in13797_2 = {s12516[0]};
    Full_Adder FA_13797(s13797, c13797, in13797_1, in13797_2, s12514[0]);
    wire[0:0] s13798, in13798_1, in13798_2;
    wire c13798;
    assign in13798_1 = {s12518[0]};
    assign in13798_2 = {s12519[0]};
    Full_Adder FA_13798(s13798, c13798, in13798_1, in13798_2, s12517[0]);
    wire[0:0] s13799, in13799_1, in13799_2;
    wire c13799;
    assign in13799_1 = {c12515};
    assign in13799_2 = {c12516};
    Full_Adder FA_13799(s13799, c13799, in13799_1, in13799_2, c12514);
    wire[0:0] s13800, in13800_1, in13800_2;
    wire c13800;
    assign in13800_1 = {c12518};
    assign in13800_2 = {c12519};
    Full_Adder FA_13800(s13800, c13800, in13800_1, in13800_2, c12517);
    wire[0:0] s13801, in13801_1, in13801_2;
    wire c13801;
    assign in13801_1 = {s12521[0]};
    assign in13801_2 = {s12522[0]};
    Full_Adder FA_13801(s13801, c13801, in13801_1, in13801_2, s12520[0]);
    wire[0:0] s13802, in13802_1, in13802_2;
    wire c13802;
    assign in13802_1 = {s12524[0]};
    assign in13802_2 = {s12525[0]};
    Full_Adder FA_13802(s13802, c13802, in13802_1, in13802_2, s12523[0]);
    wire[0:0] s13803, in13803_1, in13803_2;
    wire c13803;
    assign in13803_1 = {c12521};
    assign in13803_2 = {c12522};
    Full_Adder FA_13803(s13803, c13803, in13803_1, in13803_2, c12520);
    wire[0:0] s13804, in13804_1, in13804_2;
    wire c13804;
    assign in13804_1 = {c12524};
    assign in13804_2 = {c12525};
    Full_Adder FA_13804(s13804, c13804, in13804_1, in13804_2, c12523);
    wire[0:0] s13805, in13805_1, in13805_2;
    wire c13805;
    assign in13805_1 = {s12527[0]};
    assign in13805_2 = {s12528[0]};
    Full_Adder FA_13805(s13805, c13805, in13805_1, in13805_2, s12526[0]);
    wire[0:0] s13806, in13806_1, in13806_2;
    wire c13806;
    assign in13806_1 = {s12530[0]};
    assign in13806_2 = {s12531[0]};
    Full_Adder FA_13806(s13806, c13806, in13806_1, in13806_2, s12529[0]);
    wire[0:0] s13807, in13807_1, in13807_2;
    wire c13807;
    assign in13807_1 = {c12527};
    assign in13807_2 = {c12528};
    Full_Adder FA_13807(s13807, c13807, in13807_1, in13807_2, c12526);
    wire[0:0] s13808, in13808_1, in13808_2;
    wire c13808;
    assign in13808_1 = {c12530};
    assign in13808_2 = {c12531};
    Full_Adder FA_13808(s13808, c13808, in13808_1, in13808_2, c12529);
    wire[0:0] s13809, in13809_1, in13809_2;
    wire c13809;
    assign in13809_1 = {s12533[0]};
    assign in13809_2 = {s12534[0]};
    Full_Adder FA_13809(s13809, c13809, in13809_1, in13809_2, s12532[0]);
    wire[0:0] s13810, in13810_1, in13810_2;
    wire c13810;
    assign in13810_1 = {s12536[0]};
    assign in13810_2 = {s12537[0]};
    Full_Adder FA_13810(s13810, c13810, in13810_1, in13810_2, s12535[0]);
    wire[0:0] s13811, in13811_1, in13811_2;
    wire c13811;
    assign in13811_1 = {c12533};
    assign in13811_2 = {c12534};
    Full_Adder FA_13811(s13811, c13811, in13811_1, in13811_2, c12532);
    wire[0:0] s13812, in13812_1, in13812_2;
    wire c13812;
    assign in13812_1 = {c12536};
    assign in13812_2 = {c12537};
    Full_Adder FA_13812(s13812, c13812, in13812_1, in13812_2, c12535);
    wire[0:0] s13813, in13813_1, in13813_2;
    wire c13813;
    assign in13813_1 = {s12539[0]};
    assign in13813_2 = {s12540[0]};
    Full_Adder FA_13813(s13813, c13813, in13813_1, in13813_2, s12538[0]);
    wire[0:0] s13814, in13814_1, in13814_2;
    wire c13814;
    assign in13814_1 = {s12542[0]};
    assign in13814_2 = {s12543[0]};
    Full_Adder FA_13814(s13814, c13814, in13814_1, in13814_2, s12541[0]);
    wire[0:0] s13815, in13815_1, in13815_2;
    wire c13815;
    assign in13815_1 = {c12539};
    assign in13815_2 = {c12540};
    Full_Adder FA_13815(s13815, c13815, in13815_1, in13815_2, c12538);
    wire[0:0] s13816, in13816_1, in13816_2;
    wire c13816;
    assign in13816_1 = {c12542};
    assign in13816_2 = {c12543};
    Full_Adder FA_13816(s13816, c13816, in13816_1, in13816_2, c12541);
    wire[0:0] s13817, in13817_1, in13817_2;
    wire c13817;
    assign in13817_1 = {s12545[0]};
    assign in13817_2 = {s12546[0]};
    Full_Adder FA_13817(s13817, c13817, in13817_1, in13817_2, s12544[0]);
    wire[0:0] s13818, in13818_1, in13818_2;
    wire c13818;
    assign in13818_1 = {s12548[0]};
    assign in13818_2 = {s12549[0]};
    Full_Adder FA_13818(s13818, c13818, in13818_1, in13818_2, s12547[0]);
    wire[0:0] s13819, in13819_1, in13819_2;
    wire c13819;
    assign in13819_1 = {c12545};
    assign in13819_2 = {c12546};
    Full_Adder FA_13819(s13819, c13819, in13819_1, in13819_2, c12544);
    wire[0:0] s13820, in13820_1, in13820_2;
    wire c13820;
    assign in13820_1 = {c12548};
    assign in13820_2 = {c12549};
    Full_Adder FA_13820(s13820, c13820, in13820_1, in13820_2, c12547);
    wire[0:0] s13821, in13821_1, in13821_2;
    wire c13821;
    assign in13821_1 = {s12551[0]};
    assign in13821_2 = {s12552[0]};
    Full_Adder FA_13821(s13821, c13821, in13821_1, in13821_2, s12550[0]);
    wire[0:0] s13822, in13822_1, in13822_2;
    wire c13822;
    assign in13822_1 = {s12554[0]};
    assign in13822_2 = {s12555[0]};
    Full_Adder FA_13822(s13822, c13822, in13822_1, in13822_2, s12553[0]);
    wire[0:0] s13823, in13823_1, in13823_2;
    wire c13823;
    assign in13823_1 = {c12551};
    assign in13823_2 = {c12552};
    Full_Adder FA_13823(s13823, c13823, in13823_1, in13823_2, c12550);
    wire[0:0] s13824, in13824_1, in13824_2;
    wire c13824;
    assign in13824_1 = {c12554};
    assign in13824_2 = {c12555};
    Full_Adder FA_13824(s13824, c13824, in13824_1, in13824_2, c12553);
    wire[0:0] s13825, in13825_1, in13825_2;
    wire c13825;
    assign in13825_1 = {s12557[0]};
    assign in13825_2 = {s12558[0]};
    Full_Adder FA_13825(s13825, c13825, in13825_1, in13825_2, s12556[0]);
    wire[0:0] s13826, in13826_1, in13826_2;
    wire c13826;
    assign in13826_1 = {s12560[0]};
    assign in13826_2 = {s12561[0]};
    Full_Adder FA_13826(s13826, c13826, in13826_1, in13826_2, s12559[0]);
    wire[0:0] s13827, in13827_1, in13827_2;
    wire c13827;
    assign in13827_1 = {c12557};
    assign in13827_2 = {c12558};
    Full_Adder FA_13827(s13827, c13827, in13827_1, in13827_2, c12556);
    wire[0:0] s13828, in13828_1, in13828_2;
    wire c13828;
    assign in13828_1 = {c12560};
    assign in13828_2 = {c12561};
    Full_Adder FA_13828(s13828, c13828, in13828_1, in13828_2, c12559);
    wire[0:0] s13829, in13829_1, in13829_2;
    wire c13829;
    assign in13829_1 = {s12563[0]};
    assign in13829_2 = {s12564[0]};
    Full_Adder FA_13829(s13829, c13829, in13829_1, in13829_2, s12562[0]);
    wire[0:0] s13830, in13830_1, in13830_2;
    wire c13830;
    assign in13830_1 = {s12566[0]};
    assign in13830_2 = {s12567[0]};
    Full_Adder FA_13830(s13830, c13830, in13830_1, in13830_2, s12565[0]);
    wire[0:0] s13831, in13831_1, in13831_2;
    wire c13831;
    assign in13831_1 = {c12563};
    assign in13831_2 = {c12564};
    Full_Adder FA_13831(s13831, c13831, in13831_1, in13831_2, c12562);
    wire[0:0] s13832, in13832_1, in13832_2;
    wire c13832;
    assign in13832_1 = {c12566};
    assign in13832_2 = {c12567};
    Full_Adder FA_13832(s13832, c13832, in13832_1, in13832_2, c12565);
    wire[0:0] s13833, in13833_1, in13833_2;
    wire c13833;
    assign in13833_1 = {s12569[0]};
    assign in13833_2 = {s12570[0]};
    Full_Adder FA_13833(s13833, c13833, in13833_1, in13833_2, s12568[0]);
    wire[0:0] s13834, in13834_1, in13834_2;
    wire c13834;
    assign in13834_1 = {s12572[0]};
    assign in13834_2 = {s12573[0]};
    Full_Adder FA_13834(s13834, c13834, in13834_1, in13834_2, s12571[0]);
    wire[0:0] s13835, in13835_1, in13835_2;
    wire c13835;
    assign in13835_1 = {c12569};
    assign in13835_2 = {c12570};
    Full_Adder FA_13835(s13835, c13835, in13835_1, in13835_2, c12568);
    wire[0:0] s13836, in13836_1, in13836_2;
    wire c13836;
    assign in13836_1 = {c12572};
    assign in13836_2 = {c12573};
    Full_Adder FA_13836(s13836, c13836, in13836_1, in13836_2, c12571);
    wire[0:0] s13837, in13837_1, in13837_2;
    wire c13837;
    assign in13837_1 = {s12575[0]};
    assign in13837_2 = {s12576[0]};
    Full_Adder FA_13837(s13837, c13837, in13837_1, in13837_2, s12574[0]);
    wire[0:0] s13838, in13838_1, in13838_2;
    wire c13838;
    assign in13838_1 = {s12578[0]};
    assign in13838_2 = {s12579[0]};
    Full_Adder FA_13838(s13838, c13838, in13838_1, in13838_2, s12577[0]);
    wire[0:0] s13839, in13839_1, in13839_2;
    wire c13839;
    assign in13839_1 = {c12575};
    assign in13839_2 = {c12576};
    Full_Adder FA_13839(s13839, c13839, in13839_1, in13839_2, c12574);
    wire[0:0] s13840, in13840_1, in13840_2;
    wire c13840;
    assign in13840_1 = {c12578};
    assign in13840_2 = {c12579};
    Full_Adder FA_13840(s13840, c13840, in13840_1, in13840_2, c12577);
    wire[0:0] s13841, in13841_1, in13841_2;
    wire c13841;
    assign in13841_1 = {s12581[0]};
    assign in13841_2 = {s12582[0]};
    Full_Adder FA_13841(s13841, c13841, in13841_1, in13841_2, s12580[0]);
    wire[0:0] s13842, in13842_1, in13842_2;
    wire c13842;
    assign in13842_1 = {s12584[0]};
    assign in13842_2 = {s12585[0]};
    Full_Adder FA_13842(s13842, c13842, in13842_1, in13842_2, s12583[0]);
    wire[0:0] s13843, in13843_1, in13843_2;
    wire c13843;
    assign in13843_1 = {c12581};
    assign in13843_2 = {c12582};
    Full_Adder FA_13843(s13843, c13843, in13843_1, in13843_2, c12580);
    wire[0:0] s13844, in13844_1, in13844_2;
    wire c13844;
    assign in13844_1 = {c12584};
    assign in13844_2 = {c12585};
    Full_Adder FA_13844(s13844, c13844, in13844_1, in13844_2, c12583);
    wire[0:0] s13845, in13845_1, in13845_2;
    wire c13845;
    assign in13845_1 = {s12587[0]};
    assign in13845_2 = {s12588[0]};
    Full_Adder FA_13845(s13845, c13845, in13845_1, in13845_2, s12586[0]);
    wire[0:0] s13846, in13846_1, in13846_2;
    wire c13846;
    assign in13846_1 = {s12590[0]};
    assign in13846_2 = {s12591[0]};
    Full_Adder FA_13846(s13846, c13846, in13846_1, in13846_2, s12589[0]);
    wire[0:0] s13847, in13847_1, in13847_2;
    wire c13847;
    assign in13847_1 = {c12587};
    assign in13847_2 = {c12588};
    Full_Adder FA_13847(s13847, c13847, in13847_1, in13847_2, c12586);
    wire[0:0] s13848, in13848_1, in13848_2;
    wire c13848;
    assign in13848_1 = {c12590};
    assign in13848_2 = {c12591};
    Full_Adder FA_13848(s13848, c13848, in13848_1, in13848_2, c12589);
    wire[0:0] s13849, in13849_1, in13849_2;
    wire c13849;
    assign in13849_1 = {s12593[0]};
    assign in13849_2 = {s12594[0]};
    Full_Adder FA_13849(s13849, c13849, in13849_1, in13849_2, s12592[0]);
    wire[0:0] s13850, in13850_1, in13850_2;
    wire c13850;
    assign in13850_1 = {s12596[0]};
    assign in13850_2 = {s12597[0]};
    Full_Adder FA_13850(s13850, c13850, in13850_1, in13850_2, s12595[0]);
    wire[0:0] s13851, in13851_1, in13851_2;
    wire c13851;
    assign in13851_1 = {c12593};
    assign in13851_2 = {c12594};
    Full_Adder FA_13851(s13851, c13851, in13851_1, in13851_2, c12592);
    wire[0:0] s13852, in13852_1, in13852_2;
    wire c13852;
    assign in13852_1 = {c12596};
    assign in13852_2 = {c12597};
    Full_Adder FA_13852(s13852, c13852, in13852_1, in13852_2, c12595);
    wire[0:0] s13853, in13853_1, in13853_2;
    wire c13853;
    assign in13853_1 = {s12599[0]};
    assign in13853_2 = {s12600[0]};
    Full_Adder FA_13853(s13853, c13853, in13853_1, in13853_2, s12598[0]);
    wire[0:0] s13854, in13854_1, in13854_2;
    wire c13854;
    assign in13854_1 = {s12602[0]};
    assign in13854_2 = {s12603[0]};
    Full_Adder FA_13854(s13854, c13854, in13854_1, in13854_2, s12601[0]);
    wire[0:0] s13855, in13855_1, in13855_2;
    wire c13855;
    assign in13855_1 = {c12599};
    assign in13855_2 = {c12600};
    Full_Adder FA_13855(s13855, c13855, in13855_1, in13855_2, c12598);
    wire[0:0] s13856, in13856_1, in13856_2;
    wire c13856;
    assign in13856_1 = {c12602};
    assign in13856_2 = {c12603};
    Full_Adder FA_13856(s13856, c13856, in13856_1, in13856_2, c12601);
    wire[0:0] s13857, in13857_1, in13857_2;
    wire c13857;
    assign in13857_1 = {s12605[0]};
    assign in13857_2 = {s12606[0]};
    Full_Adder FA_13857(s13857, c13857, in13857_1, in13857_2, s12604[0]);
    wire[0:0] s13858, in13858_1, in13858_2;
    wire c13858;
    assign in13858_1 = {s12608[0]};
    assign in13858_2 = {s12609[0]};
    Full_Adder FA_13858(s13858, c13858, in13858_1, in13858_2, s12607[0]);
    wire[0:0] s13859, in13859_1, in13859_2;
    wire c13859;
    assign in13859_1 = {c12605};
    assign in13859_2 = {c12606};
    Full_Adder FA_13859(s13859, c13859, in13859_1, in13859_2, c12604);
    wire[0:0] s13860, in13860_1, in13860_2;
    wire c13860;
    assign in13860_1 = {c12608};
    assign in13860_2 = {c12609};
    Full_Adder FA_13860(s13860, c13860, in13860_1, in13860_2, c12607);
    wire[0:0] s13861, in13861_1, in13861_2;
    wire c13861;
    assign in13861_1 = {s12611[0]};
    assign in13861_2 = {s12612[0]};
    Full_Adder FA_13861(s13861, c13861, in13861_1, in13861_2, s12610[0]);
    wire[0:0] s13862, in13862_1, in13862_2;
    wire c13862;
    assign in13862_1 = {s12614[0]};
    assign in13862_2 = {s12615[0]};
    Full_Adder FA_13862(s13862, c13862, in13862_1, in13862_2, s12613[0]);
    wire[0:0] s13863, in13863_1, in13863_2;
    wire c13863;
    assign in13863_1 = {c12611};
    assign in13863_2 = {c12612};
    Full_Adder FA_13863(s13863, c13863, in13863_1, in13863_2, c12610);
    wire[0:0] s13864, in13864_1, in13864_2;
    wire c13864;
    assign in13864_1 = {c12614};
    assign in13864_2 = {c12615};
    Full_Adder FA_13864(s13864, c13864, in13864_1, in13864_2, c12613);
    wire[0:0] s13865, in13865_1, in13865_2;
    wire c13865;
    assign in13865_1 = {s12617[0]};
    assign in13865_2 = {s12618[0]};
    Full_Adder FA_13865(s13865, c13865, in13865_1, in13865_2, s12616[0]);
    wire[0:0] s13866, in13866_1, in13866_2;
    wire c13866;
    assign in13866_1 = {s12620[0]};
    assign in13866_2 = {s12621[0]};
    Full_Adder FA_13866(s13866, c13866, in13866_1, in13866_2, s12619[0]);
    wire[0:0] s13867, in13867_1, in13867_2;
    wire c13867;
    assign in13867_1 = {c12617};
    assign in13867_2 = {c12618};
    Full_Adder FA_13867(s13867, c13867, in13867_1, in13867_2, c12616);
    wire[0:0] s13868, in13868_1, in13868_2;
    wire c13868;
    assign in13868_1 = {c12620};
    assign in13868_2 = {c12621};
    Full_Adder FA_13868(s13868, c13868, in13868_1, in13868_2, c12619);
    wire[0:0] s13869, in13869_1, in13869_2;
    wire c13869;
    assign in13869_1 = {s12623[0]};
    assign in13869_2 = {s12624[0]};
    Full_Adder FA_13869(s13869, c13869, in13869_1, in13869_2, s12622[0]);
    wire[0:0] s13870, in13870_1, in13870_2;
    wire c13870;
    assign in13870_1 = {s12626[0]};
    assign in13870_2 = {s12627[0]};
    Full_Adder FA_13870(s13870, c13870, in13870_1, in13870_2, s12625[0]);
    wire[0:0] s13871, in13871_1, in13871_2;
    wire c13871;
    assign in13871_1 = {c12623};
    assign in13871_2 = {c12624};
    Full_Adder FA_13871(s13871, c13871, in13871_1, in13871_2, c12622);
    wire[0:0] s13872, in13872_1, in13872_2;
    wire c13872;
    assign in13872_1 = {c12626};
    assign in13872_2 = {c12627};
    Full_Adder FA_13872(s13872, c13872, in13872_1, in13872_2, c12625);
    wire[0:0] s13873, in13873_1, in13873_2;
    wire c13873;
    assign in13873_1 = {s12629[0]};
    assign in13873_2 = {s12630[0]};
    Full_Adder FA_13873(s13873, c13873, in13873_1, in13873_2, s12628[0]);
    wire[0:0] s13874, in13874_1, in13874_2;
    wire c13874;
    assign in13874_1 = {s12632[0]};
    assign in13874_2 = {s12633[0]};
    Full_Adder FA_13874(s13874, c13874, in13874_1, in13874_2, s12631[0]);
    wire[0:0] s13875, in13875_1, in13875_2;
    wire c13875;
    assign in13875_1 = {c12629};
    assign in13875_2 = {c12630};
    Full_Adder FA_13875(s13875, c13875, in13875_1, in13875_2, c12628);
    wire[0:0] s13876, in13876_1, in13876_2;
    wire c13876;
    assign in13876_1 = {c12632};
    assign in13876_2 = {c12633};
    Full_Adder FA_13876(s13876, c13876, in13876_1, in13876_2, c12631);
    wire[0:0] s13877, in13877_1, in13877_2;
    wire c13877;
    assign in13877_1 = {s12635[0]};
    assign in13877_2 = {s12636[0]};
    Full_Adder FA_13877(s13877, c13877, in13877_1, in13877_2, s12634[0]);
    wire[0:0] s13878, in13878_1, in13878_2;
    wire c13878;
    assign in13878_1 = {s12638[0]};
    assign in13878_2 = {s12639[0]};
    Full_Adder FA_13878(s13878, c13878, in13878_1, in13878_2, s12637[0]);
    wire[0:0] s13879, in13879_1, in13879_2;
    wire c13879;
    assign in13879_1 = {c12635};
    assign in13879_2 = {c12636};
    Full_Adder FA_13879(s13879, c13879, in13879_1, in13879_2, c12634);
    wire[0:0] s13880, in13880_1, in13880_2;
    wire c13880;
    assign in13880_1 = {c12638};
    assign in13880_2 = {c12639};
    Full_Adder FA_13880(s13880, c13880, in13880_1, in13880_2, c12637);
    wire[0:0] s13881, in13881_1, in13881_2;
    wire c13881;
    assign in13881_1 = {s12641[0]};
    assign in13881_2 = {s12642[0]};
    Full_Adder FA_13881(s13881, c13881, in13881_1, in13881_2, s12640[0]);
    wire[0:0] s13882, in13882_1, in13882_2;
    wire c13882;
    assign in13882_1 = {s12644[0]};
    assign in13882_2 = {s12645[0]};
    Full_Adder FA_13882(s13882, c13882, in13882_1, in13882_2, s12643[0]);
    wire[0:0] s13883, in13883_1, in13883_2;
    wire c13883;
    assign in13883_1 = {c12641};
    assign in13883_2 = {c12642};
    Full_Adder FA_13883(s13883, c13883, in13883_1, in13883_2, c12640);
    wire[0:0] s13884, in13884_1, in13884_2;
    wire c13884;
    assign in13884_1 = {c12644};
    assign in13884_2 = {c12645};
    Full_Adder FA_13884(s13884, c13884, in13884_1, in13884_2, c12643);
    wire[0:0] s13885, in13885_1, in13885_2;
    wire c13885;
    assign in13885_1 = {s12647[0]};
    assign in13885_2 = {s12648[0]};
    Full_Adder FA_13885(s13885, c13885, in13885_1, in13885_2, s12646[0]);
    wire[0:0] s13886, in13886_1, in13886_2;
    wire c13886;
    assign in13886_1 = {s12650[0]};
    assign in13886_2 = {s12651[0]};
    Full_Adder FA_13886(s13886, c13886, in13886_1, in13886_2, s12649[0]);
    wire[0:0] s13887, in13887_1, in13887_2;
    wire c13887;
    assign in13887_1 = {c12647};
    assign in13887_2 = {c12648};
    Full_Adder FA_13887(s13887, c13887, in13887_1, in13887_2, c12646);
    wire[0:0] s13888, in13888_1, in13888_2;
    wire c13888;
    assign in13888_1 = {c12650};
    assign in13888_2 = {c12651};
    Full_Adder FA_13888(s13888, c13888, in13888_1, in13888_2, c12649);
    wire[0:0] s13889, in13889_1, in13889_2;
    wire c13889;
    assign in13889_1 = {s12653[0]};
    assign in13889_2 = {s12654[0]};
    Full_Adder FA_13889(s13889, c13889, in13889_1, in13889_2, s12652[0]);
    wire[0:0] s13890, in13890_1, in13890_2;
    wire c13890;
    assign in13890_1 = {s12656[0]};
    assign in13890_2 = {s12657[0]};
    Full_Adder FA_13890(s13890, c13890, in13890_1, in13890_2, s12655[0]);
    wire[0:0] s13891, in13891_1, in13891_2;
    wire c13891;
    assign in13891_1 = {c12653};
    assign in13891_2 = {c12654};
    Full_Adder FA_13891(s13891, c13891, in13891_1, in13891_2, c12652);
    wire[0:0] s13892, in13892_1, in13892_2;
    wire c13892;
    assign in13892_1 = {c12656};
    assign in13892_2 = {c12657};
    Full_Adder FA_13892(s13892, c13892, in13892_1, in13892_2, c12655);
    wire[0:0] s13893, in13893_1, in13893_2;
    wire c13893;
    assign in13893_1 = {s12659[0]};
    assign in13893_2 = {s12660[0]};
    Full_Adder FA_13893(s13893, c13893, in13893_1, in13893_2, s12658[0]);
    wire[0:0] s13894, in13894_1, in13894_2;
    wire c13894;
    assign in13894_1 = {s12662[0]};
    assign in13894_2 = {s12663[0]};
    Full_Adder FA_13894(s13894, c13894, in13894_1, in13894_2, s12661[0]);
    wire[0:0] s13895, in13895_1, in13895_2;
    wire c13895;
    assign in13895_1 = {c12659};
    assign in13895_2 = {c12660};
    Full_Adder FA_13895(s13895, c13895, in13895_1, in13895_2, c12658);
    wire[0:0] s13896, in13896_1, in13896_2;
    wire c13896;
    assign in13896_1 = {c12662};
    assign in13896_2 = {c12663};
    Full_Adder FA_13896(s13896, c13896, in13896_1, in13896_2, c12661);
    wire[0:0] s13897, in13897_1, in13897_2;
    wire c13897;
    assign in13897_1 = {s12665[0]};
    assign in13897_2 = {s12666[0]};
    Full_Adder FA_13897(s13897, c13897, in13897_1, in13897_2, s12664[0]);
    wire[0:0] s13898, in13898_1, in13898_2;
    wire c13898;
    assign in13898_1 = {s12668[0]};
    assign in13898_2 = {s12669[0]};
    Full_Adder FA_13898(s13898, c13898, in13898_1, in13898_2, s12667[0]);
    wire[0:0] s13899, in13899_1, in13899_2;
    wire c13899;
    assign in13899_1 = {c12665};
    assign in13899_2 = {c12666};
    Full_Adder FA_13899(s13899, c13899, in13899_1, in13899_2, c12664);
    wire[0:0] s13900, in13900_1, in13900_2;
    wire c13900;
    assign in13900_1 = {c12668};
    assign in13900_2 = {c12669};
    Full_Adder FA_13900(s13900, c13900, in13900_1, in13900_2, c12667);
    wire[0:0] s13901, in13901_1, in13901_2;
    wire c13901;
    assign in13901_1 = {s12671[0]};
    assign in13901_2 = {s12672[0]};
    Full_Adder FA_13901(s13901, c13901, in13901_1, in13901_2, s12670[0]);
    wire[0:0] s13902, in13902_1, in13902_2;
    wire c13902;
    assign in13902_1 = {s12674[0]};
    assign in13902_2 = {s12675[0]};
    Full_Adder FA_13902(s13902, c13902, in13902_1, in13902_2, s12673[0]);
    wire[0:0] s13903, in13903_1, in13903_2;
    wire c13903;
    assign in13903_1 = {c12671};
    assign in13903_2 = {c12672};
    Full_Adder FA_13903(s13903, c13903, in13903_1, in13903_2, c12670);
    wire[0:0] s13904, in13904_1, in13904_2;
    wire c13904;
    assign in13904_1 = {c12674};
    assign in13904_2 = {c12675};
    Full_Adder FA_13904(s13904, c13904, in13904_1, in13904_2, c12673);
    wire[0:0] s13905, in13905_1, in13905_2;
    wire c13905;
    assign in13905_1 = {s12677[0]};
    assign in13905_2 = {s12678[0]};
    Full_Adder FA_13905(s13905, c13905, in13905_1, in13905_2, s12676[0]);
    wire[0:0] s13906, in13906_1, in13906_2;
    wire c13906;
    assign in13906_1 = {s12680[0]};
    assign in13906_2 = {s12681[0]};
    Full_Adder FA_13906(s13906, c13906, in13906_1, in13906_2, s12679[0]);
    wire[0:0] s13907, in13907_1, in13907_2;
    wire c13907;
    assign in13907_1 = {c12677};
    assign in13907_2 = {c12678};
    Full_Adder FA_13907(s13907, c13907, in13907_1, in13907_2, c12676);
    wire[0:0] s13908, in13908_1, in13908_2;
    wire c13908;
    assign in13908_1 = {c12680};
    assign in13908_2 = {c12681};
    Full_Adder FA_13908(s13908, c13908, in13908_1, in13908_2, c12679);
    wire[0:0] s13909, in13909_1, in13909_2;
    wire c13909;
    assign in13909_1 = {s12683[0]};
    assign in13909_2 = {s12684[0]};
    Full_Adder FA_13909(s13909, c13909, in13909_1, in13909_2, s12682[0]);
    wire[0:0] s13910, in13910_1, in13910_2;
    wire c13910;
    assign in13910_1 = {s12686[0]};
    assign in13910_2 = {s12687[0]};
    Full_Adder FA_13910(s13910, c13910, in13910_1, in13910_2, s12685[0]);
    wire[0:0] s13911, in13911_1, in13911_2;
    wire c13911;
    assign in13911_1 = {c12683};
    assign in13911_2 = {c12684};
    Full_Adder FA_13911(s13911, c13911, in13911_1, in13911_2, c12682);
    wire[0:0] s13912, in13912_1, in13912_2;
    wire c13912;
    assign in13912_1 = {c12686};
    assign in13912_2 = {c12687};
    Full_Adder FA_13912(s13912, c13912, in13912_1, in13912_2, c12685);
    wire[0:0] s13913, in13913_1, in13913_2;
    wire c13913;
    assign in13913_1 = {s12689[0]};
    assign in13913_2 = {s12690[0]};
    Full_Adder FA_13913(s13913, c13913, in13913_1, in13913_2, s12688[0]);
    wire[0:0] s13914, in13914_1, in13914_2;
    wire c13914;
    assign in13914_1 = {s12692[0]};
    assign in13914_2 = {s12693[0]};
    Full_Adder FA_13914(s13914, c13914, in13914_1, in13914_2, s12691[0]);
    wire[0:0] s13915, in13915_1, in13915_2;
    wire c13915;
    assign in13915_1 = {c12689};
    assign in13915_2 = {c12690};
    Full_Adder FA_13915(s13915, c13915, in13915_1, in13915_2, c12688);
    wire[0:0] s13916, in13916_1, in13916_2;
    wire c13916;
    assign in13916_1 = {c12692};
    assign in13916_2 = {c12693};
    Full_Adder FA_13916(s13916, c13916, in13916_1, in13916_2, c12691);
    wire[0:0] s13917, in13917_1, in13917_2;
    wire c13917;
    assign in13917_1 = {s12695[0]};
    assign in13917_2 = {s12696[0]};
    Full_Adder FA_13917(s13917, c13917, in13917_1, in13917_2, s12694[0]);
    wire[0:0] s13918, in13918_1, in13918_2;
    wire c13918;
    assign in13918_1 = {s12698[0]};
    assign in13918_2 = {s12699[0]};
    Full_Adder FA_13918(s13918, c13918, in13918_1, in13918_2, s12697[0]);
    wire[0:0] s13919, in13919_1, in13919_2;
    wire c13919;
    assign in13919_1 = {c12695};
    assign in13919_2 = {c12696};
    Full_Adder FA_13919(s13919, c13919, in13919_1, in13919_2, c12694);
    wire[0:0] s13920, in13920_1, in13920_2;
    wire c13920;
    assign in13920_1 = {c12698};
    assign in13920_2 = {c12699};
    Full_Adder FA_13920(s13920, c13920, in13920_1, in13920_2, c12697);
    wire[0:0] s13921, in13921_1, in13921_2;
    wire c13921;
    assign in13921_1 = {s12701[0]};
    assign in13921_2 = {s12702[0]};
    Full_Adder FA_13921(s13921, c13921, in13921_1, in13921_2, s12700[0]);
    wire[0:0] s13922, in13922_1, in13922_2;
    wire c13922;
    assign in13922_1 = {s12704[0]};
    assign in13922_2 = {s12705[0]};
    Full_Adder FA_13922(s13922, c13922, in13922_1, in13922_2, s12703[0]);
    wire[0:0] s13923, in13923_1, in13923_2;
    wire c13923;
    assign in13923_1 = {c12701};
    assign in13923_2 = {c12702};
    Full_Adder FA_13923(s13923, c13923, in13923_1, in13923_2, c12700);
    wire[0:0] s13924, in13924_1, in13924_2;
    wire c13924;
    assign in13924_1 = {c12704};
    assign in13924_2 = {c12705};
    Full_Adder FA_13924(s13924, c13924, in13924_1, in13924_2, c12703);
    wire[0:0] s13925, in13925_1, in13925_2;
    wire c13925;
    assign in13925_1 = {s12707[0]};
    assign in13925_2 = {s12708[0]};
    Full_Adder FA_13925(s13925, c13925, in13925_1, in13925_2, s12706[0]);
    wire[0:0] s13926, in13926_1, in13926_2;
    wire c13926;
    assign in13926_1 = {s12710[0]};
    assign in13926_2 = {s12711[0]};
    Full_Adder FA_13926(s13926, c13926, in13926_1, in13926_2, s12709[0]);
    wire[0:0] s13927, in13927_1, in13927_2;
    wire c13927;
    assign in13927_1 = {c12707};
    assign in13927_2 = {c12708};
    Full_Adder FA_13927(s13927, c13927, in13927_1, in13927_2, c12706);
    wire[0:0] s13928, in13928_1, in13928_2;
    wire c13928;
    assign in13928_1 = {c12710};
    assign in13928_2 = {c12711};
    Full_Adder FA_13928(s13928, c13928, in13928_1, in13928_2, c12709);
    wire[0:0] s13929, in13929_1, in13929_2;
    wire c13929;
    assign in13929_1 = {s12713[0]};
    assign in13929_2 = {s12714[0]};
    Full_Adder FA_13929(s13929, c13929, in13929_1, in13929_2, s12712[0]);
    wire[0:0] s13930, in13930_1, in13930_2;
    wire c13930;
    assign in13930_1 = {s12716[0]};
    assign in13930_2 = {s12717[0]};
    Full_Adder FA_13930(s13930, c13930, in13930_1, in13930_2, s12715[0]);
    wire[0:0] s13931, in13931_1, in13931_2;
    wire c13931;
    assign in13931_1 = {c12713};
    assign in13931_2 = {c12714};
    Full_Adder FA_13931(s13931, c13931, in13931_1, in13931_2, c12712);
    wire[0:0] s13932, in13932_1, in13932_2;
    wire c13932;
    assign in13932_1 = {c12716};
    assign in13932_2 = {c12717};
    Full_Adder FA_13932(s13932, c13932, in13932_1, in13932_2, c12715);
    wire[0:0] s13933, in13933_1, in13933_2;
    wire c13933;
    assign in13933_1 = {s12719[0]};
    assign in13933_2 = {s12720[0]};
    Full_Adder FA_13933(s13933, c13933, in13933_1, in13933_2, s12718[0]);
    wire[0:0] s13934, in13934_1, in13934_2;
    wire c13934;
    assign in13934_1 = {s12722[0]};
    assign in13934_2 = {s12723[0]};
    Full_Adder FA_13934(s13934, c13934, in13934_1, in13934_2, s12721[0]);
    wire[0:0] s13935, in13935_1, in13935_2;
    wire c13935;
    assign in13935_1 = {c12719};
    assign in13935_2 = {c12720};
    Full_Adder FA_13935(s13935, c13935, in13935_1, in13935_2, c12718);
    wire[0:0] s13936, in13936_1, in13936_2;
    wire c13936;
    assign in13936_1 = {c12722};
    assign in13936_2 = {c12723};
    Full_Adder FA_13936(s13936, c13936, in13936_1, in13936_2, c12721);
    wire[0:0] s13937, in13937_1, in13937_2;
    wire c13937;
    assign in13937_1 = {s12725[0]};
    assign in13937_2 = {s12726[0]};
    Full_Adder FA_13937(s13937, c13937, in13937_1, in13937_2, s12724[0]);
    wire[0:0] s13938, in13938_1, in13938_2;
    wire c13938;
    assign in13938_1 = {s12728[0]};
    assign in13938_2 = {s12729[0]};
    Full_Adder FA_13938(s13938, c13938, in13938_1, in13938_2, s12727[0]);
    wire[0:0] s13939, in13939_1, in13939_2;
    wire c13939;
    assign in13939_1 = {c12725};
    assign in13939_2 = {c12726};
    Full_Adder FA_13939(s13939, c13939, in13939_1, in13939_2, c12724);
    wire[0:0] s13940, in13940_1, in13940_2;
    wire c13940;
    assign in13940_1 = {c12728};
    assign in13940_2 = {c12729};
    Full_Adder FA_13940(s13940, c13940, in13940_1, in13940_2, c12727);
    wire[0:0] s13941, in13941_1, in13941_2;
    wire c13941;
    assign in13941_1 = {s12731[0]};
    assign in13941_2 = {s12732[0]};
    Full_Adder FA_13941(s13941, c13941, in13941_1, in13941_2, s12730[0]);
    wire[0:0] s13942, in13942_1, in13942_2;
    wire c13942;
    assign in13942_1 = {s12734[0]};
    assign in13942_2 = {s12735[0]};
    Full_Adder FA_13942(s13942, c13942, in13942_1, in13942_2, s12733[0]);
    wire[0:0] s13943, in13943_1, in13943_2;
    wire c13943;
    assign in13943_1 = {c12731};
    assign in13943_2 = {c12732};
    Full_Adder FA_13943(s13943, c13943, in13943_1, in13943_2, c12730);
    wire[0:0] s13944, in13944_1, in13944_2;
    wire c13944;
    assign in13944_1 = {c12734};
    assign in13944_2 = {c12735};
    Full_Adder FA_13944(s13944, c13944, in13944_1, in13944_2, c12733);
    wire[0:0] s13945, in13945_1, in13945_2;
    wire c13945;
    assign in13945_1 = {s12737[0]};
    assign in13945_2 = {s12738[0]};
    Full_Adder FA_13945(s13945, c13945, in13945_1, in13945_2, s12736[0]);
    wire[0:0] s13946, in13946_1, in13946_2;
    wire c13946;
    assign in13946_1 = {s12740[0]};
    assign in13946_2 = {s12741[0]};
    Full_Adder FA_13946(s13946, c13946, in13946_1, in13946_2, s12739[0]);
    wire[0:0] s13947, in13947_1, in13947_2;
    wire c13947;
    assign in13947_1 = {c12737};
    assign in13947_2 = {c12738};
    Full_Adder FA_13947(s13947, c13947, in13947_1, in13947_2, c12736);
    wire[0:0] s13948, in13948_1, in13948_2;
    wire c13948;
    assign in13948_1 = {c12740};
    assign in13948_2 = {c12741};
    Full_Adder FA_13948(s13948, c13948, in13948_1, in13948_2, c12739);
    wire[0:0] s13949, in13949_1, in13949_2;
    wire c13949;
    assign in13949_1 = {s12743[0]};
    assign in13949_2 = {s12744[0]};
    Full_Adder FA_13949(s13949, c13949, in13949_1, in13949_2, s12742[0]);
    wire[0:0] s13950, in13950_1, in13950_2;
    wire c13950;
    assign in13950_1 = {s12746[0]};
    assign in13950_2 = {s12747[0]};
    Full_Adder FA_13950(s13950, c13950, in13950_1, in13950_2, s12745[0]);
    wire[0:0] s13951, in13951_1, in13951_2;
    wire c13951;
    assign in13951_1 = {c12743};
    assign in13951_2 = {c12744};
    Full_Adder FA_13951(s13951, c13951, in13951_1, in13951_2, c12742);
    wire[0:0] s13952, in13952_1, in13952_2;
    wire c13952;
    assign in13952_1 = {c12746};
    assign in13952_2 = {c12747};
    Full_Adder FA_13952(s13952, c13952, in13952_1, in13952_2, c12745);
    wire[0:0] s13953, in13953_1, in13953_2;
    wire c13953;
    assign in13953_1 = {s12749[0]};
    assign in13953_2 = {s12750[0]};
    Full_Adder FA_13953(s13953, c13953, in13953_1, in13953_2, s12748[0]);
    wire[0:0] s13954, in13954_1, in13954_2;
    wire c13954;
    assign in13954_1 = {s12752[0]};
    assign in13954_2 = {s12753[0]};
    Full_Adder FA_13954(s13954, c13954, in13954_1, in13954_2, s12751[0]);
    wire[0:0] s13955, in13955_1, in13955_2;
    wire c13955;
    assign in13955_1 = {c12749};
    assign in13955_2 = {c12750};
    Full_Adder FA_13955(s13955, c13955, in13955_1, in13955_2, c12748);
    wire[0:0] s13956, in13956_1, in13956_2;
    wire c13956;
    assign in13956_1 = {c12752};
    assign in13956_2 = {c12753};
    Full_Adder FA_13956(s13956, c13956, in13956_1, in13956_2, c12751);
    wire[0:0] s13957, in13957_1, in13957_2;
    wire c13957;
    assign in13957_1 = {s12755[0]};
    assign in13957_2 = {s12756[0]};
    Full_Adder FA_13957(s13957, c13957, in13957_1, in13957_2, s12754[0]);
    wire[0:0] s13958, in13958_1, in13958_2;
    wire c13958;
    assign in13958_1 = {s12758[0]};
    assign in13958_2 = {s12759[0]};
    Full_Adder FA_13958(s13958, c13958, in13958_1, in13958_2, s12757[0]);
    wire[0:0] s13959, in13959_1, in13959_2;
    wire c13959;
    assign in13959_1 = {c12755};
    assign in13959_2 = {c12756};
    Full_Adder FA_13959(s13959, c13959, in13959_1, in13959_2, c12754);
    wire[0:0] s13960, in13960_1, in13960_2;
    wire c13960;
    assign in13960_1 = {c12758};
    assign in13960_2 = {c12759};
    Full_Adder FA_13960(s13960, c13960, in13960_1, in13960_2, c12757);
    wire[0:0] s13961, in13961_1, in13961_2;
    wire c13961;
    assign in13961_1 = {s12761[0]};
    assign in13961_2 = {s12762[0]};
    Full_Adder FA_13961(s13961, c13961, in13961_1, in13961_2, s12760[0]);
    wire[0:0] s13962, in13962_1, in13962_2;
    wire c13962;
    assign in13962_1 = {s12764[0]};
    assign in13962_2 = {s12765[0]};
    Full_Adder FA_13962(s13962, c13962, in13962_1, in13962_2, s12763[0]);
    wire[0:0] s13963, in13963_1, in13963_2;
    wire c13963;
    assign in13963_1 = {c12761};
    assign in13963_2 = {c12762};
    Full_Adder FA_13963(s13963, c13963, in13963_1, in13963_2, c12760);
    wire[0:0] s13964, in13964_1, in13964_2;
    wire c13964;
    assign in13964_1 = {c12764};
    assign in13964_2 = {c12765};
    Full_Adder FA_13964(s13964, c13964, in13964_1, in13964_2, c12763);
    wire[0:0] s13965, in13965_1, in13965_2;
    wire c13965;
    assign in13965_1 = {s12767[0]};
    assign in13965_2 = {s12768[0]};
    Full_Adder FA_13965(s13965, c13965, in13965_1, in13965_2, s12766[0]);
    wire[0:0] s13966, in13966_1, in13966_2;
    wire c13966;
    assign in13966_1 = {s12770[0]};
    assign in13966_2 = {s12771[0]};
    Full_Adder FA_13966(s13966, c13966, in13966_1, in13966_2, s12769[0]);
    wire[0:0] s13967, in13967_1, in13967_2;
    wire c13967;
    assign in13967_1 = {c12767};
    assign in13967_2 = {c12768};
    Full_Adder FA_13967(s13967, c13967, in13967_1, in13967_2, c12766);
    wire[0:0] s13968, in13968_1, in13968_2;
    wire c13968;
    assign in13968_1 = {c12770};
    assign in13968_2 = {c12771};
    Full_Adder FA_13968(s13968, c13968, in13968_1, in13968_2, c12769);
    wire[0:0] s13969, in13969_1, in13969_2;
    wire c13969;
    assign in13969_1 = {s12773[0]};
    assign in13969_2 = {s12774[0]};
    Full_Adder FA_13969(s13969, c13969, in13969_1, in13969_2, s12772[0]);
    wire[0:0] s13970, in13970_1, in13970_2;
    wire c13970;
    assign in13970_1 = {s12776[0]};
    assign in13970_2 = {s12777[0]};
    Full_Adder FA_13970(s13970, c13970, in13970_1, in13970_2, s12775[0]);
    wire[0:0] s13971, in13971_1, in13971_2;
    wire c13971;
    assign in13971_1 = {c12773};
    assign in13971_2 = {c12774};
    Full_Adder FA_13971(s13971, c13971, in13971_1, in13971_2, c12772);
    wire[0:0] s13972, in13972_1, in13972_2;
    wire c13972;
    assign in13972_1 = {c12776};
    assign in13972_2 = {c12777};
    Full_Adder FA_13972(s13972, c13972, in13972_1, in13972_2, c12775);
    wire[0:0] s13973, in13973_1, in13973_2;
    wire c13973;
    assign in13973_1 = {s12779[0]};
    assign in13973_2 = {s12780[0]};
    Full_Adder FA_13973(s13973, c13973, in13973_1, in13973_2, s12778[0]);
    wire[0:0] s13974, in13974_1, in13974_2;
    wire c13974;
    assign in13974_1 = {s12782[0]};
    assign in13974_2 = {s12783[0]};
    Full_Adder FA_13974(s13974, c13974, in13974_1, in13974_2, s12781[0]);
    wire[0:0] s13975, in13975_1, in13975_2;
    wire c13975;
    assign in13975_1 = {c12779};
    assign in13975_2 = {c12780};
    Full_Adder FA_13975(s13975, c13975, in13975_1, in13975_2, c12778);
    wire[0:0] s13976, in13976_1, in13976_2;
    wire c13976;
    assign in13976_1 = {c12782};
    assign in13976_2 = {c12783};
    Full_Adder FA_13976(s13976, c13976, in13976_1, in13976_2, c12781);
    wire[0:0] s13977, in13977_1, in13977_2;
    wire c13977;
    assign in13977_1 = {s12785[0]};
    assign in13977_2 = {s12786[0]};
    Full_Adder FA_13977(s13977, c13977, in13977_1, in13977_2, s12784[0]);
    wire[0:0] s13978, in13978_1, in13978_2;
    wire c13978;
    assign in13978_1 = {s12788[0]};
    assign in13978_2 = {s12789[0]};
    Full_Adder FA_13978(s13978, c13978, in13978_1, in13978_2, s12787[0]);
    wire[0:0] s13979, in13979_1, in13979_2;
    wire c13979;
    assign in13979_1 = {c12785};
    assign in13979_2 = {c12786};
    Full_Adder FA_13979(s13979, c13979, in13979_1, in13979_2, c12784);
    wire[0:0] s13980, in13980_1, in13980_2;
    wire c13980;
    assign in13980_1 = {c12788};
    assign in13980_2 = {c12789};
    Full_Adder FA_13980(s13980, c13980, in13980_1, in13980_2, c12787);
    wire[0:0] s13981, in13981_1, in13981_2;
    wire c13981;
    assign in13981_1 = {s12791[0]};
    assign in13981_2 = {s12792[0]};
    Full_Adder FA_13981(s13981, c13981, in13981_1, in13981_2, s12790[0]);
    wire[0:0] s13982, in13982_1, in13982_2;
    wire c13982;
    assign in13982_1 = {s12794[0]};
    assign in13982_2 = {s12795[0]};
    Full_Adder FA_13982(s13982, c13982, in13982_1, in13982_2, s12793[0]);
    wire[0:0] s13983, in13983_1, in13983_2;
    wire c13983;
    assign in13983_1 = {c12791};
    assign in13983_2 = {c12792};
    Full_Adder FA_13983(s13983, c13983, in13983_1, in13983_2, c12790);
    wire[0:0] s13984, in13984_1, in13984_2;
    wire c13984;
    assign in13984_1 = {c12794};
    assign in13984_2 = {c12795};
    Full_Adder FA_13984(s13984, c13984, in13984_1, in13984_2, c12793);
    wire[0:0] s13985, in13985_1, in13985_2;
    wire c13985;
    assign in13985_1 = {s12797[0]};
    assign in13985_2 = {s12798[0]};
    Full_Adder FA_13985(s13985, c13985, in13985_1, in13985_2, s12796[0]);
    wire[0:0] s13986, in13986_1, in13986_2;
    wire c13986;
    assign in13986_1 = {s12800[0]};
    assign in13986_2 = {s12801[0]};
    Full_Adder FA_13986(s13986, c13986, in13986_1, in13986_2, s12799[0]);
    wire[0:0] s13987, in13987_1, in13987_2;
    wire c13987;
    assign in13987_1 = {c12797};
    assign in13987_2 = {c12798};
    Full_Adder FA_13987(s13987, c13987, in13987_1, in13987_2, c12796);
    wire[0:0] s13988, in13988_1, in13988_2;
    wire c13988;
    assign in13988_1 = {c12800};
    assign in13988_2 = {c12801};
    Full_Adder FA_13988(s13988, c13988, in13988_1, in13988_2, c12799);
    wire[0:0] s13989, in13989_1, in13989_2;
    wire c13989;
    assign in13989_1 = {s12803[0]};
    assign in13989_2 = {s12804[0]};
    Full_Adder FA_13989(s13989, c13989, in13989_1, in13989_2, s12802[0]);
    wire[0:0] s13990, in13990_1, in13990_2;
    wire c13990;
    assign in13990_1 = {s12806[0]};
    assign in13990_2 = {s12807[0]};
    Full_Adder FA_13990(s13990, c13990, in13990_1, in13990_2, s12805[0]);
    wire[0:0] s13991, in13991_1, in13991_2;
    wire c13991;
    assign in13991_1 = {c12803};
    assign in13991_2 = {c12804};
    Full_Adder FA_13991(s13991, c13991, in13991_1, in13991_2, c12802);
    wire[0:0] s13992, in13992_1, in13992_2;
    wire c13992;
    assign in13992_1 = {c12806};
    assign in13992_2 = {c12807};
    Full_Adder FA_13992(s13992, c13992, in13992_1, in13992_2, c12805);
    wire[0:0] s13993, in13993_1, in13993_2;
    wire c13993;
    assign in13993_1 = {s12809[0]};
    assign in13993_2 = {s12810[0]};
    Full_Adder FA_13993(s13993, c13993, in13993_1, in13993_2, s12808[0]);
    wire[0:0] s13994, in13994_1, in13994_2;
    wire c13994;
    assign in13994_1 = {s12812[0]};
    assign in13994_2 = {s12813[0]};
    Full_Adder FA_13994(s13994, c13994, in13994_1, in13994_2, s12811[0]);
    wire[0:0] s13995, in13995_1, in13995_2;
    wire c13995;
    assign in13995_1 = {c12809};
    assign in13995_2 = {c12810};
    Full_Adder FA_13995(s13995, c13995, in13995_1, in13995_2, c12808);
    wire[0:0] s13996, in13996_1, in13996_2;
    wire c13996;
    assign in13996_1 = {c12812};
    assign in13996_2 = {c12813};
    Full_Adder FA_13996(s13996, c13996, in13996_1, in13996_2, c12811);
    wire[0:0] s13997, in13997_1, in13997_2;
    wire c13997;
    assign in13997_1 = {s12815[0]};
    assign in13997_2 = {s12816[0]};
    Full_Adder FA_13997(s13997, c13997, in13997_1, in13997_2, s12814[0]);
    wire[0:0] s13998, in13998_1, in13998_2;
    wire c13998;
    assign in13998_1 = {s12818[0]};
    assign in13998_2 = {s12819[0]};
    Full_Adder FA_13998(s13998, c13998, in13998_1, in13998_2, s12817[0]);
    wire[0:0] s13999, in13999_1, in13999_2;
    wire c13999;
    assign in13999_1 = {c12815};
    assign in13999_2 = {c12816};
    Full_Adder FA_13999(s13999, c13999, in13999_1, in13999_2, c12814);
    wire[0:0] s14000, in14000_1, in14000_2;
    wire c14000;
    assign in14000_1 = {c12818};
    assign in14000_2 = {c12819};
    Full_Adder FA_14000(s14000, c14000, in14000_1, in14000_2, c12817);
    wire[0:0] s14001, in14001_1, in14001_2;
    wire c14001;
    assign in14001_1 = {s12821[0]};
    assign in14001_2 = {s12822[0]};
    Full_Adder FA_14001(s14001, c14001, in14001_1, in14001_2, s12820[0]);
    wire[0:0] s14002, in14002_1, in14002_2;
    wire c14002;
    assign in14002_1 = {s12824[0]};
    assign in14002_2 = {s12825[0]};
    Full_Adder FA_14002(s14002, c14002, in14002_1, in14002_2, s12823[0]);
    wire[0:0] s14003, in14003_1, in14003_2;
    wire c14003;
    assign in14003_1 = {c12821};
    assign in14003_2 = {c12822};
    Full_Adder FA_14003(s14003, c14003, in14003_1, in14003_2, c12820);
    wire[0:0] s14004, in14004_1, in14004_2;
    wire c14004;
    assign in14004_1 = {c12824};
    assign in14004_2 = {c12825};
    Full_Adder FA_14004(s14004, c14004, in14004_1, in14004_2, c12823);
    wire[0:0] s14005, in14005_1, in14005_2;
    wire c14005;
    assign in14005_1 = {s12827[0]};
    assign in14005_2 = {s12828[0]};
    Full_Adder FA_14005(s14005, c14005, in14005_1, in14005_2, s12826[0]);
    wire[0:0] s14006, in14006_1, in14006_2;
    wire c14006;
    assign in14006_1 = {s12830[0]};
    assign in14006_2 = {s12831[0]};
    Full_Adder FA_14006(s14006, c14006, in14006_1, in14006_2, s12829[0]);
    wire[0:0] s14007, in14007_1, in14007_2;
    wire c14007;
    assign in14007_1 = {c12827};
    assign in14007_2 = {c12828};
    Full_Adder FA_14007(s14007, c14007, in14007_1, in14007_2, c12826);
    wire[0:0] s14008, in14008_1, in14008_2;
    wire c14008;
    assign in14008_1 = {c12830};
    assign in14008_2 = {c12831};
    Full_Adder FA_14008(s14008, c14008, in14008_1, in14008_2, c12829);
    wire[0:0] s14009, in14009_1, in14009_2;
    wire c14009;
    assign in14009_1 = {s12833[0]};
    assign in14009_2 = {s12834[0]};
    Full_Adder FA_14009(s14009, c14009, in14009_1, in14009_2, s12832[0]);
    wire[0:0] s14010, in14010_1, in14010_2;
    wire c14010;
    assign in14010_1 = {s12836[0]};
    assign in14010_2 = {s12837[0]};
    Full_Adder FA_14010(s14010, c14010, in14010_1, in14010_2, s12835[0]);
    wire[0:0] s14011, in14011_1, in14011_2;
    wire c14011;
    assign in14011_1 = {c12833};
    assign in14011_2 = {c12834};
    Full_Adder FA_14011(s14011, c14011, in14011_1, in14011_2, c12832);
    wire[0:0] s14012, in14012_1, in14012_2;
    wire c14012;
    assign in14012_1 = {c12836};
    assign in14012_2 = {c12837};
    Full_Adder FA_14012(s14012, c14012, in14012_1, in14012_2, c12835);
    wire[0:0] s14013, in14013_1, in14013_2;
    wire c14013;
    assign in14013_1 = {s12839[0]};
    assign in14013_2 = {s12840[0]};
    Full_Adder FA_14013(s14013, c14013, in14013_1, in14013_2, s12838[0]);
    wire[0:0] s14014, in14014_1, in14014_2;
    wire c14014;
    assign in14014_1 = {s12842[0]};
    assign in14014_2 = {s12843[0]};
    Full_Adder FA_14014(s14014, c14014, in14014_1, in14014_2, s12841[0]);
    wire[0:0] s14015, in14015_1, in14015_2;
    wire c14015;
    assign in14015_1 = {c12839};
    assign in14015_2 = {c12840};
    Full_Adder FA_14015(s14015, c14015, in14015_1, in14015_2, c12838);
    wire[0:0] s14016, in14016_1, in14016_2;
    wire c14016;
    assign in14016_1 = {c12842};
    assign in14016_2 = {c12843};
    Full_Adder FA_14016(s14016, c14016, in14016_1, in14016_2, c12841);
    wire[0:0] s14017, in14017_1, in14017_2;
    wire c14017;
    assign in14017_1 = {s12845[0]};
    assign in14017_2 = {s12846[0]};
    Full_Adder FA_14017(s14017, c14017, in14017_1, in14017_2, s12844[0]);
    wire[0:0] s14018, in14018_1, in14018_2;
    wire c14018;
    assign in14018_1 = {s12848[0]};
    assign in14018_2 = {s12849[0]};
    Full_Adder FA_14018(s14018, c14018, in14018_1, in14018_2, s12847[0]);
    wire[0:0] s14019, in14019_1, in14019_2;
    wire c14019;
    assign in14019_1 = {c12845};
    assign in14019_2 = {c12846};
    Full_Adder FA_14019(s14019, c14019, in14019_1, in14019_2, c12844);
    wire[0:0] s14020, in14020_1, in14020_2;
    wire c14020;
    assign in14020_1 = {c12848};
    assign in14020_2 = {c12849};
    Full_Adder FA_14020(s14020, c14020, in14020_1, in14020_2, c12847);
    wire[0:0] s14021, in14021_1, in14021_2;
    wire c14021;
    assign in14021_1 = {s12851[0]};
    assign in14021_2 = {s12852[0]};
    Full_Adder FA_14021(s14021, c14021, in14021_1, in14021_2, s12850[0]);
    wire[0:0] s14022, in14022_1, in14022_2;
    wire c14022;
    assign in14022_1 = {s12854[0]};
    assign in14022_2 = {s12855[0]};
    Full_Adder FA_14022(s14022, c14022, in14022_1, in14022_2, s12853[0]);
    wire[0:0] s14023, in14023_1, in14023_2;
    wire c14023;
    assign in14023_1 = {c12851};
    assign in14023_2 = {c12852};
    Full_Adder FA_14023(s14023, c14023, in14023_1, in14023_2, c12850);
    wire[0:0] s14024, in14024_1, in14024_2;
    wire c14024;
    assign in14024_1 = {c12854};
    assign in14024_2 = {c12855};
    Full_Adder FA_14024(s14024, c14024, in14024_1, in14024_2, c12853);
    wire[0:0] s14025, in14025_1, in14025_2;
    wire c14025;
    assign in14025_1 = {s12857[0]};
    assign in14025_2 = {s12858[0]};
    Full_Adder FA_14025(s14025, c14025, in14025_1, in14025_2, s12856[0]);
    wire[0:0] s14026, in14026_1, in14026_2;
    wire c14026;
    assign in14026_1 = {s12860[0]};
    assign in14026_2 = {s12861[0]};
    Full_Adder FA_14026(s14026, c14026, in14026_1, in14026_2, s12859[0]);
    wire[0:0] s14027, in14027_1, in14027_2;
    wire c14027;
    assign in14027_1 = {c12857};
    assign in14027_2 = {c12858};
    Full_Adder FA_14027(s14027, c14027, in14027_1, in14027_2, c12856);
    wire[0:0] s14028, in14028_1, in14028_2;
    wire c14028;
    assign in14028_1 = {c12860};
    assign in14028_2 = {c12861};
    Full_Adder FA_14028(s14028, c14028, in14028_1, in14028_2, c12859);
    wire[0:0] s14029, in14029_1, in14029_2;
    wire c14029;
    assign in14029_1 = {s12863[0]};
    assign in14029_2 = {s12864[0]};
    Full_Adder FA_14029(s14029, c14029, in14029_1, in14029_2, s12862[0]);
    wire[0:0] s14030, in14030_1, in14030_2;
    wire c14030;
    assign in14030_1 = {s12866[0]};
    assign in14030_2 = {s12867[0]};
    Full_Adder FA_14030(s14030, c14030, in14030_1, in14030_2, s12865[0]);
    wire[0:0] s14031, in14031_1, in14031_2;
    wire c14031;
    assign in14031_1 = {c12863};
    assign in14031_2 = {c12864};
    Full_Adder FA_14031(s14031, c14031, in14031_1, in14031_2, c12862);
    wire[0:0] s14032, in14032_1, in14032_2;
    wire c14032;
    assign in14032_1 = {c12866};
    assign in14032_2 = {c12867};
    Full_Adder FA_14032(s14032, c14032, in14032_1, in14032_2, c12865);
    wire[0:0] s14033, in14033_1, in14033_2;
    wire c14033;
    assign in14033_1 = {s12869[0]};
    assign in14033_2 = {s12870[0]};
    Full_Adder FA_14033(s14033, c14033, in14033_1, in14033_2, s12868[0]);
    wire[0:0] s14034, in14034_1, in14034_2;
    wire c14034;
    assign in14034_1 = {s12872[0]};
    assign in14034_2 = {s12873[0]};
    Full_Adder FA_14034(s14034, c14034, in14034_1, in14034_2, s12871[0]);
    wire[0:0] s14035, in14035_1, in14035_2;
    wire c14035;
    assign in14035_1 = {c12869};
    assign in14035_2 = {c12870};
    Full_Adder FA_14035(s14035, c14035, in14035_1, in14035_2, c12868);
    wire[0:0] s14036, in14036_1, in14036_2;
    wire c14036;
    assign in14036_1 = {c12872};
    assign in14036_2 = {c12873};
    Full_Adder FA_14036(s14036, c14036, in14036_1, in14036_2, c12871);
    wire[0:0] s14037, in14037_1, in14037_2;
    wire c14037;
    assign in14037_1 = {s12875[0]};
    assign in14037_2 = {s12876[0]};
    Full_Adder FA_14037(s14037, c14037, in14037_1, in14037_2, s12874[0]);
    wire[0:0] s14038, in14038_1, in14038_2;
    wire c14038;
    assign in14038_1 = {s12878[0]};
    assign in14038_2 = {s12879[0]};
    Full_Adder FA_14038(s14038, c14038, in14038_1, in14038_2, s12877[0]);
    wire[0:0] s14039, in14039_1, in14039_2;
    wire c14039;
    assign in14039_1 = {c12875};
    assign in14039_2 = {c12876};
    Full_Adder FA_14039(s14039, c14039, in14039_1, in14039_2, c12874);
    wire[0:0] s14040, in14040_1, in14040_2;
    wire c14040;
    assign in14040_1 = {c12878};
    assign in14040_2 = {c12879};
    Full_Adder FA_14040(s14040, c14040, in14040_1, in14040_2, c12877);
    wire[0:0] s14041, in14041_1, in14041_2;
    wire c14041;
    assign in14041_1 = {s12881[0]};
    assign in14041_2 = {s12882[0]};
    Full_Adder FA_14041(s14041, c14041, in14041_1, in14041_2, s12880[0]);
    wire[0:0] s14042, in14042_1, in14042_2;
    wire c14042;
    assign in14042_1 = {s12884[0]};
    assign in14042_2 = {s12885[0]};
    Full_Adder FA_14042(s14042, c14042, in14042_1, in14042_2, s12883[0]);
    wire[0:0] s14043, in14043_1, in14043_2;
    wire c14043;
    assign in14043_1 = {c12881};
    assign in14043_2 = {c12882};
    Full_Adder FA_14043(s14043, c14043, in14043_1, in14043_2, c12880);
    wire[0:0] s14044, in14044_1, in14044_2;
    wire c14044;
    assign in14044_1 = {c12884};
    assign in14044_2 = {c12885};
    Full_Adder FA_14044(s14044, c14044, in14044_1, in14044_2, c12883);
    wire[0:0] s14045, in14045_1, in14045_2;
    wire c14045;
    assign in14045_1 = {s12887[0]};
    assign in14045_2 = {s12888[0]};
    Full_Adder FA_14045(s14045, c14045, in14045_1, in14045_2, s12886[0]);
    wire[0:0] s14046, in14046_1, in14046_2;
    wire c14046;
    assign in14046_1 = {s12890[0]};
    assign in14046_2 = {s12891[0]};
    Full_Adder FA_14046(s14046, c14046, in14046_1, in14046_2, s12889[0]);
    wire[0:0] s14047, in14047_1, in14047_2;
    wire c14047;
    assign in14047_1 = {c12887};
    assign in14047_2 = {c12888};
    Full_Adder FA_14047(s14047, c14047, in14047_1, in14047_2, c12886);
    wire[0:0] s14048, in14048_1, in14048_2;
    wire c14048;
    assign in14048_1 = {c12890};
    assign in14048_2 = {c12891};
    Full_Adder FA_14048(s14048, c14048, in14048_1, in14048_2, c12889);
    wire[0:0] s14049, in14049_1, in14049_2;
    wire c14049;
    assign in14049_1 = {s12893[0]};
    assign in14049_2 = {s12894[0]};
    Full_Adder FA_14049(s14049, c14049, in14049_1, in14049_2, s12892[0]);
    wire[0:0] s14050, in14050_1, in14050_2;
    wire c14050;
    assign in14050_1 = {s12896[0]};
    assign in14050_2 = {s12897[0]};
    Full_Adder FA_14050(s14050, c14050, in14050_1, in14050_2, s12895[0]);
    wire[0:0] s14051, in14051_1, in14051_2;
    wire c14051;
    assign in14051_1 = {c12893};
    assign in14051_2 = {c12894};
    Full_Adder FA_14051(s14051, c14051, in14051_1, in14051_2, c12892);
    wire[0:0] s14052, in14052_1, in14052_2;
    wire c14052;
    assign in14052_1 = {c12896};
    assign in14052_2 = {c12897};
    Full_Adder FA_14052(s14052, c14052, in14052_1, in14052_2, c12895);
    wire[0:0] s14053, in14053_1, in14053_2;
    wire c14053;
    assign in14053_1 = {s12899[0]};
    assign in14053_2 = {s12900[0]};
    Full_Adder FA_14053(s14053, c14053, in14053_1, in14053_2, s12898[0]);
    wire[0:0] s14054, in14054_1, in14054_2;
    wire c14054;
    assign in14054_1 = {s12902[0]};
    assign in14054_2 = {s12903[0]};
    Full_Adder FA_14054(s14054, c14054, in14054_1, in14054_2, s12901[0]);
    wire[0:0] s14055, in14055_1, in14055_2;
    wire c14055;
    assign in14055_1 = {c12899};
    assign in14055_2 = {c12900};
    Full_Adder FA_14055(s14055, c14055, in14055_1, in14055_2, c12898);
    wire[0:0] s14056, in14056_1, in14056_2;
    wire c14056;
    assign in14056_1 = {c12902};
    assign in14056_2 = {c12903};
    Full_Adder FA_14056(s14056, c14056, in14056_1, in14056_2, c12901);
    wire[0:0] s14057, in14057_1, in14057_2;
    wire c14057;
    assign in14057_1 = {s12905[0]};
    assign in14057_2 = {s12906[0]};
    Full_Adder FA_14057(s14057, c14057, in14057_1, in14057_2, s12904[0]);
    wire[0:0] s14058, in14058_1, in14058_2;
    wire c14058;
    assign in14058_1 = {s12908[0]};
    assign in14058_2 = {s12909[0]};
    Full_Adder FA_14058(s14058, c14058, in14058_1, in14058_2, s12907[0]);
    wire[0:0] s14059, in14059_1, in14059_2;
    wire c14059;
    assign in14059_1 = {c12905};
    assign in14059_2 = {c12906};
    Full_Adder FA_14059(s14059, c14059, in14059_1, in14059_2, c12904);
    wire[0:0] s14060, in14060_1, in14060_2;
    wire c14060;
    assign in14060_1 = {c12908};
    assign in14060_2 = {c12909};
    Full_Adder FA_14060(s14060, c14060, in14060_1, in14060_2, c12907);
    wire[0:0] s14061, in14061_1, in14061_2;
    wire c14061;
    assign in14061_1 = {s12911[0]};
    assign in14061_2 = {s12912[0]};
    Full_Adder FA_14061(s14061, c14061, in14061_1, in14061_2, s12910[0]);
    wire[0:0] s14062, in14062_1, in14062_2;
    wire c14062;
    assign in14062_1 = {s12914[0]};
    assign in14062_2 = {s12915[0]};
    Full_Adder FA_14062(s14062, c14062, in14062_1, in14062_2, s12913[0]);
    wire[0:0] s14063, in14063_1, in14063_2;
    wire c14063;
    assign in14063_1 = {c12911};
    assign in14063_2 = {c12912};
    Full_Adder FA_14063(s14063, c14063, in14063_1, in14063_2, c12910);
    wire[0:0] s14064, in14064_1, in14064_2;
    wire c14064;
    assign in14064_1 = {c12914};
    assign in14064_2 = {c12915};
    Full_Adder FA_14064(s14064, c14064, in14064_1, in14064_2, c12913);
    wire[0:0] s14065, in14065_1, in14065_2;
    wire c14065;
    assign in14065_1 = {s12917[0]};
    assign in14065_2 = {s12918[0]};
    Full_Adder FA_14065(s14065, c14065, in14065_1, in14065_2, s12916[0]);
    wire[0:0] s14066, in14066_1, in14066_2;
    wire c14066;
    assign in14066_1 = {s12920[0]};
    assign in14066_2 = {s12921[0]};
    Full_Adder FA_14066(s14066, c14066, in14066_1, in14066_2, s12919[0]);
    wire[0:0] s14067, in14067_1, in14067_2;
    wire c14067;
    assign in14067_1 = {c12917};
    assign in14067_2 = {c12918};
    Full_Adder FA_14067(s14067, c14067, in14067_1, in14067_2, c12916);
    wire[0:0] s14068, in14068_1, in14068_2;
    wire c14068;
    assign in14068_1 = {c12920};
    assign in14068_2 = {c12921};
    Full_Adder FA_14068(s14068, c14068, in14068_1, in14068_2, c12919);
    wire[0:0] s14069, in14069_1, in14069_2;
    wire c14069;
    assign in14069_1 = {s12923[0]};
    assign in14069_2 = {s12924[0]};
    Full_Adder FA_14069(s14069, c14069, in14069_1, in14069_2, s12922[0]);
    wire[0:0] s14070, in14070_1, in14070_2;
    wire c14070;
    assign in14070_1 = {s12926[0]};
    assign in14070_2 = {s12927[0]};
    Full_Adder FA_14070(s14070, c14070, in14070_1, in14070_2, s12925[0]);
    wire[0:0] s14071, in14071_1, in14071_2;
    wire c14071;
    assign in14071_1 = {c12923};
    assign in14071_2 = {c12924};
    Full_Adder FA_14071(s14071, c14071, in14071_1, in14071_2, c12922);
    wire[0:0] s14072, in14072_1, in14072_2;
    wire c14072;
    assign in14072_1 = {c12926};
    assign in14072_2 = {c12927};
    Full_Adder FA_14072(s14072, c14072, in14072_1, in14072_2, c12925);
    wire[0:0] s14073, in14073_1, in14073_2;
    wire c14073;
    assign in14073_1 = {s12929[0]};
    assign in14073_2 = {s12930[0]};
    Full_Adder FA_14073(s14073, c14073, in14073_1, in14073_2, s12928[0]);
    wire[0:0] s14074, in14074_1, in14074_2;
    wire c14074;
    assign in14074_1 = {s12932[0]};
    assign in14074_2 = {s12933[0]};
    Full_Adder FA_14074(s14074, c14074, in14074_1, in14074_2, s12931[0]);
    wire[0:0] s14075, in14075_1, in14075_2;
    wire c14075;
    assign in14075_1 = {c12929};
    assign in14075_2 = {c12930};
    Full_Adder FA_14075(s14075, c14075, in14075_1, in14075_2, c12928);
    wire[0:0] s14076, in14076_1, in14076_2;
    wire c14076;
    assign in14076_1 = {c12932};
    assign in14076_2 = {c12933};
    Full_Adder FA_14076(s14076, c14076, in14076_1, in14076_2, c12931);
    wire[0:0] s14077, in14077_1, in14077_2;
    wire c14077;
    assign in14077_1 = {s12935[0]};
    assign in14077_2 = {s12936[0]};
    Full_Adder FA_14077(s14077, c14077, in14077_1, in14077_2, s12934[0]);
    wire[0:0] s14078, in14078_1, in14078_2;
    wire c14078;
    assign in14078_1 = {s12938[0]};
    assign in14078_2 = {s12939[0]};
    Full_Adder FA_14078(s14078, c14078, in14078_1, in14078_2, s12937[0]);
    wire[0:0] s14079, in14079_1, in14079_2;
    wire c14079;
    assign in14079_1 = {c12935};
    assign in14079_2 = {c12936};
    Full_Adder FA_14079(s14079, c14079, in14079_1, in14079_2, c12934);
    wire[0:0] s14080, in14080_1, in14080_2;
    wire c14080;
    assign in14080_1 = {c12938};
    assign in14080_2 = {c12939};
    Full_Adder FA_14080(s14080, c14080, in14080_1, in14080_2, c12937);
    wire[0:0] s14081, in14081_1, in14081_2;
    wire c14081;
    assign in14081_1 = {s12941[0]};
    assign in14081_2 = {s12942[0]};
    Full_Adder FA_14081(s14081, c14081, in14081_1, in14081_2, s12940[0]);
    wire[0:0] s14082, in14082_1, in14082_2;
    wire c14082;
    assign in14082_1 = {s12944[0]};
    assign in14082_2 = {s12945[0]};
    Full_Adder FA_14082(s14082, c14082, in14082_1, in14082_2, s12943[0]);
    wire[0:0] s14083, in14083_1, in14083_2;
    wire c14083;
    assign in14083_1 = {c12941};
    assign in14083_2 = {c12942};
    Full_Adder FA_14083(s14083, c14083, in14083_1, in14083_2, c12940);
    wire[0:0] s14084, in14084_1, in14084_2;
    wire c14084;
    assign in14084_1 = {c12944};
    assign in14084_2 = {c12945};
    Full_Adder FA_14084(s14084, c14084, in14084_1, in14084_2, c12943);
    wire[0:0] s14085, in14085_1, in14085_2;
    wire c14085;
    assign in14085_1 = {s12947[0]};
    assign in14085_2 = {s12948[0]};
    Full_Adder FA_14085(s14085, c14085, in14085_1, in14085_2, s12946[0]);
    wire[0:0] s14086, in14086_1, in14086_2;
    wire c14086;
    assign in14086_1 = {s12950[0]};
    assign in14086_2 = {s12951[0]};
    Full_Adder FA_14086(s14086, c14086, in14086_1, in14086_2, s12949[0]);
    wire[0:0] s14087, in14087_1, in14087_2;
    wire c14087;
    assign in14087_1 = {c12947};
    assign in14087_2 = {c12948};
    Full_Adder FA_14087(s14087, c14087, in14087_1, in14087_2, c12946);
    wire[0:0] s14088, in14088_1, in14088_2;
    wire c14088;
    assign in14088_1 = {c12950};
    assign in14088_2 = {c12951};
    Full_Adder FA_14088(s14088, c14088, in14088_1, in14088_2, c12949);
    wire[0:0] s14089, in14089_1, in14089_2;
    wire c14089;
    assign in14089_1 = {s12953[0]};
    assign in14089_2 = {s12954[0]};
    Full_Adder FA_14089(s14089, c14089, in14089_1, in14089_2, s12952[0]);
    wire[0:0] s14090, in14090_1, in14090_2;
    wire c14090;
    assign in14090_1 = {s12956[0]};
    assign in14090_2 = {s12957[0]};
    Full_Adder FA_14090(s14090, c14090, in14090_1, in14090_2, s12955[0]);
    wire[0:0] s14091, in14091_1, in14091_2;
    wire c14091;
    assign in14091_1 = {c12953};
    assign in14091_2 = {c12954};
    Full_Adder FA_14091(s14091, c14091, in14091_1, in14091_2, c12952);
    wire[0:0] s14092, in14092_1, in14092_2;
    wire c14092;
    assign in14092_1 = {c12956};
    assign in14092_2 = {c12957};
    Full_Adder FA_14092(s14092, c14092, in14092_1, in14092_2, c12955);
    wire[0:0] s14093, in14093_1, in14093_2;
    wire c14093;
    assign in14093_1 = {s12959[0]};
    assign in14093_2 = {s12960[0]};
    Full_Adder FA_14093(s14093, c14093, in14093_1, in14093_2, s12958[0]);
    wire[0:0] s14094, in14094_1, in14094_2;
    wire c14094;
    assign in14094_1 = {s12962[0]};
    assign in14094_2 = {s12963[0]};
    Full_Adder FA_14094(s14094, c14094, in14094_1, in14094_2, s12961[0]);
    wire[0:0] s14095, in14095_1, in14095_2;
    wire c14095;
    assign in14095_1 = {c12959};
    assign in14095_2 = {c12960};
    Full_Adder FA_14095(s14095, c14095, in14095_1, in14095_2, c12958);
    wire[0:0] s14096, in14096_1, in14096_2;
    wire c14096;
    assign in14096_1 = {c12962};
    assign in14096_2 = {c12963};
    Full_Adder FA_14096(s14096, c14096, in14096_1, in14096_2, c12961);
    wire[0:0] s14097, in14097_1, in14097_2;
    wire c14097;
    assign in14097_1 = {s12965[0]};
    assign in14097_2 = {s12966[0]};
    Full_Adder FA_14097(s14097, c14097, in14097_1, in14097_2, s12964[0]);
    wire[0:0] s14098, in14098_1, in14098_2;
    wire c14098;
    assign in14098_1 = {s12968[0]};
    assign in14098_2 = {s12969[0]};
    Full_Adder FA_14098(s14098, c14098, in14098_1, in14098_2, s12967[0]);
    wire[0:0] s14099, in14099_1, in14099_2;
    wire c14099;
    assign in14099_1 = {c12965};
    assign in14099_2 = {c12966};
    Full_Adder FA_14099(s14099, c14099, in14099_1, in14099_2, c12964);
    wire[0:0] s14100, in14100_1, in14100_2;
    wire c14100;
    assign in14100_1 = {c12968};
    assign in14100_2 = {c12969};
    Full_Adder FA_14100(s14100, c14100, in14100_1, in14100_2, c12967);
    wire[0:0] s14101, in14101_1, in14101_2;
    wire c14101;
    assign in14101_1 = {s12971[0]};
    assign in14101_2 = {s12972[0]};
    Full_Adder FA_14101(s14101, c14101, in14101_1, in14101_2, s12970[0]);
    wire[0:0] s14102, in14102_1, in14102_2;
    wire c14102;
    assign in14102_1 = {s12974[0]};
    assign in14102_2 = {s12975[0]};
    Full_Adder FA_14102(s14102, c14102, in14102_1, in14102_2, s12973[0]);
    wire[0:0] s14103, in14103_1, in14103_2;
    wire c14103;
    assign in14103_1 = {c12971};
    assign in14103_2 = {c12972};
    Full_Adder FA_14103(s14103, c14103, in14103_1, in14103_2, c12970);
    wire[0:0] s14104, in14104_1, in14104_2;
    wire c14104;
    assign in14104_1 = {c12974};
    assign in14104_2 = {c12975};
    Full_Adder FA_14104(s14104, c14104, in14104_1, in14104_2, c12973);
    wire[0:0] s14105, in14105_1, in14105_2;
    wire c14105;
    assign in14105_1 = {s12977[0]};
    assign in14105_2 = {s12978[0]};
    Full_Adder FA_14105(s14105, c14105, in14105_1, in14105_2, s12976[0]);
    wire[0:0] s14106, in14106_1, in14106_2;
    wire c14106;
    assign in14106_1 = {s12980[0]};
    assign in14106_2 = {s12981[0]};
    Full_Adder FA_14106(s14106, c14106, in14106_1, in14106_2, s12979[0]);
    wire[0:0] s14107, in14107_1, in14107_2;
    wire c14107;
    assign in14107_1 = {c12977};
    assign in14107_2 = {c12978};
    Full_Adder FA_14107(s14107, c14107, in14107_1, in14107_2, c12976);
    wire[0:0] s14108, in14108_1, in14108_2;
    wire c14108;
    assign in14108_1 = {c12980};
    assign in14108_2 = {c12981};
    Full_Adder FA_14108(s14108, c14108, in14108_1, in14108_2, c12979);
    wire[0:0] s14109, in14109_1, in14109_2;
    wire c14109;
    assign in14109_1 = {s12983[0]};
    assign in14109_2 = {s12984[0]};
    Full_Adder FA_14109(s14109, c14109, in14109_1, in14109_2, s12982[0]);
    wire[0:0] s14110, in14110_1, in14110_2;
    wire c14110;
    assign in14110_1 = {s12986[0]};
    assign in14110_2 = {s12987[0]};
    Full_Adder FA_14110(s14110, c14110, in14110_1, in14110_2, s12985[0]);
    wire[0:0] s14111, in14111_1, in14111_2;
    wire c14111;
    assign in14111_1 = {c12983};
    assign in14111_2 = {c12984};
    Full_Adder FA_14111(s14111, c14111, in14111_1, in14111_2, c12982);
    wire[0:0] s14112, in14112_1, in14112_2;
    wire c14112;
    assign in14112_1 = {c12986};
    assign in14112_2 = {c12987};
    Full_Adder FA_14112(s14112, c14112, in14112_1, in14112_2, c12985);
    wire[0:0] s14113, in14113_1, in14113_2;
    wire c14113;
    assign in14113_1 = {s12989[0]};
    assign in14113_2 = {s12990[0]};
    Full_Adder FA_14113(s14113, c14113, in14113_1, in14113_2, s12988[0]);
    wire[0:0] s14114, in14114_1, in14114_2;
    wire c14114;
    assign in14114_1 = {s12992[0]};
    assign in14114_2 = {s12993[0]};
    Full_Adder FA_14114(s14114, c14114, in14114_1, in14114_2, s12991[0]);
    wire[0:0] s14115, in14115_1, in14115_2;
    wire c14115;
    assign in14115_1 = {c12989};
    assign in14115_2 = {c12990};
    Full_Adder FA_14115(s14115, c14115, in14115_1, in14115_2, c12988);
    wire[0:0] s14116, in14116_1, in14116_2;
    wire c14116;
    assign in14116_1 = {c12992};
    assign in14116_2 = {c12993};
    Full_Adder FA_14116(s14116, c14116, in14116_1, in14116_2, c12991);
    wire[0:0] s14117, in14117_1, in14117_2;
    wire c14117;
    assign in14117_1 = {s12995[0]};
    assign in14117_2 = {s12996[0]};
    Full_Adder FA_14117(s14117, c14117, in14117_1, in14117_2, s12994[0]);
    wire[0:0] s14118, in14118_1, in14118_2;
    wire c14118;
    assign in14118_1 = {s12998[0]};
    assign in14118_2 = {s12999[0]};
    Full_Adder FA_14118(s14118, c14118, in14118_1, in14118_2, s12997[0]);
    wire[0:0] s14119, in14119_1, in14119_2;
    wire c14119;
    assign in14119_1 = {c12995};
    assign in14119_2 = {c12996};
    Full_Adder FA_14119(s14119, c14119, in14119_1, in14119_2, c12994);
    wire[0:0] s14120, in14120_1, in14120_2;
    wire c14120;
    assign in14120_1 = {c12998};
    assign in14120_2 = {c12999};
    Full_Adder FA_14120(s14120, c14120, in14120_1, in14120_2, c12997);
    wire[0:0] s14121, in14121_1, in14121_2;
    wire c14121;
    assign in14121_1 = {s13001[0]};
    assign in14121_2 = {s13002[0]};
    Full_Adder FA_14121(s14121, c14121, in14121_1, in14121_2, s13000[0]);
    wire[0:0] s14122, in14122_1, in14122_2;
    wire c14122;
    assign in14122_1 = {s13004[0]};
    assign in14122_2 = {s13005[0]};
    Full_Adder FA_14122(s14122, c14122, in14122_1, in14122_2, s13003[0]);
    wire[0:0] s14123, in14123_1, in14123_2;
    wire c14123;
    assign in14123_1 = {c13001};
    assign in14123_2 = {c13002};
    Full_Adder FA_14123(s14123, c14123, in14123_1, in14123_2, c13000);
    wire[0:0] s14124, in14124_1, in14124_2;
    wire c14124;
    assign in14124_1 = {c13004};
    assign in14124_2 = {c13005};
    Full_Adder FA_14124(s14124, c14124, in14124_1, in14124_2, c13003);
    wire[0:0] s14125, in14125_1, in14125_2;
    wire c14125;
    assign in14125_1 = {s13007[0]};
    assign in14125_2 = {s13008[0]};
    Full_Adder FA_14125(s14125, c14125, in14125_1, in14125_2, s13006[0]);
    wire[0:0] s14126, in14126_1, in14126_2;
    wire c14126;
    assign in14126_1 = {s13010[0]};
    assign in14126_2 = {s13011[0]};
    Full_Adder FA_14126(s14126, c14126, in14126_1, in14126_2, s13009[0]);
    wire[0:0] s14127, in14127_1, in14127_2;
    wire c14127;
    assign in14127_1 = {c13007};
    assign in14127_2 = {c13008};
    Full_Adder FA_14127(s14127, c14127, in14127_1, in14127_2, c13006);
    wire[0:0] s14128, in14128_1, in14128_2;
    wire c14128;
    assign in14128_1 = {c13010};
    assign in14128_2 = {c13011};
    Full_Adder FA_14128(s14128, c14128, in14128_1, in14128_2, c13009);
    wire[0:0] s14129, in14129_1, in14129_2;
    wire c14129;
    assign in14129_1 = {s13013[0]};
    assign in14129_2 = {s13014[0]};
    Full_Adder FA_14129(s14129, c14129, in14129_1, in14129_2, s13012[0]);
    wire[0:0] s14130, in14130_1, in14130_2;
    wire c14130;
    assign in14130_1 = {s13016[0]};
    assign in14130_2 = {s13017[0]};
    Full_Adder FA_14130(s14130, c14130, in14130_1, in14130_2, s13015[0]);
    wire[0:0] s14131, in14131_1, in14131_2;
    wire c14131;
    assign in14131_1 = {c13013};
    assign in14131_2 = {c13014};
    Full_Adder FA_14131(s14131, c14131, in14131_1, in14131_2, c13012);
    wire[0:0] s14132, in14132_1, in14132_2;
    wire c14132;
    assign in14132_1 = {c13016};
    assign in14132_2 = {c13017};
    Full_Adder FA_14132(s14132, c14132, in14132_1, in14132_2, c13015);
    wire[0:0] s14133, in14133_1, in14133_2;
    wire c14133;
    assign in14133_1 = {s13019[0]};
    assign in14133_2 = {s13020[0]};
    Full_Adder FA_14133(s14133, c14133, in14133_1, in14133_2, s13018[0]);
    wire[0:0] s14134, in14134_1, in14134_2;
    wire c14134;
    assign in14134_1 = {s13022[0]};
    assign in14134_2 = {s13023[0]};
    Full_Adder FA_14134(s14134, c14134, in14134_1, in14134_2, s13021[0]);
    wire[0:0] s14135, in14135_1, in14135_2;
    wire c14135;
    assign in14135_1 = {c13019};
    assign in14135_2 = {c13020};
    Full_Adder FA_14135(s14135, c14135, in14135_1, in14135_2, c13018);
    wire[0:0] s14136, in14136_1, in14136_2;
    wire c14136;
    assign in14136_1 = {c13022};
    assign in14136_2 = {c13023};
    Full_Adder FA_14136(s14136, c14136, in14136_1, in14136_2, c13021);
    wire[0:0] s14137, in14137_1, in14137_2;
    wire c14137;
    assign in14137_1 = {s13025[0]};
    assign in14137_2 = {s13026[0]};
    Full_Adder FA_14137(s14137, c14137, in14137_1, in14137_2, s13024[0]);
    wire[0:0] s14138, in14138_1, in14138_2;
    wire c14138;
    assign in14138_1 = {s13028[0]};
    assign in14138_2 = {s13029[0]};
    Full_Adder FA_14138(s14138, c14138, in14138_1, in14138_2, s13027[0]);
    wire[0:0] s14139, in14139_1, in14139_2;
    wire c14139;
    assign in14139_1 = {c13025};
    assign in14139_2 = {c13026};
    Full_Adder FA_14139(s14139, c14139, in14139_1, in14139_2, c13024);
    wire[0:0] s14140, in14140_1, in14140_2;
    wire c14140;
    assign in14140_1 = {c13028};
    assign in14140_2 = {c13029};
    Full_Adder FA_14140(s14140, c14140, in14140_1, in14140_2, c13027);
    wire[0:0] s14141, in14141_1, in14141_2;
    wire c14141;
    assign in14141_1 = {s13031[0]};
    assign in14141_2 = {s13032[0]};
    Full_Adder FA_14141(s14141, c14141, in14141_1, in14141_2, s13030[0]);
    wire[0:0] s14142, in14142_1, in14142_2;
    wire c14142;
    assign in14142_1 = {s13034[0]};
    assign in14142_2 = {s13035[0]};
    Full_Adder FA_14142(s14142, c14142, in14142_1, in14142_2, s13033[0]);
    wire[0:0] s14143, in14143_1, in14143_2;
    wire c14143;
    assign in14143_1 = {c13031};
    assign in14143_2 = {c13032};
    Full_Adder FA_14143(s14143, c14143, in14143_1, in14143_2, c13030);
    wire[0:0] s14144, in14144_1, in14144_2;
    wire c14144;
    assign in14144_1 = {c13034};
    assign in14144_2 = {c13035};
    Full_Adder FA_14144(s14144, c14144, in14144_1, in14144_2, c13033);
    wire[0:0] s14145, in14145_1, in14145_2;
    wire c14145;
    assign in14145_1 = {s13037[0]};
    assign in14145_2 = {s13038[0]};
    Full_Adder FA_14145(s14145, c14145, in14145_1, in14145_2, s13036[0]);
    wire[0:0] s14146, in14146_1, in14146_2;
    wire c14146;
    assign in14146_1 = {s13040[0]};
    assign in14146_2 = {s13041[0]};
    Full_Adder FA_14146(s14146, c14146, in14146_1, in14146_2, s13039[0]);
    wire[0:0] s14147, in14147_1, in14147_2;
    wire c14147;
    assign in14147_1 = {c13037};
    assign in14147_2 = {c13038};
    Full_Adder FA_14147(s14147, c14147, in14147_1, in14147_2, c13036);
    wire[0:0] s14148, in14148_1, in14148_2;
    wire c14148;
    assign in14148_1 = {c13040};
    assign in14148_2 = {c13041};
    Full_Adder FA_14148(s14148, c14148, in14148_1, in14148_2, c13039);
    wire[0:0] s14149, in14149_1, in14149_2;
    wire c14149;
    assign in14149_1 = {s13043[0]};
    assign in14149_2 = {s13044[0]};
    Full_Adder FA_14149(s14149, c14149, in14149_1, in14149_2, s13042[0]);
    wire[0:0] s14150, in14150_1, in14150_2;
    wire c14150;
    assign in14150_1 = {s13046[0]};
    assign in14150_2 = {s13047[0]};
    Full_Adder FA_14150(s14150, c14150, in14150_1, in14150_2, s13045[0]);
    wire[0:0] s14151, in14151_1, in14151_2;
    wire c14151;
    assign in14151_1 = {c13043};
    assign in14151_2 = {c13044};
    Full_Adder FA_14151(s14151, c14151, in14151_1, in14151_2, c13042);
    wire[0:0] s14152, in14152_1, in14152_2;
    wire c14152;
    assign in14152_1 = {c13046};
    assign in14152_2 = {c13047};
    Full_Adder FA_14152(s14152, c14152, in14152_1, in14152_2, c13045);
    wire[0:0] s14153, in14153_1, in14153_2;
    wire c14153;
    assign in14153_1 = {s13049[0]};
    assign in14153_2 = {s13050[0]};
    Full_Adder FA_14153(s14153, c14153, in14153_1, in14153_2, s13048[0]);
    wire[0:0] s14154, in14154_1, in14154_2;
    wire c14154;
    assign in14154_1 = {s13052[0]};
    assign in14154_2 = {s13053[0]};
    Full_Adder FA_14154(s14154, c14154, in14154_1, in14154_2, s13051[0]);
    wire[0:0] s14155, in14155_1, in14155_2;
    wire c14155;
    assign in14155_1 = {c13049};
    assign in14155_2 = {c13050};
    Full_Adder FA_14155(s14155, c14155, in14155_1, in14155_2, c13048);
    wire[0:0] s14156, in14156_1, in14156_2;
    wire c14156;
    assign in14156_1 = {c13052};
    assign in14156_2 = {c13053};
    Full_Adder FA_14156(s14156, c14156, in14156_1, in14156_2, c13051);
    wire[0:0] s14157, in14157_1, in14157_2;
    wire c14157;
    assign in14157_1 = {s13055[0]};
    assign in14157_2 = {s13056[0]};
    Full_Adder FA_14157(s14157, c14157, in14157_1, in14157_2, s13054[0]);
    wire[0:0] s14158, in14158_1, in14158_2;
    wire c14158;
    assign in14158_1 = {s13058[0]};
    assign in14158_2 = {s13059[0]};
    Full_Adder FA_14158(s14158, c14158, in14158_1, in14158_2, s13057[0]);
    wire[0:0] s14159, in14159_1, in14159_2;
    wire c14159;
    assign in14159_1 = {c13055};
    assign in14159_2 = {c13056};
    Full_Adder FA_14159(s14159, c14159, in14159_1, in14159_2, c13054);
    wire[0:0] s14160, in14160_1, in14160_2;
    wire c14160;
    assign in14160_1 = {c13058};
    assign in14160_2 = {c13059};
    Full_Adder FA_14160(s14160, c14160, in14160_1, in14160_2, c13057);
    wire[0:0] s14161, in14161_1, in14161_2;
    wire c14161;
    assign in14161_1 = {s13061[0]};
    assign in14161_2 = {s13062[0]};
    Full_Adder FA_14161(s14161, c14161, in14161_1, in14161_2, s13060[0]);
    wire[0:0] s14162, in14162_1, in14162_2;
    wire c14162;
    assign in14162_1 = {s13064[0]};
    assign in14162_2 = {s13065[0]};
    Full_Adder FA_14162(s14162, c14162, in14162_1, in14162_2, s13063[0]);
    wire[0:0] s14163, in14163_1, in14163_2;
    wire c14163;
    assign in14163_1 = {c13061};
    assign in14163_2 = {c13062};
    Full_Adder FA_14163(s14163, c14163, in14163_1, in14163_2, c13060);
    wire[0:0] s14164, in14164_1, in14164_2;
    wire c14164;
    assign in14164_1 = {c13064};
    assign in14164_2 = {c13065};
    Full_Adder FA_14164(s14164, c14164, in14164_1, in14164_2, c13063);
    wire[0:0] s14165, in14165_1, in14165_2;
    wire c14165;
    assign in14165_1 = {s13067[0]};
    assign in14165_2 = {s13068[0]};
    Full_Adder FA_14165(s14165, c14165, in14165_1, in14165_2, s13066[0]);
    wire[0:0] s14166, in14166_1, in14166_2;
    wire c14166;
    assign in14166_1 = {s13070[0]};
    assign in14166_2 = {s13071[0]};
    Full_Adder FA_14166(s14166, c14166, in14166_1, in14166_2, s13069[0]);
    wire[0:0] s14167, in14167_1, in14167_2;
    wire c14167;
    assign in14167_1 = {c13067};
    assign in14167_2 = {c13068};
    Full_Adder FA_14167(s14167, c14167, in14167_1, in14167_2, c13066);
    wire[0:0] s14168, in14168_1, in14168_2;
    wire c14168;
    assign in14168_1 = {c13070};
    assign in14168_2 = {c13071};
    Full_Adder FA_14168(s14168, c14168, in14168_1, in14168_2, c13069);
    wire[0:0] s14169, in14169_1, in14169_2;
    wire c14169;
    assign in14169_1 = {s13073[0]};
    assign in14169_2 = {s13074[0]};
    Full_Adder FA_14169(s14169, c14169, in14169_1, in14169_2, s13072[0]);
    wire[0:0] s14170, in14170_1, in14170_2;
    wire c14170;
    assign in14170_1 = {s13076[0]};
    assign in14170_2 = {s13077[0]};
    Full_Adder FA_14170(s14170, c14170, in14170_1, in14170_2, s13075[0]);
    wire[0:0] s14171, in14171_1, in14171_2;
    wire c14171;
    assign in14171_1 = {c13073};
    assign in14171_2 = {c13074};
    Full_Adder FA_14171(s14171, c14171, in14171_1, in14171_2, c13072);
    wire[0:0] s14172, in14172_1, in14172_2;
    wire c14172;
    assign in14172_1 = {c13076};
    assign in14172_2 = {c13077};
    Full_Adder FA_14172(s14172, c14172, in14172_1, in14172_2, c13075);
    wire[0:0] s14173, in14173_1, in14173_2;
    wire c14173;
    assign in14173_1 = {s13079[0]};
    assign in14173_2 = {s13080[0]};
    Full_Adder FA_14173(s14173, c14173, in14173_1, in14173_2, s13078[0]);
    wire[0:0] s14174, in14174_1, in14174_2;
    wire c14174;
    assign in14174_1 = {s13082[0]};
    assign in14174_2 = {s13083[0]};
    Full_Adder FA_14174(s14174, c14174, in14174_1, in14174_2, s13081[0]);
    wire[0:0] s14175, in14175_1, in14175_2;
    wire c14175;
    assign in14175_1 = {c13079};
    assign in14175_2 = {c13080};
    Full_Adder FA_14175(s14175, c14175, in14175_1, in14175_2, c13078);
    wire[0:0] s14176, in14176_1, in14176_2;
    wire c14176;
    assign in14176_1 = {c13082};
    assign in14176_2 = {c13083};
    Full_Adder FA_14176(s14176, c14176, in14176_1, in14176_2, c13081);
    wire[0:0] s14177, in14177_1, in14177_2;
    wire c14177;
    assign in14177_1 = {s13085[0]};
    assign in14177_2 = {s13086[0]};
    Full_Adder FA_14177(s14177, c14177, in14177_1, in14177_2, s13084[0]);
    wire[0:0] s14178, in14178_1, in14178_2;
    wire c14178;
    assign in14178_1 = {s13088[0]};
    assign in14178_2 = {s13089[0]};
    Full_Adder FA_14178(s14178, c14178, in14178_1, in14178_2, s13087[0]);
    wire[0:0] s14179, in14179_1, in14179_2;
    wire c14179;
    assign in14179_1 = {c13085};
    assign in14179_2 = {c13086};
    Full_Adder FA_14179(s14179, c14179, in14179_1, in14179_2, c13084);
    wire[0:0] s14180, in14180_1, in14180_2;
    wire c14180;
    assign in14180_1 = {c13088};
    assign in14180_2 = {c13089};
    Full_Adder FA_14180(s14180, c14180, in14180_1, in14180_2, c13087);
    wire[0:0] s14181, in14181_1, in14181_2;
    wire c14181;
    assign in14181_1 = {s13091[0]};
    assign in14181_2 = {s13092[0]};
    Full_Adder FA_14181(s14181, c14181, in14181_1, in14181_2, s13090[0]);
    wire[0:0] s14182, in14182_1, in14182_2;
    wire c14182;
    assign in14182_1 = {s13094[0]};
    assign in14182_2 = {s13095[0]};
    Full_Adder FA_14182(s14182, c14182, in14182_1, in14182_2, s13093[0]);
    wire[0:0] s14183, in14183_1, in14183_2;
    wire c14183;
    assign in14183_1 = {c13091};
    assign in14183_2 = {c13092};
    Full_Adder FA_14183(s14183, c14183, in14183_1, in14183_2, c13090);
    wire[0:0] s14184, in14184_1, in14184_2;
    wire c14184;
    assign in14184_1 = {c13094};
    assign in14184_2 = {c13095};
    Full_Adder FA_14184(s14184, c14184, in14184_1, in14184_2, c13093);
    wire[0:0] s14185, in14185_1, in14185_2;
    wire c14185;
    assign in14185_1 = {s13097[0]};
    assign in14185_2 = {s13098[0]};
    Full_Adder FA_14185(s14185, c14185, in14185_1, in14185_2, s13096[0]);
    wire[0:0] s14186, in14186_1, in14186_2;
    wire c14186;
    assign in14186_1 = {s13100[0]};
    assign in14186_2 = {s13101[0]};
    Full_Adder FA_14186(s14186, c14186, in14186_1, in14186_2, s13099[0]);
    wire[0:0] s14187, in14187_1, in14187_2;
    wire c14187;
    assign in14187_1 = {c13097};
    assign in14187_2 = {c13098};
    Full_Adder FA_14187(s14187, c14187, in14187_1, in14187_2, c13096);
    wire[0:0] s14188, in14188_1, in14188_2;
    wire c14188;
    assign in14188_1 = {c13100};
    assign in14188_2 = {c13101};
    Full_Adder FA_14188(s14188, c14188, in14188_1, in14188_2, c13099);
    wire[0:0] s14189, in14189_1, in14189_2;
    wire c14189;
    assign in14189_1 = {s13103[0]};
    assign in14189_2 = {s13104[0]};
    Full_Adder FA_14189(s14189, c14189, in14189_1, in14189_2, s13102[0]);
    wire[0:0] s14190, in14190_1, in14190_2;
    wire c14190;
    assign in14190_1 = {s13106[0]};
    assign in14190_2 = {s13107[0]};
    Full_Adder FA_14190(s14190, c14190, in14190_1, in14190_2, s13105[0]);
    wire[0:0] s14191, in14191_1, in14191_2;
    wire c14191;
    assign in14191_1 = {c13103};
    assign in14191_2 = {c13104};
    Full_Adder FA_14191(s14191, c14191, in14191_1, in14191_2, c13102);
    wire[0:0] s14192, in14192_1, in14192_2;
    wire c14192;
    assign in14192_1 = {c13106};
    assign in14192_2 = {c13107};
    Full_Adder FA_14192(s14192, c14192, in14192_1, in14192_2, c13105);
    wire[0:0] s14193, in14193_1, in14193_2;
    wire c14193;
    assign in14193_1 = {s13109[0]};
    assign in14193_2 = {s13110[0]};
    Full_Adder FA_14193(s14193, c14193, in14193_1, in14193_2, s13108[0]);
    wire[0:0] s14194, in14194_1, in14194_2;
    wire c14194;
    assign in14194_1 = {s13112[0]};
    assign in14194_2 = {s13113[0]};
    Full_Adder FA_14194(s14194, c14194, in14194_1, in14194_2, s13111[0]);
    wire[0:0] s14195, in14195_1, in14195_2;
    wire c14195;
    assign in14195_1 = {c13109};
    assign in14195_2 = {c13110};
    Full_Adder FA_14195(s14195, c14195, in14195_1, in14195_2, c13108);
    wire[0:0] s14196, in14196_1, in14196_2;
    wire c14196;
    assign in14196_1 = {c13112};
    assign in14196_2 = {c13113};
    Full_Adder FA_14196(s14196, c14196, in14196_1, in14196_2, c13111);
    wire[0:0] s14197, in14197_1, in14197_2;
    wire c14197;
    assign in14197_1 = {s13115[0]};
    assign in14197_2 = {s13116[0]};
    Full_Adder FA_14197(s14197, c14197, in14197_1, in14197_2, s13114[0]);
    wire[0:0] s14198, in14198_1, in14198_2;
    wire c14198;
    assign in14198_1 = {s13118[0]};
    assign in14198_2 = {s13119[0]};
    Full_Adder FA_14198(s14198, c14198, in14198_1, in14198_2, s13117[0]);
    wire[0:0] s14199, in14199_1, in14199_2;
    wire c14199;
    assign in14199_1 = {c13115};
    assign in14199_2 = {c13116};
    Full_Adder FA_14199(s14199, c14199, in14199_1, in14199_2, c13114);
    wire[0:0] s14200, in14200_1, in14200_2;
    wire c14200;
    assign in14200_1 = {c13118};
    assign in14200_2 = {c13119};
    Full_Adder FA_14200(s14200, c14200, in14200_1, in14200_2, c13117);
    wire[0:0] s14201, in14201_1, in14201_2;
    wire c14201;
    assign in14201_1 = {s13121[0]};
    assign in14201_2 = {s13122[0]};
    Full_Adder FA_14201(s14201, c14201, in14201_1, in14201_2, s13120[0]);
    wire[0:0] s14202, in14202_1, in14202_2;
    wire c14202;
    assign in14202_1 = {s13124[0]};
    assign in14202_2 = {s13125[0]};
    Full_Adder FA_14202(s14202, c14202, in14202_1, in14202_2, s13123[0]);
    wire[0:0] s14203, in14203_1, in14203_2;
    wire c14203;
    assign in14203_1 = {c13121};
    assign in14203_2 = {c13122};
    Full_Adder FA_14203(s14203, c14203, in14203_1, in14203_2, c13120);
    wire[0:0] s14204, in14204_1, in14204_2;
    wire c14204;
    assign in14204_1 = {c13124};
    assign in14204_2 = {c13125};
    Full_Adder FA_14204(s14204, c14204, in14204_1, in14204_2, c13123);
    wire[0:0] s14205, in14205_1, in14205_2;
    wire c14205;
    assign in14205_1 = {s13127[0]};
    assign in14205_2 = {s13128[0]};
    Full_Adder FA_14205(s14205, c14205, in14205_1, in14205_2, s13126[0]);
    wire[0:0] s14206, in14206_1, in14206_2;
    wire c14206;
    assign in14206_1 = {s13130[0]};
    assign in14206_2 = {s13131[0]};
    Full_Adder FA_14206(s14206, c14206, in14206_1, in14206_2, s13129[0]);
    wire[0:0] s14207, in14207_1, in14207_2;
    wire c14207;
    assign in14207_1 = {c13127};
    assign in14207_2 = {c13128};
    Full_Adder FA_14207(s14207, c14207, in14207_1, in14207_2, c13126);
    wire[0:0] s14208, in14208_1, in14208_2;
    wire c14208;
    assign in14208_1 = {c13130};
    assign in14208_2 = {c13131};
    Full_Adder FA_14208(s14208, c14208, in14208_1, in14208_2, c13129);
    wire[0:0] s14209, in14209_1, in14209_2;
    wire c14209;
    assign in14209_1 = {s13133[0]};
    assign in14209_2 = {s13134[0]};
    Full_Adder FA_14209(s14209, c14209, in14209_1, in14209_2, s13132[0]);
    wire[0:0] s14210, in14210_1, in14210_2;
    wire c14210;
    assign in14210_1 = {s13136[0]};
    assign in14210_2 = {s13137[0]};
    Full_Adder FA_14210(s14210, c14210, in14210_1, in14210_2, s13135[0]);
    wire[0:0] s14211, in14211_1, in14211_2;
    wire c14211;
    assign in14211_1 = {c13133};
    assign in14211_2 = {c13134};
    Full_Adder FA_14211(s14211, c14211, in14211_1, in14211_2, c13132);
    wire[0:0] s14212, in14212_1, in14212_2;
    wire c14212;
    assign in14212_1 = {c13136};
    assign in14212_2 = {c13137};
    Full_Adder FA_14212(s14212, c14212, in14212_1, in14212_2, c13135);
    wire[0:0] s14213, in14213_1, in14213_2;
    wire c14213;
    assign in14213_1 = {s13139[0]};
    assign in14213_2 = {s13140[0]};
    Full_Adder FA_14213(s14213, c14213, in14213_1, in14213_2, s13138[0]);
    wire[0:0] s14214, in14214_1, in14214_2;
    wire c14214;
    assign in14214_1 = {s13142[0]};
    assign in14214_2 = {s13143[0]};
    Full_Adder FA_14214(s14214, c14214, in14214_1, in14214_2, s13141[0]);
    wire[0:0] s14215, in14215_1, in14215_2;
    wire c14215;
    assign in14215_1 = {c13139};
    assign in14215_2 = {c13140};
    Full_Adder FA_14215(s14215, c14215, in14215_1, in14215_2, c13138);
    wire[0:0] s14216, in14216_1, in14216_2;
    wire c14216;
    assign in14216_1 = {c13142};
    assign in14216_2 = {c13143};
    Full_Adder FA_14216(s14216, c14216, in14216_1, in14216_2, c13141);
    wire[0:0] s14217, in14217_1, in14217_2;
    wire c14217;
    assign in14217_1 = {s13145[0]};
    assign in14217_2 = {s13146[0]};
    Full_Adder FA_14217(s14217, c14217, in14217_1, in14217_2, s13144[0]);
    wire[0:0] s14218, in14218_1, in14218_2;
    wire c14218;
    assign in14218_1 = {s13148[0]};
    assign in14218_2 = {s13149[0]};
    Full_Adder FA_14218(s14218, c14218, in14218_1, in14218_2, s13147[0]);
    wire[0:0] s14219, in14219_1, in14219_2;
    wire c14219;
    assign in14219_1 = {c13145};
    assign in14219_2 = {c13146};
    Full_Adder FA_14219(s14219, c14219, in14219_1, in14219_2, c13144);
    wire[0:0] s14220, in14220_1, in14220_2;
    wire c14220;
    assign in14220_1 = {c13148};
    assign in14220_2 = {c13149};
    Full_Adder FA_14220(s14220, c14220, in14220_1, in14220_2, c13147);
    wire[0:0] s14221, in14221_1, in14221_2;
    wire c14221;
    assign in14221_1 = {s13151[0]};
    assign in14221_2 = {s13152[0]};
    Full_Adder FA_14221(s14221, c14221, in14221_1, in14221_2, s13150[0]);
    wire[0:0] s14222, in14222_1, in14222_2;
    wire c14222;
    assign in14222_1 = {s13154[0]};
    assign in14222_2 = {s13155[0]};
    Full_Adder FA_14222(s14222, c14222, in14222_1, in14222_2, s13153[0]);
    wire[0:0] s14223, in14223_1, in14223_2;
    wire c14223;
    assign in14223_1 = {c13151};
    assign in14223_2 = {c13152};
    Full_Adder FA_14223(s14223, c14223, in14223_1, in14223_2, c13150);
    wire[0:0] s14224, in14224_1, in14224_2;
    wire c14224;
    assign in14224_1 = {c13154};
    assign in14224_2 = {c13155};
    Full_Adder FA_14224(s14224, c14224, in14224_1, in14224_2, c13153);
    wire[0:0] s14225, in14225_1, in14225_2;
    wire c14225;
    assign in14225_1 = {s13157[0]};
    assign in14225_2 = {s13158[0]};
    Full_Adder FA_14225(s14225, c14225, in14225_1, in14225_2, s13156[0]);
    wire[0:0] s14226, in14226_1, in14226_2;
    wire c14226;
    assign in14226_1 = {s13160[0]};
    assign in14226_2 = {s13161[0]};
    Full_Adder FA_14226(s14226, c14226, in14226_1, in14226_2, s13159[0]);
    wire[0:0] s14227, in14227_1, in14227_2;
    wire c14227;
    assign in14227_1 = {c13157};
    assign in14227_2 = {c13158};
    Full_Adder FA_14227(s14227, c14227, in14227_1, in14227_2, c13156);
    wire[0:0] s14228, in14228_1, in14228_2;
    wire c14228;
    assign in14228_1 = {c13160};
    assign in14228_2 = {c13161};
    Full_Adder FA_14228(s14228, c14228, in14228_1, in14228_2, c13159);
    wire[0:0] s14229, in14229_1, in14229_2;
    wire c14229;
    assign in14229_1 = {s13163[0]};
    assign in14229_2 = {s13164[0]};
    Full_Adder FA_14229(s14229, c14229, in14229_1, in14229_2, s13162[0]);
    wire[0:0] s14230, in14230_1, in14230_2;
    wire c14230;
    assign in14230_1 = {s13166[0]};
    assign in14230_2 = {s13167[0]};
    Full_Adder FA_14230(s14230, c14230, in14230_1, in14230_2, s13165[0]);
    wire[0:0] s14231, in14231_1, in14231_2;
    wire c14231;
    assign in14231_1 = {c13163};
    assign in14231_2 = {c13164};
    Full_Adder FA_14231(s14231, c14231, in14231_1, in14231_2, c13162);
    wire[0:0] s14232, in14232_1, in14232_2;
    wire c14232;
    assign in14232_1 = {c13166};
    assign in14232_2 = {c13167};
    Full_Adder FA_14232(s14232, c14232, in14232_1, in14232_2, c13165);
    wire[0:0] s14233, in14233_1, in14233_2;
    wire c14233;
    assign in14233_1 = {s13169[0]};
    assign in14233_2 = {s13170[0]};
    Full_Adder FA_14233(s14233, c14233, in14233_1, in14233_2, s13168[0]);
    wire[0:0] s14234, in14234_1, in14234_2;
    wire c14234;
    assign in14234_1 = {s13172[0]};
    assign in14234_2 = {s13173[0]};
    Full_Adder FA_14234(s14234, c14234, in14234_1, in14234_2, s13171[0]);
    wire[0:0] s14235, in14235_1, in14235_2;
    wire c14235;
    assign in14235_1 = {c13169};
    assign in14235_2 = {c13170};
    Full_Adder FA_14235(s14235, c14235, in14235_1, in14235_2, c13168);
    wire[0:0] s14236, in14236_1, in14236_2;
    wire c14236;
    assign in14236_1 = {c13172};
    assign in14236_2 = {c13173};
    Full_Adder FA_14236(s14236, c14236, in14236_1, in14236_2, c13171);
    wire[0:0] s14237, in14237_1, in14237_2;
    wire c14237;
    assign in14237_1 = {s13175[0]};
    assign in14237_2 = {s13176[0]};
    Full_Adder FA_14237(s14237, c14237, in14237_1, in14237_2, s13174[0]);
    wire[0:0] s14238, in14238_1, in14238_2;
    wire c14238;
    assign in14238_1 = {s13178[0]};
    assign in14238_2 = {s13179[0]};
    Full_Adder FA_14238(s14238, c14238, in14238_1, in14238_2, s13177[0]);
    wire[0:0] s14239, in14239_1, in14239_2;
    wire c14239;
    assign in14239_1 = {c13175};
    assign in14239_2 = {c13176};
    Full_Adder FA_14239(s14239, c14239, in14239_1, in14239_2, c13174);
    wire[0:0] s14240, in14240_1, in14240_2;
    wire c14240;
    assign in14240_1 = {c13178};
    assign in14240_2 = {c13179};
    Full_Adder FA_14240(s14240, c14240, in14240_1, in14240_2, c13177);
    wire[0:0] s14241, in14241_1, in14241_2;
    wire c14241;
    assign in14241_1 = {s13181[0]};
    assign in14241_2 = {s13182[0]};
    Full_Adder FA_14241(s14241, c14241, in14241_1, in14241_2, s13180[0]);
    wire[0:0] s14242, in14242_1, in14242_2;
    wire c14242;
    assign in14242_1 = {s13184[0]};
    assign in14242_2 = {s13185[0]};
    Full_Adder FA_14242(s14242, c14242, in14242_1, in14242_2, s13183[0]);
    wire[0:0] s14243, in14243_1, in14243_2;
    wire c14243;
    assign in14243_1 = {c13181};
    assign in14243_2 = {c13182};
    Full_Adder FA_14243(s14243, c14243, in14243_1, in14243_2, c13180);
    wire[0:0] s14244, in14244_1, in14244_2;
    wire c14244;
    assign in14244_1 = {c13184};
    assign in14244_2 = {c13185};
    Full_Adder FA_14244(s14244, c14244, in14244_1, in14244_2, c13183);
    wire[0:0] s14245, in14245_1, in14245_2;
    wire c14245;
    assign in14245_1 = {s13187[0]};
    assign in14245_2 = {s13188[0]};
    Full_Adder FA_14245(s14245, c14245, in14245_1, in14245_2, s13186[0]);
    wire[0:0] s14246, in14246_1, in14246_2;
    wire c14246;
    assign in14246_1 = {s13190[0]};
    assign in14246_2 = {s13191[0]};
    Full_Adder FA_14246(s14246, c14246, in14246_1, in14246_2, s13189[0]);
    wire[0:0] s14247, in14247_1, in14247_2;
    wire c14247;
    assign in14247_1 = {c13187};
    assign in14247_2 = {c13188};
    Full_Adder FA_14247(s14247, c14247, in14247_1, in14247_2, c13186);
    wire[0:0] s14248, in14248_1, in14248_2;
    wire c14248;
    assign in14248_1 = {c13190};
    assign in14248_2 = {c13191};
    Full_Adder FA_14248(s14248, c14248, in14248_1, in14248_2, c13189);
    wire[0:0] s14249, in14249_1, in14249_2;
    wire c14249;
    assign in14249_1 = {s13193[0]};
    assign in14249_2 = {s13194[0]};
    Full_Adder FA_14249(s14249, c14249, in14249_1, in14249_2, s13192[0]);
    wire[0:0] s14250, in14250_1, in14250_2;
    wire c14250;
    assign in14250_1 = {s13196[0]};
    assign in14250_2 = {s13197[0]};
    Full_Adder FA_14250(s14250, c14250, in14250_1, in14250_2, s13195[0]);
    wire[0:0] s14251, in14251_1, in14251_2;
    wire c14251;
    assign in14251_1 = {c13193};
    assign in14251_2 = {c13194};
    Full_Adder FA_14251(s14251, c14251, in14251_1, in14251_2, c13192);
    wire[0:0] s14252, in14252_1, in14252_2;
    wire c14252;
    assign in14252_1 = {c13196};
    assign in14252_2 = {c13197};
    Full_Adder FA_14252(s14252, c14252, in14252_1, in14252_2, c13195);
    wire[0:0] s14253, in14253_1, in14253_2;
    wire c14253;
    assign in14253_1 = {s13199[0]};
    assign in14253_2 = {s13200[0]};
    Full_Adder FA_14253(s14253, c14253, in14253_1, in14253_2, s13198[0]);
    wire[0:0] s14254, in14254_1, in14254_2;
    wire c14254;
    assign in14254_1 = {s13202[0]};
    assign in14254_2 = {s13203[0]};
    Full_Adder FA_14254(s14254, c14254, in14254_1, in14254_2, s13201[0]);
    wire[0:0] s14255, in14255_1, in14255_2;
    wire c14255;
    assign in14255_1 = {c13199};
    assign in14255_2 = {c13200};
    Full_Adder FA_14255(s14255, c14255, in14255_1, in14255_2, c13198);
    wire[0:0] s14256, in14256_1, in14256_2;
    wire c14256;
    assign in14256_1 = {c13202};
    assign in14256_2 = {c13203};
    Full_Adder FA_14256(s14256, c14256, in14256_1, in14256_2, c13201);
    wire[0:0] s14257, in14257_1, in14257_2;
    wire c14257;
    assign in14257_1 = {s13205[0]};
    assign in14257_2 = {s13206[0]};
    Full_Adder FA_14257(s14257, c14257, in14257_1, in14257_2, s13204[0]);
    wire[0:0] s14258, in14258_1, in14258_2;
    wire c14258;
    assign in14258_1 = {s13208[0]};
    assign in14258_2 = {s13209[0]};
    Full_Adder FA_14258(s14258, c14258, in14258_1, in14258_2, s13207[0]);
    wire[0:0] s14259, in14259_1, in14259_2;
    wire c14259;
    assign in14259_1 = {c13205};
    assign in14259_2 = {c13206};
    Full_Adder FA_14259(s14259, c14259, in14259_1, in14259_2, c13204);
    wire[0:0] s14260, in14260_1, in14260_2;
    wire c14260;
    assign in14260_1 = {c13208};
    assign in14260_2 = {c13209};
    Full_Adder FA_14260(s14260, c14260, in14260_1, in14260_2, c13207);
    wire[0:0] s14261, in14261_1, in14261_2;
    wire c14261;
    assign in14261_1 = {s13211[0]};
    assign in14261_2 = {s13212[0]};
    Full_Adder FA_14261(s14261, c14261, in14261_1, in14261_2, s13210[0]);
    wire[0:0] s14262, in14262_1, in14262_2;
    wire c14262;
    assign in14262_1 = {s13214[0]};
    assign in14262_2 = {s13215[0]};
    Full_Adder FA_14262(s14262, c14262, in14262_1, in14262_2, s13213[0]);
    wire[0:0] s14263, in14263_1, in14263_2;
    wire c14263;
    assign in14263_1 = {c13211};
    assign in14263_2 = {c13212};
    Full_Adder FA_14263(s14263, c14263, in14263_1, in14263_2, c13210);
    wire[0:0] s14264, in14264_1, in14264_2;
    wire c14264;
    assign in14264_1 = {c13214};
    assign in14264_2 = {c13215};
    Full_Adder FA_14264(s14264, c14264, in14264_1, in14264_2, c13213);
    wire[0:0] s14265, in14265_1, in14265_2;
    wire c14265;
    assign in14265_1 = {s13217[0]};
    assign in14265_2 = {s13218[0]};
    Full_Adder FA_14265(s14265, c14265, in14265_1, in14265_2, s13216[0]);
    wire[0:0] s14266, in14266_1, in14266_2;
    wire c14266;
    assign in14266_1 = {s13220[0]};
    assign in14266_2 = {s13221[0]};
    Full_Adder FA_14266(s14266, c14266, in14266_1, in14266_2, s13219[0]);
    wire[0:0] s14267, in14267_1, in14267_2;
    wire c14267;
    assign in14267_1 = {c13217};
    assign in14267_2 = {c13218};
    Full_Adder FA_14267(s14267, c14267, in14267_1, in14267_2, c13216);
    wire[0:0] s14268, in14268_1, in14268_2;
    wire c14268;
    assign in14268_1 = {c13220};
    assign in14268_2 = {c13221};
    Full_Adder FA_14268(s14268, c14268, in14268_1, in14268_2, c13219);
    wire[0:0] s14269, in14269_1, in14269_2;
    wire c14269;
    assign in14269_1 = {s13223[0]};
    assign in14269_2 = {s13224[0]};
    Full_Adder FA_14269(s14269, c14269, in14269_1, in14269_2, s13222[0]);
    wire[0:0] s14270, in14270_1, in14270_2;
    wire c14270;
    assign in14270_1 = {s13226[0]};
    assign in14270_2 = {s13227[0]};
    Full_Adder FA_14270(s14270, c14270, in14270_1, in14270_2, s13225[0]);
    wire[0:0] s14271, in14271_1, in14271_2;
    wire c14271;
    assign in14271_1 = {c13223};
    assign in14271_2 = {c13224};
    Full_Adder FA_14271(s14271, c14271, in14271_1, in14271_2, c13222);
    wire[0:0] s14272, in14272_1, in14272_2;
    wire c14272;
    assign in14272_1 = {c13226};
    assign in14272_2 = {c13227};
    Full_Adder FA_14272(s14272, c14272, in14272_1, in14272_2, c13225);
    wire[0:0] s14273, in14273_1, in14273_2;
    wire c14273;
    assign in14273_1 = {s13229[0]};
    assign in14273_2 = {s13230[0]};
    Full_Adder FA_14273(s14273, c14273, in14273_1, in14273_2, s13228[0]);
    wire[0:0] s14274, in14274_1, in14274_2;
    wire c14274;
    assign in14274_1 = {s13232[0]};
    assign in14274_2 = {s13233[0]};
    Full_Adder FA_14274(s14274, c14274, in14274_1, in14274_2, s13231[0]);
    wire[0:0] s14275, in14275_1, in14275_2;
    wire c14275;
    assign in14275_1 = {c13229};
    assign in14275_2 = {c13230};
    Full_Adder FA_14275(s14275, c14275, in14275_1, in14275_2, c13228);
    wire[0:0] s14276, in14276_1, in14276_2;
    wire c14276;
    assign in14276_1 = {c13232};
    assign in14276_2 = {c13233};
    Full_Adder FA_14276(s14276, c14276, in14276_1, in14276_2, c13231);
    wire[0:0] s14277, in14277_1, in14277_2;
    wire c14277;
    assign in14277_1 = {s13235[0]};
    assign in14277_2 = {s13236[0]};
    Full_Adder FA_14277(s14277, c14277, in14277_1, in14277_2, s13234[0]);
    wire[0:0] s14278, in14278_1, in14278_2;
    wire c14278;
    assign in14278_1 = {s13238[0]};
    assign in14278_2 = {s13239[0]};
    Full_Adder FA_14278(s14278, c14278, in14278_1, in14278_2, s13237[0]);
    wire[0:0] s14279, in14279_1, in14279_2;
    wire c14279;
    assign in14279_1 = {c13235};
    assign in14279_2 = {c13236};
    Full_Adder FA_14279(s14279, c14279, in14279_1, in14279_2, c13234);
    wire[0:0] s14280, in14280_1, in14280_2;
    wire c14280;
    assign in14280_1 = {c13238};
    assign in14280_2 = {c13239};
    Full_Adder FA_14280(s14280, c14280, in14280_1, in14280_2, c13237);
    wire[0:0] s14281, in14281_1, in14281_2;
    wire c14281;
    assign in14281_1 = {s13241[0]};
    assign in14281_2 = {s13242[0]};
    Full_Adder FA_14281(s14281, c14281, in14281_1, in14281_2, s13240[0]);
    wire[0:0] s14282, in14282_1, in14282_2;
    wire c14282;
    assign in14282_1 = {s13244[0]};
    assign in14282_2 = {s13245[0]};
    Full_Adder FA_14282(s14282, c14282, in14282_1, in14282_2, s13243[0]);
    wire[0:0] s14283, in14283_1, in14283_2;
    wire c14283;
    assign in14283_1 = {c13241};
    assign in14283_2 = {c13242};
    Full_Adder FA_14283(s14283, c14283, in14283_1, in14283_2, c13240);
    wire[0:0] s14284, in14284_1, in14284_2;
    wire c14284;
    assign in14284_1 = {c13244};
    assign in14284_2 = {c13245};
    Full_Adder FA_14284(s14284, c14284, in14284_1, in14284_2, c13243);
    wire[0:0] s14285, in14285_1, in14285_2;
    wire c14285;
    assign in14285_1 = {s13247[0]};
    assign in14285_2 = {s13248[0]};
    Full_Adder FA_14285(s14285, c14285, in14285_1, in14285_2, s13246[0]);
    wire[0:0] s14286, in14286_1, in14286_2;
    wire c14286;
    assign in14286_1 = {s13250[0]};
    assign in14286_2 = {s13251[0]};
    Full_Adder FA_14286(s14286, c14286, in14286_1, in14286_2, s13249[0]);
    wire[0:0] s14287, in14287_1, in14287_2;
    wire c14287;
    assign in14287_1 = {c13247};
    assign in14287_2 = {c13248};
    Full_Adder FA_14287(s14287, c14287, in14287_1, in14287_2, c13246);
    wire[0:0] s14288, in14288_1, in14288_2;
    wire c14288;
    assign in14288_1 = {c13250};
    assign in14288_2 = {c13251};
    Full_Adder FA_14288(s14288, c14288, in14288_1, in14288_2, c13249);
    wire[0:0] s14289, in14289_1, in14289_2;
    wire c14289;
    assign in14289_1 = {s13253[0]};
    assign in14289_2 = {s13254[0]};
    Full_Adder FA_14289(s14289, c14289, in14289_1, in14289_2, s13252[0]);
    wire[0:0] s14290, in14290_1, in14290_2;
    wire c14290;
    assign in14290_1 = {s13256[0]};
    assign in14290_2 = {s13257[0]};
    Full_Adder FA_14290(s14290, c14290, in14290_1, in14290_2, s13255[0]);
    wire[0:0] s14291, in14291_1, in14291_2;
    wire c14291;
    assign in14291_1 = {c13253};
    assign in14291_2 = {c13254};
    Full_Adder FA_14291(s14291, c14291, in14291_1, in14291_2, c13252);
    wire[0:0] s14292, in14292_1, in14292_2;
    wire c14292;
    assign in14292_1 = {c13256};
    assign in14292_2 = {c13257};
    Full_Adder FA_14292(s14292, c14292, in14292_1, in14292_2, c13255);
    wire[0:0] s14293, in14293_1, in14293_2;
    wire c14293;
    assign in14293_1 = {s13259[0]};
    assign in14293_2 = {s13260[0]};
    Full_Adder FA_14293(s14293, c14293, in14293_1, in14293_2, s13258[0]);
    wire[0:0] s14294, in14294_1, in14294_2;
    wire c14294;
    assign in14294_1 = {s13262[0]};
    assign in14294_2 = {s13263[0]};
    Full_Adder FA_14294(s14294, c14294, in14294_1, in14294_2, s13261[0]);
    wire[0:0] s14295, in14295_1, in14295_2;
    wire c14295;
    assign in14295_1 = {c13259};
    assign in14295_2 = {c13260};
    Full_Adder FA_14295(s14295, c14295, in14295_1, in14295_2, c13258);
    wire[0:0] s14296, in14296_1, in14296_2;
    wire c14296;
    assign in14296_1 = {c13262};
    assign in14296_2 = {c13263};
    Full_Adder FA_14296(s14296, c14296, in14296_1, in14296_2, c13261);
    wire[0:0] s14297, in14297_1, in14297_2;
    wire c14297;
    assign in14297_1 = {s13265[0]};
    assign in14297_2 = {s13266[0]};
    Full_Adder FA_14297(s14297, c14297, in14297_1, in14297_2, s13264[0]);
    wire[0:0] s14298, in14298_1, in14298_2;
    wire c14298;
    assign in14298_1 = {s13268[0]};
    assign in14298_2 = {s13269[0]};
    Full_Adder FA_14298(s14298, c14298, in14298_1, in14298_2, s13267[0]);
    wire[0:0] s14299, in14299_1, in14299_2;
    wire c14299;
    assign in14299_1 = {c13265};
    assign in14299_2 = {c13266};
    Full_Adder FA_14299(s14299, c14299, in14299_1, in14299_2, c13264);
    wire[0:0] s14300, in14300_1, in14300_2;
    wire c14300;
    assign in14300_1 = {c13268};
    assign in14300_2 = {c13269};
    Full_Adder FA_14300(s14300, c14300, in14300_1, in14300_2, c13267);
    wire[0:0] s14301, in14301_1, in14301_2;
    wire c14301;
    assign in14301_1 = {s13271[0]};
    assign in14301_2 = {s13272[0]};
    Full_Adder FA_14301(s14301, c14301, in14301_1, in14301_2, s13270[0]);
    wire[0:0] s14302, in14302_1, in14302_2;
    wire c14302;
    assign in14302_1 = {s13274[0]};
    assign in14302_2 = {s13275[0]};
    Full_Adder FA_14302(s14302, c14302, in14302_1, in14302_2, s13273[0]);
    wire[0:0] s14303, in14303_1, in14303_2;
    wire c14303;
    assign in14303_1 = {c13271};
    assign in14303_2 = {c13272};
    Full_Adder FA_14303(s14303, c14303, in14303_1, in14303_2, c13270);
    wire[0:0] s14304, in14304_1, in14304_2;
    wire c14304;
    assign in14304_1 = {c13274};
    assign in14304_2 = {c13275};
    Full_Adder FA_14304(s14304, c14304, in14304_1, in14304_2, c13273);
    wire[0:0] s14305, in14305_1, in14305_2;
    wire c14305;
    assign in14305_1 = {s13277[0]};
    assign in14305_2 = {s13278[0]};
    Full_Adder FA_14305(s14305, c14305, in14305_1, in14305_2, s13276[0]);
    wire[0:0] s14306, in14306_1, in14306_2;
    wire c14306;
    assign in14306_1 = {s13280[0]};
    assign in14306_2 = {s13281[0]};
    Full_Adder FA_14306(s14306, c14306, in14306_1, in14306_2, s13279[0]);
    wire[0:0] s14307, in14307_1, in14307_2;
    wire c14307;
    assign in14307_1 = {c13277};
    assign in14307_2 = {c13278};
    Full_Adder FA_14307(s14307, c14307, in14307_1, in14307_2, c13276);
    wire[0:0] s14308, in14308_1, in14308_2;
    wire c14308;
    assign in14308_1 = {c13280};
    assign in14308_2 = {c13281};
    Full_Adder FA_14308(s14308, c14308, in14308_1, in14308_2, c13279);
    wire[0:0] s14309, in14309_1, in14309_2;
    wire c14309;
    assign in14309_1 = {s13283[0]};
    assign in14309_2 = {s13284[0]};
    Full_Adder FA_14309(s14309, c14309, in14309_1, in14309_2, s13282[0]);
    wire[0:0] s14310, in14310_1, in14310_2;
    wire c14310;
    assign in14310_1 = {s13286[0]};
    assign in14310_2 = {s13287[0]};
    Full_Adder FA_14310(s14310, c14310, in14310_1, in14310_2, s13285[0]);
    wire[0:0] s14311, in14311_1, in14311_2;
    wire c14311;
    assign in14311_1 = {c13283};
    assign in14311_2 = {c13284};
    Full_Adder FA_14311(s14311, c14311, in14311_1, in14311_2, c13282);
    wire[0:0] s14312, in14312_1, in14312_2;
    wire c14312;
    assign in14312_1 = {c13286};
    assign in14312_2 = {c13287};
    Full_Adder FA_14312(s14312, c14312, in14312_1, in14312_2, c13285);
    wire[0:0] s14313, in14313_1, in14313_2;
    wire c14313;
    assign in14313_1 = {s13289[0]};
    assign in14313_2 = {s13290[0]};
    Full_Adder FA_14313(s14313, c14313, in14313_1, in14313_2, s13288[0]);
    wire[0:0] s14314, in14314_1, in14314_2;
    wire c14314;
    assign in14314_1 = {s13292[0]};
    assign in14314_2 = {s13293[0]};
    Full_Adder FA_14314(s14314, c14314, in14314_1, in14314_2, s13291[0]);
    wire[0:0] s14315, in14315_1, in14315_2;
    wire c14315;
    assign in14315_1 = {c13289};
    assign in14315_2 = {c13290};
    Full_Adder FA_14315(s14315, c14315, in14315_1, in14315_2, c13288);
    wire[0:0] s14316, in14316_1, in14316_2;
    wire c14316;
    assign in14316_1 = {c13292};
    assign in14316_2 = {c13293};
    Full_Adder FA_14316(s14316, c14316, in14316_1, in14316_2, c13291);
    wire[0:0] s14317, in14317_1, in14317_2;
    wire c14317;
    assign in14317_1 = {s13295[0]};
    assign in14317_2 = {s13296[0]};
    Full_Adder FA_14317(s14317, c14317, in14317_1, in14317_2, s13294[0]);
    wire[0:0] s14318, in14318_1, in14318_2;
    wire c14318;
    assign in14318_1 = {s13298[0]};
    assign in14318_2 = {s13299[0]};
    Full_Adder FA_14318(s14318, c14318, in14318_1, in14318_2, s13297[0]);
    wire[0:0] s14319, in14319_1, in14319_2;
    wire c14319;
    assign in14319_1 = {c13295};
    assign in14319_2 = {c13296};
    Full_Adder FA_14319(s14319, c14319, in14319_1, in14319_2, c13294);
    wire[0:0] s14320, in14320_1, in14320_2;
    wire c14320;
    assign in14320_1 = {c13298};
    assign in14320_2 = {c13299};
    Full_Adder FA_14320(s14320, c14320, in14320_1, in14320_2, c13297);
    wire[0:0] s14321, in14321_1, in14321_2;
    wire c14321;
    assign in14321_1 = {s13301[0]};
    assign in14321_2 = {s13302[0]};
    Full_Adder FA_14321(s14321, c14321, in14321_1, in14321_2, s13300[0]);
    wire[0:0] s14322, in14322_1, in14322_2;
    wire c14322;
    assign in14322_1 = {s13304[0]};
    assign in14322_2 = {s13305[0]};
    Full_Adder FA_14322(s14322, c14322, in14322_1, in14322_2, s13303[0]);
    wire[0:0] s14323, in14323_1, in14323_2;
    wire c14323;
    assign in14323_1 = {c13301};
    assign in14323_2 = {c13302};
    Full_Adder FA_14323(s14323, c14323, in14323_1, in14323_2, c13300);
    wire[0:0] s14324, in14324_1, in14324_2;
    wire c14324;
    assign in14324_1 = {c13304};
    assign in14324_2 = {c13305};
    Full_Adder FA_14324(s14324, c14324, in14324_1, in14324_2, c13303);
    wire[0:0] s14325, in14325_1, in14325_2;
    wire c14325;
    assign in14325_1 = {s13307[0]};
    assign in14325_2 = {s13308[0]};
    Full_Adder FA_14325(s14325, c14325, in14325_1, in14325_2, s13306[0]);
    wire[0:0] s14326, in14326_1, in14326_2;
    wire c14326;
    assign in14326_1 = {s13310[0]};
    assign in14326_2 = {s13311[0]};
    Full_Adder FA_14326(s14326, c14326, in14326_1, in14326_2, s13309[0]);
    wire[0:0] s14327, in14327_1, in14327_2;
    wire c14327;
    assign in14327_1 = {c13307};
    assign in14327_2 = {c13308};
    Full_Adder FA_14327(s14327, c14327, in14327_1, in14327_2, c13306);
    wire[0:0] s14328, in14328_1, in14328_2;
    wire c14328;
    assign in14328_1 = {c13310};
    assign in14328_2 = {c13311};
    Full_Adder FA_14328(s14328, c14328, in14328_1, in14328_2, c13309);
    wire[0:0] s14329, in14329_1, in14329_2;
    wire c14329;
    assign in14329_1 = {s13313[0]};
    assign in14329_2 = {s13314[0]};
    Full_Adder FA_14329(s14329, c14329, in14329_1, in14329_2, s13312[0]);
    wire[0:0] s14330, in14330_1, in14330_2;
    wire c14330;
    assign in14330_1 = {s13316[0]};
    assign in14330_2 = {s13317[0]};
    Full_Adder FA_14330(s14330, c14330, in14330_1, in14330_2, s13315[0]);
    wire[0:0] s14331, in14331_1, in14331_2;
    wire c14331;
    assign in14331_1 = {c13313};
    assign in14331_2 = {c13314};
    Full_Adder FA_14331(s14331, c14331, in14331_1, in14331_2, c13312);
    wire[0:0] s14332, in14332_1, in14332_2;
    wire c14332;
    assign in14332_1 = {c13316};
    assign in14332_2 = {c13317};
    Full_Adder FA_14332(s14332, c14332, in14332_1, in14332_2, c13315);
    wire[0:0] s14333, in14333_1, in14333_2;
    wire c14333;
    assign in14333_1 = {s13319[0]};
    assign in14333_2 = {s13320[0]};
    Full_Adder FA_14333(s14333, c14333, in14333_1, in14333_2, s13318[0]);
    wire[0:0] s14334, in14334_1, in14334_2;
    wire c14334;
    assign in14334_1 = {s13322[0]};
    assign in14334_2 = {s13323[0]};
    Full_Adder FA_14334(s14334, c14334, in14334_1, in14334_2, s13321[0]);
    wire[0:0] s14335, in14335_1, in14335_2;
    wire c14335;
    assign in14335_1 = {c13319};
    assign in14335_2 = {c13320};
    Full_Adder FA_14335(s14335, c14335, in14335_1, in14335_2, c13318);
    wire[0:0] s14336, in14336_1, in14336_2;
    wire c14336;
    assign in14336_1 = {c13322};
    assign in14336_2 = {c13323};
    Full_Adder FA_14336(s14336, c14336, in14336_1, in14336_2, c13321);
    wire[0:0] s14337, in14337_1, in14337_2;
    wire c14337;
    assign in14337_1 = {s13325[0]};
    assign in14337_2 = {s13326[0]};
    Full_Adder FA_14337(s14337, c14337, in14337_1, in14337_2, s13324[0]);
    wire[0:0] s14338, in14338_1, in14338_2;
    wire c14338;
    assign in14338_1 = {s13328[0]};
    assign in14338_2 = {s13329[0]};
    Full_Adder FA_14338(s14338, c14338, in14338_1, in14338_2, s13327[0]);
    wire[0:0] s14339, in14339_1, in14339_2;
    wire c14339;
    assign in14339_1 = {c13325};
    assign in14339_2 = {c13326};
    Full_Adder FA_14339(s14339, c14339, in14339_1, in14339_2, c13324);
    wire[0:0] s14340, in14340_1, in14340_2;
    wire c14340;
    assign in14340_1 = {c13328};
    assign in14340_2 = {c13329};
    Full_Adder FA_14340(s14340, c14340, in14340_1, in14340_2, c13327);
    wire[0:0] s14341, in14341_1, in14341_2;
    wire c14341;
    assign in14341_1 = {s13331[0]};
    assign in14341_2 = {s13332[0]};
    Full_Adder FA_14341(s14341, c14341, in14341_1, in14341_2, s13330[0]);
    wire[0:0] s14342, in14342_1, in14342_2;
    wire c14342;
    assign in14342_1 = {s13334[0]};
    assign in14342_2 = {s13335[0]};
    Full_Adder FA_14342(s14342, c14342, in14342_1, in14342_2, s13333[0]);
    wire[0:0] s14343, in14343_1, in14343_2;
    wire c14343;
    assign in14343_1 = {c13331};
    assign in14343_2 = {c13332};
    Full_Adder FA_14343(s14343, c14343, in14343_1, in14343_2, c13330);
    wire[0:0] s14344, in14344_1, in14344_2;
    wire c14344;
    assign in14344_1 = {c13334};
    assign in14344_2 = {c13335};
    Full_Adder FA_14344(s14344, c14344, in14344_1, in14344_2, c13333);
    wire[0:0] s14345, in14345_1, in14345_2;
    wire c14345;
    assign in14345_1 = {s13337[0]};
    assign in14345_2 = {s13338[0]};
    Full_Adder FA_14345(s14345, c14345, in14345_1, in14345_2, s13336[0]);
    wire[0:0] s14346, in14346_1, in14346_2;
    wire c14346;
    assign in14346_1 = {s13340[0]};
    assign in14346_2 = {s13341[0]};
    Full_Adder FA_14346(s14346, c14346, in14346_1, in14346_2, s13339[0]);
    wire[0:0] s14347, in14347_1, in14347_2;
    wire c14347;
    assign in14347_1 = {c13337};
    assign in14347_2 = {c13338};
    Full_Adder FA_14347(s14347, c14347, in14347_1, in14347_2, c13336);
    wire[0:0] s14348, in14348_1, in14348_2;
    wire c14348;
    assign in14348_1 = {c13340};
    assign in14348_2 = {c13341};
    Full_Adder FA_14348(s14348, c14348, in14348_1, in14348_2, c13339);
    wire[0:0] s14349, in14349_1, in14349_2;
    wire c14349;
    assign in14349_1 = {s13343[0]};
    assign in14349_2 = {s13344[0]};
    Full_Adder FA_14349(s14349, c14349, in14349_1, in14349_2, s13342[0]);
    wire[0:0] s14350, in14350_1, in14350_2;
    wire c14350;
    assign in14350_1 = {s13346[0]};
    assign in14350_2 = {s13347[0]};
    Full_Adder FA_14350(s14350, c14350, in14350_1, in14350_2, s13345[0]);
    wire[0:0] s14351, in14351_1, in14351_2;
    wire c14351;
    assign in14351_1 = {c13343};
    assign in14351_2 = {c13344};
    Full_Adder FA_14351(s14351, c14351, in14351_1, in14351_2, c13342);
    wire[0:0] s14352, in14352_1, in14352_2;
    wire c14352;
    assign in14352_1 = {c13346};
    assign in14352_2 = {c13347};
    Full_Adder FA_14352(s14352, c14352, in14352_1, in14352_2, c13345);
    wire[0:0] s14353, in14353_1, in14353_2;
    wire c14353;
    assign in14353_1 = {s13349[0]};
    assign in14353_2 = {s13350[0]};
    Full_Adder FA_14353(s14353, c14353, in14353_1, in14353_2, s13348[0]);
    wire[0:0] s14354, in14354_1, in14354_2;
    wire c14354;
    assign in14354_1 = {s13352[0]};
    assign in14354_2 = {s13353[0]};
    Full_Adder FA_14354(s14354, c14354, in14354_1, in14354_2, s13351[0]);
    wire[0:0] s14355, in14355_1, in14355_2;
    wire c14355;
    assign in14355_1 = {c13349};
    assign in14355_2 = {c13350};
    Full_Adder FA_14355(s14355, c14355, in14355_1, in14355_2, c13348);
    wire[0:0] s14356, in14356_1, in14356_2;
    wire c14356;
    assign in14356_1 = {c13352};
    assign in14356_2 = {c13353};
    Full_Adder FA_14356(s14356, c14356, in14356_1, in14356_2, c13351);
    wire[0:0] s14357, in14357_1, in14357_2;
    wire c14357;
    assign in14357_1 = {s13355[0]};
    assign in14357_2 = {s13356[0]};
    Full_Adder FA_14357(s14357, c14357, in14357_1, in14357_2, s13354[0]);
    wire[0:0] s14358, in14358_1, in14358_2;
    wire c14358;
    assign in14358_1 = {s13358[0]};
    assign in14358_2 = {s13359[0]};
    Full_Adder FA_14358(s14358, c14358, in14358_1, in14358_2, s13357[0]);
    wire[0:0] s14359, in14359_1, in14359_2;
    wire c14359;
    assign in14359_1 = {c13355};
    assign in14359_2 = {c13356};
    Full_Adder FA_14359(s14359, c14359, in14359_1, in14359_2, c13354);
    wire[0:0] s14360, in14360_1, in14360_2;
    wire c14360;
    assign in14360_1 = {c13358};
    assign in14360_2 = {c13359};
    Full_Adder FA_14360(s14360, c14360, in14360_1, in14360_2, c13357);
    wire[0:0] s14361, in14361_1, in14361_2;
    wire c14361;
    assign in14361_1 = {s13361[0]};
    assign in14361_2 = {s13362[0]};
    Full_Adder FA_14361(s14361, c14361, in14361_1, in14361_2, s13360[0]);
    wire[0:0] s14362, in14362_1, in14362_2;
    wire c14362;
    assign in14362_1 = {s13364[0]};
    assign in14362_2 = {s13365[0]};
    Full_Adder FA_14362(s14362, c14362, in14362_1, in14362_2, s13363[0]);
    wire[0:0] s14363, in14363_1, in14363_2;
    wire c14363;
    assign in14363_1 = {c13361};
    assign in14363_2 = {c13362};
    Full_Adder FA_14363(s14363, c14363, in14363_1, in14363_2, c13360);
    wire[0:0] s14364, in14364_1, in14364_2;
    wire c14364;
    assign in14364_1 = {c13364};
    assign in14364_2 = {c13365};
    Full_Adder FA_14364(s14364, c14364, in14364_1, in14364_2, c13363);
    wire[0:0] s14365, in14365_1, in14365_2;
    wire c14365;
    assign in14365_1 = {s13367[0]};
    assign in14365_2 = {s13368[0]};
    Full_Adder FA_14365(s14365, c14365, in14365_1, in14365_2, s13366[0]);
    wire[0:0] s14366, in14366_1, in14366_2;
    wire c14366;
    assign in14366_1 = {s13370[0]};
    assign in14366_2 = {s13371[0]};
    Full_Adder FA_14366(s14366, c14366, in14366_1, in14366_2, s13369[0]);
    wire[0:0] s14367, in14367_1, in14367_2;
    wire c14367;
    assign in14367_1 = {c13367};
    assign in14367_2 = {c13368};
    Full_Adder FA_14367(s14367, c14367, in14367_1, in14367_2, c13366);
    wire[0:0] s14368, in14368_1, in14368_2;
    wire c14368;
    assign in14368_1 = {c13370};
    assign in14368_2 = {c13371};
    Full_Adder FA_14368(s14368, c14368, in14368_1, in14368_2, c13369);
    wire[0:0] s14369, in14369_1, in14369_2;
    wire c14369;
    assign in14369_1 = {s13373[0]};
    assign in14369_2 = {s13374[0]};
    Full_Adder FA_14369(s14369, c14369, in14369_1, in14369_2, s13372[0]);
    wire[0:0] s14370, in14370_1, in14370_2;
    wire c14370;
    assign in14370_1 = {s13376[0]};
    assign in14370_2 = {s13377[0]};
    Full_Adder FA_14370(s14370, c14370, in14370_1, in14370_2, s13375[0]);
    wire[0:0] s14371, in14371_1, in14371_2;
    wire c14371;
    assign in14371_1 = {c13373};
    assign in14371_2 = {c13374};
    Full_Adder FA_14371(s14371, c14371, in14371_1, in14371_2, c13372);
    wire[0:0] s14372, in14372_1, in14372_2;
    wire c14372;
    assign in14372_1 = {c13376};
    assign in14372_2 = {c13377};
    Full_Adder FA_14372(s14372, c14372, in14372_1, in14372_2, c13375);
    wire[0:0] s14373, in14373_1, in14373_2;
    wire c14373;
    assign in14373_1 = {s13379[0]};
    assign in14373_2 = {s13380[0]};
    Full_Adder FA_14373(s14373, c14373, in14373_1, in14373_2, s13378[0]);
    wire[0:0] s14374, in14374_1, in14374_2;
    wire c14374;
    assign in14374_1 = {s13382[0]};
    assign in14374_2 = {s13383[0]};
    Full_Adder FA_14374(s14374, c14374, in14374_1, in14374_2, s13381[0]);
    wire[0:0] s14375, in14375_1, in14375_2;
    wire c14375;
    assign in14375_1 = {c13379};
    assign in14375_2 = {c13380};
    Full_Adder FA_14375(s14375, c14375, in14375_1, in14375_2, c13378);
    wire[0:0] s14376, in14376_1, in14376_2;
    wire c14376;
    assign in14376_1 = {c13382};
    assign in14376_2 = {c13383};
    Full_Adder FA_14376(s14376, c14376, in14376_1, in14376_2, c13381);
    wire[0:0] s14377, in14377_1, in14377_2;
    wire c14377;
    assign in14377_1 = {s13385[0]};
    assign in14377_2 = {s13386[0]};
    Full_Adder FA_14377(s14377, c14377, in14377_1, in14377_2, s13384[0]);
    wire[0:0] s14378, in14378_1, in14378_2;
    wire c14378;
    assign in14378_1 = {s13388[0]};
    assign in14378_2 = {s13389[0]};
    Full_Adder FA_14378(s14378, c14378, in14378_1, in14378_2, s13387[0]);
    wire[0:0] s14379, in14379_1, in14379_2;
    wire c14379;
    assign in14379_1 = {c13385};
    assign in14379_2 = {c13386};
    Full_Adder FA_14379(s14379, c14379, in14379_1, in14379_2, c13384);
    wire[0:0] s14380, in14380_1, in14380_2;
    wire c14380;
    assign in14380_1 = {c13388};
    assign in14380_2 = {c13389};
    Full_Adder FA_14380(s14380, c14380, in14380_1, in14380_2, c13387);
    wire[0:0] s14381, in14381_1, in14381_2;
    wire c14381;
    assign in14381_1 = {s13391[0]};
    assign in14381_2 = {s13392[0]};
    Full_Adder FA_14381(s14381, c14381, in14381_1, in14381_2, s13390[0]);
    wire[0:0] s14382, in14382_1, in14382_2;
    wire c14382;
    assign in14382_1 = {s13394[0]};
    assign in14382_2 = {s13395[0]};
    Full_Adder FA_14382(s14382, c14382, in14382_1, in14382_2, s13393[0]);
    wire[0:0] s14383, in14383_1, in14383_2;
    wire c14383;
    assign in14383_1 = {c13391};
    assign in14383_2 = {c13392};
    Full_Adder FA_14383(s14383, c14383, in14383_1, in14383_2, c13390);
    wire[0:0] s14384, in14384_1, in14384_2;
    wire c14384;
    assign in14384_1 = {c13394};
    assign in14384_2 = {c13395};
    Full_Adder FA_14384(s14384, c14384, in14384_1, in14384_2, c13393);
    wire[0:0] s14385, in14385_1, in14385_2;
    wire c14385;
    assign in14385_1 = {s13397[0]};
    assign in14385_2 = {s13398[0]};
    Full_Adder FA_14385(s14385, c14385, in14385_1, in14385_2, s13396[0]);
    wire[0:0] s14386, in14386_1, in14386_2;
    wire c14386;
    assign in14386_1 = {s13400[0]};
    assign in14386_2 = {s13401[0]};
    Full_Adder FA_14386(s14386, c14386, in14386_1, in14386_2, s13399[0]);
    wire[0:0] s14387, in14387_1, in14387_2;
    wire c14387;
    assign in14387_1 = {c13397};
    assign in14387_2 = {c13398};
    Full_Adder FA_14387(s14387, c14387, in14387_1, in14387_2, c13396);
    wire[0:0] s14388, in14388_1, in14388_2;
    wire c14388;
    assign in14388_1 = {c13400};
    assign in14388_2 = {c13401};
    Full_Adder FA_14388(s14388, c14388, in14388_1, in14388_2, c13399);
    wire[0:0] s14389, in14389_1, in14389_2;
    wire c14389;
    assign in14389_1 = {s13403[0]};
    assign in14389_2 = {s13404[0]};
    Full_Adder FA_14389(s14389, c14389, in14389_1, in14389_2, s13402[0]);
    wire[0:0] s14390, in14390_1, in14390_2;
    wire c14390;
    assign in14390_1 = {s13406[0]};
    assign in14390_2 = {s13407[0]};
    Full_Adder FA_14390(s14390, c14390, in14390_1, in14390_2, s13405[0]);
    wire[0:0] s14391, in14391_1, in14391_2;
    wire c14391;
    assign in14391_1 = {c13403};
    assign in14391_2 = {c13404};
    Full_Adder FA_14391(s14391, c14391, in14391_1, in14391_2, c13402);
    wire[0:0] s14392, in14392_1, in14392_2;
    wire c14392;
    assign in14392_1 = {c13406};
    assign in14392_2 = {c13407};
    Full_Adder FA_14392(s14392, c14392, in14392_1, in14392_2, c13405);
    wire[0:0] s14393, in14393_1, in14393_2;
    wire c14393;
    assign in14393_1 = {s13409[0]};
    assign in14393_2 = {s13410[0]};
    Full_Adder FA_14393(s14393, c14393, in14393_1, in14393_2, s13408[0]);
    wire[0:0] s14394, in14394_1, in14394_2;
    wire c14394;
    assign in14394_1 = {s13412[0]};
    assign in14394_2 = {s13413[0]};
    Full_Adder FA_14394(s14394, c14394, in14394_1, in14394_2, s13411[0]);
    wire[0:0] s14395, in14395_1, in14395_2;
    wire c14395;
    assign in14395_1 = {c13409};
    assign in14395_2 = {c13410};
    Full_Adder FA_14395(s14395, c14395, in14395_1, in14395_2, c13408);
    wire[0:0] s14396, in14396_1, in14396_2;
    wire c14396;
    assign in14396_1 = {c13412};
    assign in14396_2 = {c13413};
    Full_Adder FA_14396(s14396, c14396, in14396_1, in14396_2, c13411);
    wire[0:0] s14397, in14397_1, in14397_2;
    wire c14397;
    assign in14397_1 = {s13415[0]};
    assign in14397_2 = {s13416[0]};
    Full_Adder FA_14397(s14397, c14397, in14397_1, in14397_2, s13414[0]);
    wire[0:0] s14398, in14398_1, in14398_2;
    wire c14398;
    assign in14398_1 = {s13418[0]};
    assign in14398_2 = {s13419[0]};
    Full_Adder FA_14398(s14398, c14398, in14398_1, in14398_2, s13417[0]);
    wire[0:0] s14399, in14399_1, in14399_2;
    wire c14399;
    assign in14399_1 = {c13415};
    assign in14399_2 = {c13416};
    Full_Adder FA_14399(s14399, c14399, in14399_1, in14399_2, c13414);
    wire[0:0] s14400, in14400_1, in14400_2;
    wire c14400;
    assign in14400_1 = {c13418};
    assign in14400_2 = {c13419};
    Full_Adder FA_14400(s14400, c14400, in14400_1, in14400_2, c13417);
    wire[0:0] s14401, in14401_1, in14401_2;
    wire c14401;
    assign in14401_1 = {s13421[0]};
    assign in14401_2 = {s13422[0]};
    Full_Adder FA_14401(s14401, c14401, in14401_1, in14401_2, s13420[0]);
    wire[0:0] s14402, in14402_1, in14402_2;
    wire c14402;
    assign in14402_1 = {s13424[0]};
    assign in14402_2 = {s13425[0]};
    Full_Adder FA_14402(s14402, c14402, in14402_1, in14402_2, s13423[0]);
    wire[0:0] s14403, in14403_1, in14403_2;
    wire c14403;
    assign in14403_1 = {c13421};
    assign in14403_2 = {c13422};
    Full_Adder FA_14403(s14403, c14403, in14403_1, in14403_2, c13420);
    wire[0:0] s14404, in14404_1, in14404_2;
    wire c14404;
    assign in14404_1 = {c13424};
    assign in14404_2 = {c13425};
    Full_Adder FA_14404(s14404, c14404, in14404_1, in14404_2, c13423);
    wire[0:0] s14405, in14405_1, in14405_2;
    wire c14405;
    assign in14405_1 = {s13427[0]};
    assign in14405_2 = {s13428[0]};
    Full_Adder FA_14405(s14405, c14405, in14405_1, in14405_2, s13426[0]);
    wire[0:0] s14406, in14406_1, in14406_2;
    wire c14406;
    assign in14406_1 = {s13430[0]};
    assign in14406_2 = {s13431[0]};
    Full_Adder FA_14406(s14406, c14406, in14406_1, in14406_2, s13429[0]);
    wire[0:0] s14407, in14407_1, in14407_2;
    wire c14407;
    assign in14407_1 = {c13427};
    assign in14407_2 = {c13428};
    Full_Adder FA_14407(s14407, c14407, in14407_1, in14407_2, c13426);
    wire[0:0] s14408, in14408_1, in14408_2;
    wire c14408;
    assign in14408_1 = {c13430};
    assign in14408_2 = {c13431};
    Full_Adder FA_14408(s14408, c14408, in14408_1, in14408_2, c13429);
    wire[0:0] s14409, in14409_1, in14409_2;
    wire c14409;
    assign in14409_1 = {s13433[0]};
    assign in14409_2 = {s13434[0]};
    Full_Adder FA_14409(s14409, c14409, in14409_1, in14409_2, s13432[0]);
    wire[0:0] s14410, in14410_1, in14410_2;
    wire c14410;
    assign in14410_1 = {s13436[0]};
    assign in14410_2 = {s13437[0]};
    Full_Adder FA_14410(s14410, c14410, in14410_1, in14410_2, s13435[0]);
    wire[0:0] s14411, in14411_1, in14411_2;
    wire c14411;
    assign in14411_1 = {c13433};
    assign in14411_2 = {c13434};
    Full_Adder FA_14411(s14411, c14411, in14411_1, in14411_2, c13432);
    wire[0:0] s14412, in14412_1, in14412_2;
    wire c14412;
    assign in14412_1 = {c13436};
    assign in14412_2 = {c13437};
    Full_Adder FA_14412(s14412, c14412, in14412_1, in14412_2, c13435);
    wire[0:0] s14413, in14413_1, in14413_2;
    wire c14413;
    assign in14413_1 = {s13439[0]};
    assign in14413_2 = {s13440[0]};
    Full_Adder FA_14413(s14413, c14413, in14413_1, in14413_2, s13438[0]);
    wire[0:0] s14414, in14414_1, in14414_2;
    wire c14414;
    assign in14414_1 = {s13442[0]};
    assign in14414_2 = {s13443[0]};
    Full_Adder FA_14414(s14414, c14414, in14414_1, in14414_2, s13441[0]);
    wire[0:0] s14415, in14415_1, in14415_2;
    wire c14415;
    assign in14415_1 = {c13439};
    assign in14415_2 = {c13440};
    Full_Adder FA_14415(s14415, c14415, in14415_1, in14415_2, c13438);
    wire[0:0] s14416, in14416_1, in14416_2;
    wire c14416;
    assign in14416_1 = {c13442};
    assign in14416_2 = {c13443};
    Full_Adder FA_14416(s14416, c14416, in14416_1, in14416_2, c13441);
    wire[0:0] s14417, in14417_1, in14417_2;
    wire c14417;
    assign in14417_1 = {s13445[0]};
    assign in14417_2 = {s13446[0]};
    Full_Adder FA_14417(s14417, c14417, in14417_1, in14417_2, s13444[0]);
    wire[0:0] s14418, in14418_1, in14418_2;
    wire c14418;
    assign in14418_1 = {s13448[0]};
    assign in14418_2 = {s13449[0]};
    Full_Adder FA_14418(s14418, c14418, in14418_1, in14418_2, s13447[0]);
    wire[0:0] s14419, in14419_1, in14419_2;
    wire c14419;
    assign in14419_1 = {c13445};
    assign in14419_2 = {c13446};
    Full_Adder FA_14419(s14419, c14419, in14419_1, in14419_2, c13444);
    wire[0:0] s14420, in14420_1, in14420_2;
    wire c14420;
    assign in14420_1 = {c13448};
    assign in14420_2 = {c13449};
    Full_Adder FA_14420(s14420, c14420, in14420_1, in14420_2, c13447);
    wire[0:0] s14421, in14421_1, in14421_2;
    wire c14421;
    assign in14421_1 = {s13451[0]};
    assign in14421_2 = {s13452[0]};
    Full_Adder FA_14421(s14421, c14421, in14421_1, in14421_2, s13450[0]);
    wire[0:0] s14422, in14422_1, in14422_2;
    wire c14422;
    assign in14422_1 = {s13454[0]};
    assign in14422_2 = {s13455[0]};
    Full_Adder FA_14422(s14422, c14422, in14422_1, in14422_2, s13453[0]);
    wire[0:0] s14423, in14423_1, in14423_2;
    wire c14423;
    assign in14423_1 = {c13451};
    assign in14423_2 = {c13452};
    Full_Adder FA_14423(s14423, c14423, in14423_1, in14423_2, c13450);
    wire[0:0] s14424, in14424_1, in14424_2;
    wire c14424;
    assign in14424_1 = {c13454};
    assign in14424_2 = {c13455};
    Full_Adder FA_14424(s14424, c14424, in14424_1, in14424_2, c13453);
    wire[0:0] s14425, in14425_1, in14425_2;
    wire c14425;
    assign in14425_1 = {s13457[0]};
    assign in14425_2 = {s13458[0]};
    Full_Adder FA_14425(s14425, c14425, in14425_1, in14425_2, s13456[0]);
    wire[0:0] s14426, in14426_1, in14426_2;
    wire c14426;
    assign in14426_1 = {s13460[0]};
    assign in14426_2 = {s13461[0]};
    Full_Adder FA_14426(s14426, c14426, in14426_1, in14426_2, s13459[0]);
    wire[0:0] s14427, in14427_1, in14427_2;
    wire c14427;
    assign in14427_1 = {c13457};
    assign in14427_2 = {c13458};
    Full_Adder FA_14427(s14427, c14427, in14427_1, in14427_2, c13456);
    wire[0:0] s14428, in14428_1, in14428_2;
    wire c14428;
    assign in14428_1 = {c13460};
    assign in14428_2 = {c13461};
    Full_Adder FA_14428(s14428, c14428, in14428_1, in14428_2, c13459);
    wire[0:0] s14429, in14429_1, in14429_2;
    wire c14429;
    assign in14429_1 = {s13463[0]};
    assign in14429_2 = {s13464[0]};
    Full_Adder FA_14429(s14429, c14429, in14429_1, in14429_2, s13462[0]);
    wire[0:0] s14430, in14430_1, in14430_2;
    wire c14430;
    assign in14430_1 = {s13466[0]};
    assign in14430_2 = {s13467[0]};
    Full_Adder FA_14430(s14430, c14430, in14430_1, in14430_2, s13465[0]);
    wire[0:0] s14431, in14431_1, in14431_2;
    wire c14431;
    assign in14431_1 = {c13463};
    assign in14431_2 = {c13464};
    Full_Adder FA_14431(s14431, c14431, in14431_1, in14431_2, c13462);
    wire[0:0] s14432, in14432_1, in14432_2;
    wire c14432;
    assign in14432_1 = {c13466};
    assign in14432_2 = {c13467};
    Full_Adder FA_14432(s14432, c14432, in14432_1, in14432_2, c13465);
    wire[0:0] s14433, in14433_1, in14433_2;
    wire c14433;
    assign in14433_1 = {s13469[0]};
    assign in14433_2 = {s13470[0]};
    Full_Adder FA_14433(s14433, c14433, in14433_1, in14433_2, s13468[0]);
    wire[0:0] s14434, in14434_1, in14434_2;
    wire c14434;
    assign in14434_1 = {s13472[0]};
    assign in14434_2 = {s13473[0]};
    Full_Adder FA_14434(s14434, c14434, in14434_1, in14434_2, s13471[0]);
    wire[0:0] s14435, in14435_1, in14435_2;
    wire c14435;
    assign in14435_1 = {c13469};
    assign in14435_2 = {c13470};
    Full_Adder FA_14435(s14435, c14435, in14435_1, in14435_2, c13468);
    wire[0:0] s14436, in14436_1, in14436_2;
    wire c14436;
    assign in14436_1 = {c13472};
    assign in14436_2 = {c13473};
    Full_Adder FA_14436(s14436, c14436, in14436_1, in14436_2, c13471);
    wire[0:0] s14437, in14437_1, in14437_2;
    wire c14437;
    assign in14437_1 = {s13475[0]};
    assign in14437_2 = {s13476[0]};
    Full_Adder FA_14437(s14437, c14437, in14437_1, in14437_2, s13474[0]);
    wire[0:0] s14438, in14438_1, in14438_2;
    wire c14438;
    assign in14438_1 = {s13478[0]};
    assign in14438_2 = {s13479[0]};
    Full_Adder FA_14438(s14438, c14438, in14438_1, in14438_2, s13477[0]);
    wire[0:0] s14439, in14439_1, in14439_2;
    wire c14439;
    assign in14439_1 = {c13475};
    assign in14439_2 = {c13476};
    Full_Adder FA_14439(s14439, c14439, in14439_1, in14439_2, c13474);
    wire[0:0] s14440, in14440_1, in14440_2;
    wire c14440;
    assign in14440_1 = {c13478};
    assign in14440_2 = {c13479};
    Full_Adder FA_14440(s14440, c14440, in14440_1, in14440_2, c13477);
    wire[0:0] s14441, in14441_1, in14441_2;
    wire c14441;
    assign in14441_1 = {s13481[0]};
    assign in14441_2 = {s13482[0]};
    Full_Adder FA_14441(s14441, c14441, in14441_1, in14441_2, s13480[0]);
    wire[0:0] s14442, in14442_1, in14442_2;
    wire c14442;
    assign in14442_1 = {s13484[0]};
    assign in14442_2 = {s13485[0]};
    Full_Adder FA_14442(s14442, c14442, in14442_1, in14442_2, s13483[0]);
    wire[0:0] s14443, in14443_1, in14443_2;
    wire c14443;
    assign in14443_1 = {c13481};
    assign in14443_2 = {c13482};
    Full_Adder FA_14443(s14443, c14443, in14443_1, in14443_2, c13480);
    wire[0:0] s14444, in14444_1, in14444_2;
    wire c14444;
    assign in14444_1 = {c13484};
    assign in14444_2 = {c13485};
    Full_Adder FA_14444(s14444, c14444, in14444_1, in14444_2, c13483);
    wire[0:0] s14445, in14445_1, in14445_2;
    wire c14445;
    assign in14445_1 = {s13487[0]};
    assign in14445_2 = {s13488[0]};
    Full_Adder FA_14445(s14445, c14445, in14445_1, in14445_2, s13486[0]);
    wire[0:0] s14446, in14446_1, in14446_2;
    wire c14446;
    assign in14446_1 = {s13490[0]};
    assign in14446_2 = {s13491[0]};
    Full_Adder FA_14446(s14446, c14446, in14446_1, in14446_2, s13489[0]);
    wire[0:0] s14447, in14447_1, in14447_2;
    wire c14447;
    assign in14447_1 = {c13487};
    assign in14447_2 = {c13488};
    Full_Adder FA_14447(s14447, c14447, in14447_1, in14447_2, c13486);
    wire[0:0] s14448, in14448_1, in14448_2;
    wire c14448;
    assign in14448_1 = {c13490};
    assign in14448_2 = {c13491};
    Full_Adder FA_14448(s14448, c14448, in14448_1, in14448_2, c13489);
    wire[0:0] s14449, in14449_1, in14449_2;
    wire c14449;
    assign in14449_1 = {s13493[0]};
    assign in14449_2 = {s13494[0]};
    Full_Adder FA_14449(s14449, c14449, in14449_1, in14449_2, s13492[0]);
    wire[0:0] s14450, in14450_1, in14450_2;
    wire c14450;
    assign in14450_1 = {s13496[0]};
    assign in14450_2 = {s13497[0]};
    Full_Adder FA_14450(s14450, c14450, in14450_1, in14450_2, s13495[0]);
    wire[0:0] s14451, in14451_1, in14451_2;
    wire c14451;
    assign in14451_1 = {c13493};
    assign in14451_2 = {c13494};
    Full_Adder FA_14451(s14451, c14451, in14451_1, in14451_2, c13492);
    wire[0:0] s14452, in14452_1, in14452_2;
    wire c14452;
    assign in14452_1 = {c13496};
    assign in14452_2 = {c13497};
    Full_Adder FA_14452(s14452, c14452, in14452_1, in14452_2, c13495);
    wire[0:0] s14453, in14453_1, in14453_2;
    wire c14453;
    assign in14453_1 = {s13499[0]};
    assign in14453_2 = {s13500[0]};
    Full_Adder FA_14453(s14453, c14453, in14453_1, in14453_2, s13498[0]);
    wire[0:0] s14454, in14454_1, in14454_2;
    wire c14454;
    assign in14454_1 = {s13502[0]};
    assign in14454_2 = {s13503[0]};
    Full_Adder FA_14454(s14454, c14454, in14454_1, in14454_2, s13501[0]);
    wire[0:0] s14455, in14455_1, in14455_2;
    wire c14455;
    assign in14455_1 = {c13499};
    assign in14455_2 = {c13500};
    Full_Adder FA_14455(s14455, c14455, in14455_1, in14455_2, c13498);
    wire[0:0] s14456, in14456_1, in14456_2;
    wire c14456;
    assign in14456_1 = {c13502};
    assign in14456_2 = {c13503};
    Full_Adder FA_14456(s14456, c14456, in14456_1, in14456_2, c13501);
    wire[0:0] s14457, in14457_1, in14457_2;
    wire c14457;
    assign in14457_1 = {s13505[0]};
    assign in14457_2 = {s13506[0]};
    Full_Adder FA_14457(s14457, c14457, in14457_1, in14457_2, s13504[0]);
    wire[0:0] s14458, in14458_1, in14458_2;
    wire c14458;
    assign in14458_1 = {s13508[0]};
    assign in14458_2 = {s13509[0]};
    Full_Adder FA_14458(s14458, c14458, in14458_1, in14458_2, s13507[0]);
    wire[0:0] s14459, in14459_1, in14459_2;
    wire c14459;
    assign in14459_1 = {c13505};
    assign in14459_2 = {c13506};
    Full_Adder FA_14459(s14459, c14459, in14459_1, in14459_2, c13504);
    wire[0:0] s14460, in14460_1, in14460_2;
    wire c14460;
    assign in14460_1 = {c13508};
    assign in14460_2 = {c13509};
    Full_Adder FA_14460(s14460, c14460, in14460_1, in14460_2, c13507);
    wire[0:0] s14461, in14461_1, in14461_2;
    wire c14461;
    assign in14461_1 = {s13511[0]};
    assign in14461_2 = {s13512[0]};
    Full_Adder FA_14461(s14461, c14461, in14461_1, in14461_2, s13510[0]);
    wire[0:0] s14462, in14462_1, in14462_2;
    wire c14462;
    assign in14462_1 = {s13514[0]};
    assign in14462_2 = {s13515[0]};
    Full_Adder FA_14462(s14462, c14462, in14462_1, in14462_2, s13513[0]);
    wire[0:0] s14463, in14463_1, in14463_2;
    wire c14463;
    assign in14463_1 = {c13511};
    assign in14463_2 = {c13512};
    Full_Adder FA_14463(s14463, c14463, in14463_1, in14463_2, c13510);
    wire[0:0] s14464, in14464_1, in14464_2;
    wire c14464;
    assign in14464_1 = {c13514};
    assign in14464_2 = {c13515};
    Full_Adder FA_14464(s14464, c14464, in14464_1, in14464_2, c13513);
    wire[0:0] s14465, in14465_1, in14465_2;
    wire c14465;
    assign in14465_1 = {s13517[0]};
    assign in14465_2 = {s13518[0]};
    Full_Adder FA_14465(s14465, c14465, in14465_1, in14465_2, s13516[0]);
    wire[0:0] s14466, in14466_1, in14466_2;
    wire c14466;
    assign in14466_1 = {s13520[0]};
    assign in14466_2 = {s13521[0]};
    Full_Adder FA_14466(s14466, c14466, in14466_1, in14466_2, s13519[0]);
    wire[0:0] s14467, in14467_1, in14467_2;
    wire c14467;
    assign in14467_1 = {c13517};
    assign in14467_2 = {c13518};
    Full_Adder FA_14467(s14467, c14467, in14467_1, in14467_2, c13516);
    wire[0:0] s14468, in14468_1, in14468_2;
    wire c14468;
    assign in14468_1 = {c13520};
    assign in14468_2 = {c13521};
    Full_Adder FA_14468(s14468, c14468, in14468_1, in14468_2, c13519);
    wire[0:0] s14469, in14469_1, in14469_2;
    wire c14469;
    assign in14469_1 = {s13523[0]};
    assign in14469_2 = {s13524[0]};
    Full_Adder FA_14469(s14469, c14469, in14469_1, in14469_2, s13522[0]);
    wire[0:0] s14470, in14470_1, in14470_2;
    wire c14470;
    assign in14470_1 = {s13526[0]};
    assign in14470_2 = {s13527[0]};
    Full_Adder FA_14470(s14470, c14470, in14470_1, in14470_2, s13525[0]);
    wire[0:0] s14471, in14471_1, in14471_2;
    wire c14471;
    assign in14471_1 = {c13523};
    assign in14471_2 = {c13524};
    Full_Adder FA_14471(s14471, c14471, in14471_1, in14471_2, c13522);
    wire[0:0] s14472, in14472_1, in14472_2;
    wire c14472;
    assign in14472_1 = {c13526};
    assign in14472_2 = {c13527};
    Full_Adder FA_14472(s14472, c14472, in14472_1, in14472_2, c13525);
    wire[0:0] s14473, in14473_1, in14473_2;
    wire c14473;
    assign in14473_1 = {s13529[0]};
    assign in14473_2 = {s13530[0]};
    Full_Adder FA_14473(s14473, c14473, in14473_1, in14473_2, s13528[0]);
    wire[0:0] s14474, in14474_1, in14474_2;
    wire c14474;
    assign in14474_1 = {s13532[0]};
    assign in14474_2 = {s13533[0]};
    Full_Adder FA_14474(s14474, c14474, in14474_1, in14474_2, s13531[0]);
    wire[0:0] s14475, in14475_1, in14475_2;
    wire c14475;
    assign in14475_1 = {c13529};
    assign in14475_2 = {c13530};
    Full_Adder FA_14475(s14475, c14475, in14475_1, in14475_2, c13528);
    wire[0:0] s14476, in14476_1, in14476_2;
    wire c14476;
    assign in14476_1 = {c13532};
    assign in14476_2 = {c13533};
    Full_Adder FA_14476(s14476, c14476, in14476_1, in14476_2, c13531);
    wire[0:0] s14477, in14477_1, in14477_2;
    wire c14477;
    assign in14477_1 = {s13535[0]};
    assign in14477_2 = {s13536[0]};
    Full_Adder FA_14477(s14477, c14477, in14477_1, in14477_2, s13534[0]);
    wire[0:0] s14478, in14478_1, in14478_2;
    wire c14478;
    assign in14478_1 = {s13538[0]};
    assign in14478_2 = {s13539[0]};
    Full_Adder FA_14478(s14478, c14478, in14478_1, in14478_2, s13537[0]);
    wire[0:0] s14479, in14479_1, in14479_2;
    wire c14479;
    assign in14479_1 = {c13535};
    assign in14479_2 = {c13536};
    Full_Adder FA_14479(s14479, c14479, in14479_1, in14479_2, c13534);
    wire[0:0] s14480, in14480_1, in14480_2;
    wire c14480;
    assign in14480_1 = {c13538};
    assign in14480_2 = {c13539};
    Full_Adder FA_14480(s14480, c14480, in14480_1, in14480_2, c13537);
    wire[0:0] s14481, in14481_1, in14481_2;
    wire c14481;
    assign in14481_1 = {s13541[0]};
    assign in14481_2 = {s13542[0]};
    Full_Adder FA_14481(s14481, c14481, in14481_1, in14481_2, s13540[0]);
    wire[0:0] s14482, in14482_1, in14482_2;
    wire c14482;
    assign in14482_1 = {s13544[0]};
    assign in14482_2 = {s13545[0]};
    Full_Adder FA_14482(s14482, c14482, in14482_1, in14482_2, s13543[0]);
    wire[0:0] s14483, in14483_1, in14483_2;
    wire c14483;
    assign in14483_1 = {c13541};
    assign in14483_2 = {c13542};
    Full_Adder FA_14483(s14483, c14483, in14483_1, in14483_2, c13540);
    wire[0:0] s14484, in14484_1, in14484_2;
    wire c14484;
    assign in14484_1 = {c13544};
    assign in14484_2 = {c13545};
    Full_Adder FA_14484(s14484, c14484, in14484_1, in14484_2, c13543);
    wire[0:0] s14485, in14485_1, in14485_2;
    wire c14485;
    assign in14485_1 = {s13547[0]};
    assign in14485_2 = {s13548[0]};
    Full_Adder FA_14485(s14485, c14485, in14485_1, in14485_2, s13546[0]);
    wire[0:0] s14486, in14486_1, in14486_2;
    wire c14486;
    assign in14486_1 = {s13550[0]};
    assign in14486_2 = {s13551[0]};
    Full_Adder FA_14486(s14486, c14486, in14486_1, in14486_2, s13549[0]);
    wire[0:0] s14487, in14487_1, in14487_2;
    wire c14487;
    assign in14487_1 = {c13547};
    assign in14487_2 = {c13548};
    Full_Adder FA_14487(s14487, c14487, in14487_1, in14487_2, c13546);
    wire[0:0] s14488, in14488_1, in14488_2;
    wire c14488;
    assign in14488_1 = {c13550};
    assign in14488_2 = {c13551};
    Full_Adder FA_14488(s14488, c14488, in14488_1, in14488_2, c13549);
    wire[0:0] s14489, in14489_1, in14489_2;
    wire c14489;
    assign in14489_1 = {s13553[0]};
    assign in14489_2 = {s13554[0]};
    Full_Adder FA_14489(s14489, c14489, in14489_1, in14489_2, s13552[0]);
    wire[0:0] s14490, in14490_1, in14490_2;
    wire c14490;
    assign in14490_1 = {s13556[0]};
    assign in14490_2 = {s13557[0]};
    Full_Adder FA_14490(s14490, c14490, in14490_1, in14490_2, s13555[0]);
    wire[0:0] s14491, in14491_1, in14491_2;
    wire c14491;
    assign in14491_1 = {c13552};
    assign in14491_2 = {c13553};
    Full_Adder FA_14491(s14491, c14491, in14491_1, in14491_2, pp127[112]);
    wire[0:0] s14492, in14492_1, in14492_2;
    wire c14492;
    assign in14492_1 = {c13555};
    assign in14492_2 = {c13556};
    Full_Adder FA_14492(s14492, c14492, in14492_1, in14492_2, c13554);
    wire[0:0] s14493, in14493_1, in14493_2;
    wire c14493;
    assign in14493_1 = {s13558[0]};
    assign in14493_2 = {s13559[0]};
    Full_Adder FA_14493(s14493, c14493, in14493_1, in14493_2, c13557);
    wire[0:0] s14494, in14494_1, in14494_2;
    wire c14494;
    assign in14494_1 = {s13561[0]};
    assign in14494_2 = {s13562[0]};
    Full_Adder FA_14494(s14494, c14494, in14494_1, in14494_2, s13560[0]);
    wire[0:0] s14495, in14495_1, in14495_2;
    wire c14495;
    assign in14495_1 = {pp126[114]};
    assign in14495_2 = {pp127[113]};
    Full_Adder FA_14495(s14495, c14495, in14495_1, in14495_2, pp125[115]);
    wire[0:0] s14496, in14496_1, in14496_2;
    wire c14496;
    assign in14496_1 = {c13559};
    assign in14496_2 = {c13560};
    Full_Adder FA_14496(s14496, c14496, in14496_1, in14496_2, c13558);
    wire[0:0] s14497, in14497_1, in14497_2;
    wire c14497;
    assign in14497_1 = {c13562};
    assign in14497_2 = {s13563[0]};
    Full_Adder FA_14497(s14497, c14497, in14497_1, in14497_2, c13561);
    wire[0:0] s14498, in14498_1, in14498_2;
    wire c14498;
    assign in14498_1 = {s13565[0]};
    assign in14498_2 = {s13566[0]};
    Full_Adder FA_14498(s14498, c14498, in14498_1, in14498_2, s13564[0]);
    wire[0:0] s14499, in14499_1, in14499_2;
    wire c14499;
    assign in14499_1 = {pp124[117]};
    assign in14499_2 = {pp125[116]};
    Full_Adder FA_14499(s14499, c14499, in14499_1, in14499_2, pp123[118]);
    wire[0:0] s14500, in14500_1, in14500_2;
    wire c14500;
    assign in14500_1 = {pp127[114]};
    assign in14500_2 = {c13563};
    Full_Adder FA_14500(s14500, c14500, in14500_1, in14500_2, pp126[115]);
    wire[0:0] s14501, in14501_1, in14501_2;
    wire c14501;
    assign in14501_1 = {c13565};
    assign in14501_2 = {c13566};
    Full_Adder FA_14501(s14501, c14501, in14501_1, in14501_2, c13564);
    wire[0:0] s14502, in14502_1, in14502_2;
    wire c14502;
    assign in14502_1 = {s13568[0]};
    assign in14502_2 = {s13569[0]};
    Full_Adder FA_14502(s14502, c14502, in14502_1, in14502_2, s13567[0]);
    wire[0:0] s14503, in14503_1, in14503_2;
    wire c14503;
    assign in14503_1 = {pp122[120]};
    assign in14503_2 = {pp123[119]};
    Full_Adder FA_14503(s14503, c14503, in14503_1, in14503_2, pp121[121]);
    wire[0:0] s14504, in14504_1, in14504_2;
    wire c14504;
    assign in14504_1 = {pp125[117]};
    assign in14504_2 = {pp126[116]};
    Full_Adder FA_14504(s14504, c14504, in14504_1, in14504_2, pp124[118]);
    wire[0:0] s14505, in14505_1, in14505_2;
    wire c14505;
    assign in14505_1 = {c13567};
    assign in14505_2 = {c13568};
    Full_Adder FA_14505(s14505, c14505, in14505_1, in14505_2, pp127[115]);
    wire[0:0] s14506, in14506_1, in14506_2;
    wire c14506;
    assign in14506_1 = {s13570[0]};
    assign in14506_2 = {s13571[0]};
    Full_Adder FA_14506(s14506, c14506, in14506_1, in14506_2, c13569);
    wire[0:0] s14507, in14507_1, in14507_2;
    wire c14507;
    assign in14507_1 = {pp120[123]};
    assign in14507_2 = {pp121[122]};
    Full_Adder FA_14507(s14507, c14507, in14507_1, in14507_2, pp119[124]);
    wire[0:0] s14508, in14508_1, in14508_2;
    wire c14508;
    assign in14508_1 = {pp123[120]};
    assign in14508_2 = {pp124[119]};
    Full_Adder FA_14508(s14508, c14508, in14508_1, in14508_2, pp122[121]);
    wire[0:0] s14509, in14509_1, in14509_2;
    wire c14509;
    assign in14509_1 = {pp126[117]};
    assign in14509_2 = {pp127[116]};
    Full_Adder FA_14509(s14509, c14509, in14509_1, in14509_2, pp125[118]);
    wire[0:0] s14510, in14510_1, in14510_2;
    wire c14510;
    assign in14510_1 = {c13571};
    assign in14510_2 = {s13572[0]};
    Full_Adder FA_14510(s14510, c14510, in14510_1, in14510_2, c13570);
    wire[0:0] s14511, in14511_1, in14511_2;
    wire c14511;
    assign in14511_1 = {pp118[126]};
    assign in14511_2 = {pp119[125]};
    Full_Adder FA_14511(s14511, c14511, in14511_1, in14511_2, pp117[127]);
    wire[0:0] s14512, in14512_1, in14512_2;
    wire c14512;
    assign in14512_1 = {pp121[123]};
    assign in14512_2 = {pp122[122]};
    Full_Adder FA_14512(s14512, c14512, in14512_1, in14512_2, pp120[124]);
    wire[0:0] s14513, in14513_1, in14513_2;
    wire c14513;
    assign in14513_1 = {pp124[120]};
    assign in14513_2 = {pp125[119]};
    Full_Adder FA_14513(s14513, c14513, in14513_1, in14513_2, pp123[121]);
    wire[0:0] s14514, in14514_1, in14514_2;
    wire c14514;
    assign in14514_1 = {pp127[117]};
    assign in14514_2 = {c13572};
    Full_Adder FA_14514(s14514, c14514, in14514_1, in14514_2, pp126[118]);
    wire[0:0] s14515, in14515_1, in14515_2;
    wire c14515;
    assign in14515_1 = {pp119[126]};
    assign in14515_2 = {pp120[125]};
    Full_Adder FA_14515(s14515, c14515, in14515_1, in14515_2, pp118[127]);
    wire[0:0] s14516, in14516_1, in14516_2;
    wire c14516;
    assign in14516_1 = {pp122[123]};
    assign in14516_2 = {pp123[122]};
    Full_Adder FA_14516(s14516, c14516, in14516_1, in14516_2, pp121[124]);
    wire[0:0] s14517, in14517_1, in14517_2;
    wire c14517;
    assign in14517_1 = {pp125[120]};
    assign in14517_2 = {pp126[119]};
    Full_Adder FA_14517(s14517, c14517, in14517_1, in14517_2, pp124[121]);
    wire[0:0] s14518, in14518_1, in14518_2;
    wire c14518;
    assign in14518_1 = {pp120[126]};
    assign in14518_2 = {pp121[125]};
    Full_Adder FA_14518(s14518, c14518, in14518_1, in14518_2, pp119[127]);
    wire[0:0] s14519, in14519_1, in14519_2;
    wire c14519;
    assign in14519_1 = {pp123[123]};
    assign in14519_2 = {pp124[122]};
    Full_Adder FA_14519(s14519, c14519, in14519_1, in14519_2, pp122[124]);
    wire[0:0] s14520, in14520_1, in14520_2;
    wire c14520;
    assign in14520_1 = {pp121[126]};
    assign in14520_2 = {pp122[125]};
    Full_Adder FA_14520(s14520, c14520, in14520_1, in14520_2, pp120[127]);

    /*Stage 8*/
    wire[0:0] s14521, in14521_1, in14521_2;
    wire c14521;
    assign in14521_1 = {pp0[6]};
    assign in14521_2 = {pp1[5]};
    Half_Adder HA_14521(s14521, c14521, in14521_1, in14521_2);
    wire[0:0] s14522, in14522_1, in14522_2;
    wire c14522;
    assign in14522_1 = {pp1[6]};
    assign in14522_2 = {pp2[5]};
    Full_Adder FA_14522(s14522, c14522, in14522_1, in14522_2, pp0[7]);
    wire[0:0] s14523, in14523_1, in14523_2;
    wire c14523;
    assign in14523_1 = {pp3[4]};
    assign in14523_2 = {pp4[3]};
    Half_Adder HA_14523(s14523, c14523, in14523_1, in14523_2);
    wire[0:0] s14524, in14524_1, in14524_2;
    wire c14524;
    assign in14524_1 = {pp3[5]};
    assign in14524_2 = {pp4[4]};
    Full_Adder FA_14524(s14524, c14524, in14524_1, in14524_2, pp2[6]);
    wire[0:0] s14525, in14525_1, in14525_2;
    wire c14525;
    assign in14525_1 = {pp6[2]};
    assign in14525_2 = {pp7[1]};
    Full_Adder FA_14525(s14525, c14525, in14525_1, in14525_2, pp5[3]);
    wire[0:0] s14526, in14526_1, in14526_2;
    wire c14526;
    assign in14526_1 = {pp6[3]};
    assign in14526_2 = {pp7[2]};
    Full_Adder FA_14526(s14526, c14526, in14526_1, in14526_2, pp5[4]);
    wire[0:0] s14527, in14527_1, in14527_2;
    wire c14527;
    assign in14527_1 = {pp9[0]};
    assign in14527_2 = {c13573};
    Full_Adder FA_14527(s14527, c14527, in14527_1, in14527_2, pp8[1]);
    wire[0:0] s14528, in14528_1, in14528_2;
    wire c14528;
    assign in14528_1 = {pp9[1]};
    assign in14528_2 = {pp10[0]};
    Full_Adder FA_14528(s14528, c14528, in14528_1, in14528_2, pp8[2]);
    wire[0:0] s14529, in14529_1, in14529_2;
    wire c14529;
    assign in14529_1 = {c13575};
    assign in14529_2 = {s13576[0]};
    Full_Adder FA_14529(s14529, c14529, in14529_1, in14529_2, c13574);
    wire[0:0] s14530, in14530_1, in14530_2;
    wire c14530;
    assign in14530_1 = {c13576};
    assign in14530_2 = {c13577};
    Full_Adder FA_14530(s14530, c14530, in14530_1, in14530_2, pp11[0]);
    wire[0:0] s14531, in14531_1, in14531_2;
    wire c14531;
    assign in14531_1 = {s13579[0]};
    assign in14531_2 = {s13580[0]};
    Full_Adder FA_14531(s14531, c14531, in14531_1, in14531_2, c13578);
    wire[0:0] s14532, in14532_1, in14532_2;
    wire c14532;
    assign in14532_1 = {c13580};
    assign in14532_2 = {c13581};
    Full_Adder FA_14532(s14532, c14532, in14532_1, in14532_2, c13579);
    wire[0:0] s14533, in14533_1, in14533_2;
    wire c14533;
    assign in14533_1 = {s13583[0]};
    assign in14533_2 = {s13584[0]};
    Full_Adder FA_14533(s14533, c14533, in14533_1, in14533_2, c13582);
    wire[0:0] s14534, in14534_1, in14534_2;
    wire c14534;
    assign in14534_1 = {c13584};
    assign in14534_2 = {c13585};
    Full_Adder FA_14534(s14534, c14534, in14534_1, in14534_2, c13583);
    wire[0:0] s14535, in14535_1, in14535_2;
    wire c14535;
    assign in14535_1 = {s13587[0]};
    assign in14535_2 = {s13588[0]};
    Full_Adder FA_14535(s14535, c14535, in14535_1, in14535_2, c13586);
    wire[0:0] s14536, in14536_1, in14536_2;
    wire c14536;
    assign in14536_1 = {c13588};
    assign in14536_2 = {c13589};
    Full_Adder FA_14536(s14536, c14536, in14536_1, in14536_2, c13587);
    wire[0:0] s14537, in14537_1, in14537_2;
    wire c14537;
    assign in14537_1 = {s13591[0]};
    assign in14537_2 = {s13592[0]};
    Full_Adder FA_14537(s14537, c14537, in14537_1, in14537_2, c13590);
    wire[0:0] s14538, in14538_1, in14538_2;
    wire c14538;
    assign in14538_1 = {c13592};
    assign in14538_2 = {c13593};
    Full_Adder FA_14538(s14538, c14538, in14538_1, in14538_2, c13591);
    wire[0:0] s14539, in14539_1, in14539_2;
    wire c14539;
    assign in14539_1 = {s13595[0]};
    assign in14539_2 = {s13596[0]};
    Full_Adder FA_14539(s14539, c14539, in14539_1, in14539_2, c13594);
    wire[0:0] s14540, in14540_1, in14540_2;
    wire c14540;
    assign in14540_1 = {c13596};
    assign in14540_2 = {c13597};
    Full_Adder FA_14540(s14540, c14540, in14540_1, in14540_2, c13595);
    wire[0:0] s14541, in14541_1, in14541_2;
    wire c14541;
    assign in14541_1 = {s13599[0]};
    assign in14541_2 = {s13600[0]};
    Full_Adder FA_14541(s14541, c14541, in14541_1, in14541_2, c13598);
    wire[0:0] s14542, in14542_1, in14542_2;
    wire c14542;
    assign in14542_1 = {c13600};
    assign in14542_2 = {c13601};
    Full_Adder FA_14542(s14542, c14542, in14542_1, in14542_2, c13599);
    wire[0:0] s14543, in14543_1, in14543_2;
    wire c14543;
    assign in14543_1 = {s13603[0]};
    assign in14543_2 = {s13604[0]};
    Full_Adder FA_14543(s14543, c14543, in14543_1, in14543_2, c13602);
    wire[0:0] s14544, in14544_1, in14544_2;
    wire c14544;
    assign in14544_1 = {c13604};
    assign in14544_2 = {c13605};
    Full_Adder FA_14544(s14544, c14544, in14544_1, in14544_2, c13603);
    wire[0:0] s14545, in14545_1, in14545_2;
    wire c14545;
    assign in14545_1 = {s13607[0]};
    assign in14545_2 = {s13608[0]};
    Full_Adder FA_14545(s14545, c14545, in14545_1, in14545_2, c13606);
    wire[0:0] s14546, in14546_1, in14546_2;
    wire c14546;
    assign in14546_1 = {c13608};
    assign in14546_2 = {c13609};
    Full_Adder FA_14546(s14546, c14546, in14546_1, in14546_2, c13607);
    wire[0:0] s14547, in14547_1, in14547_2;
    wire c14547;
    assign in14547_1 = {s13611[0]};
    assign in14547_2 = {s13612[0]};
    Full_Adder FA_14547(s14547, c14547, in14547_1, in14547_2, c13610);
    wire[0:0] s14548, in14548_1, in14548_2;
    wire c14548;
    assign in14548_1 = {c13612};
    assign in14548_2 = {c13613};
    Full_Adder FA_14548(s14548, c14548, in14548_1, in14548_2, c13611);
    wire[0:0] s14549, in14549_1, in14549_2;
    wire c14549;
    assign in14549_1 = {s13615[0]};
    assign in14549_2 = {s13616[0]};
    Full_Adder FA_14549(s14549, c14549, in14549_1, in14549_2, c13614);
    wire[0:0] s14550, in14550_1, in14550_2;
    wire c14550;
    assign in14550_1 = {c13616};
    assign in14550_2 = {c13617};
    Full_Adder FA_14550(s14550, c14550, in14550_1, in14550_2, c13615);
    wire[0:0] s14551, in14551_1, in14551_2;
    wire c14551;
    assign in14551_1 = {s13619[0]};
    assign in14551_2 = {s13620[0]};
    Full_Adder FA_14551(s14551, c14551, in14551_1, in14551_2, c13618);
    wire[0:0] s14552, in14552_1, in14552_2;
    wire c14552;
    assign in14552_1 = {c13620};
    assign in14552_2 = {c13621};
    Full_Adder FA_14552(s14552, c14552, in14552_1, in14552_2, c13619);
    wire[0:0] s14553, in14553_1, in14553_2;
    wire c14553;
    assign in14553_1 = {s13623[0]};
    assign in14553_2 = {s13624[0]};
    Full_Adder FA_14553(s14553, c14553, in14553_1, in14553_2, c13622);
    wire[0:0] s14554, in14554_1, in14554_2;
    wire c14554;
    assign in14554_1 = {c13624};
    assign in14554_2 = {c13625};
    Full_Adder FA_14554(s14554, c14554, in14554_1, in14554_2, c13623);
    wire[0:0] s14555, in14555_1, in14555_2;
    wire c14555;
    assign in14555_1 = {s13627[0]};
    assign in14555_2 = {s13628[0]};
    Full_Adder FA_14555(s14555, c14555, in14555_1, in14555_2, c13626);
    wire[0:0] s14556, in14556_1, in14556_2;
    wire c14556;
    assign in14556_1 = {c13628};
    assign in14556_2 = {c13629};
    Full_Adder FA_14556(s14556, c14556, in14556_1, in14556_2, c13627);
    wire[0:0] s14557, in14557_1, in14557_2;
    wire c14557;
    assign in14557_1 = {s13631[0]};
    assign in14557_2 = {s13632[0]};
    Full_Adder FA_14557(s14557, c14557, in14557_1, in14557_2, c13630);
    wire[0:0] s14558, in14558_1, in14558_2;
    wire c14558;
    assign in14558_1 = {c13632};
    assign in14558_2 = {c13633};
    Full_Adder FA_14558(s14558, c14558, in14558_1, in14558_2, c13631);
    wire[0:0] s14559, in14559_1, in14559_2;
    wire c14559;
    assign in14559_1 = {s13635[0]};
    assign in14559_2 = {s13636[0]};
    Full_Adder FA_14559(s14559, c14559, in14559_1, in14559_2, c13634);
    wire[0:0] s14560, in14560_1, in14560_2;
    wire c14560;
    assign in14560_1 = {c13636};
    assign in14560_2 = {c13637};
    Full_Adder FA_14560(s14560, c14560, in14560_1, in14560_2, c13635);
    wire[0:0] s14561, in14561_1, in14561_2;
    wire c14561;
    assign in14561_1 = {s13639[0]};
    assign in14561_2 = {s13640[0]};
    Full_Adder FA_14561(s14561, c14561, in14561_1, in14561_2, c13638);
    wire[0:0] s14562, in14562_1, in14562_2;
    wire c14562;
    assign in14562_1 = {c13640};
    assign in14562_2 = {c13641};
    Full_Adder FA_14562(s14562, c14562, in14562_1, in14562_2, c13639);
    wire[0:0] s14563, in14563_1, in14563_2;
    wire c14563;
    assign in14563_1 = {s13643[0]};
    assign in14563_2 = {s13644[0]};
    Full_Adder FA_14563(s14563, c14563, in14563_1, in14563_2, c13642);
    wire[0:0] s14564, in14564_1, in14564_2;
    wire c14564;
    assign in14564_1 = {c13644};
    assign in14564_2 = {c13645};
    Full_Adder FA_14564(s14564, c14564, in14564_1, in14564_2, c13643);
    wire[0:0] s14565, in14565_1, in14565_2;
    wire c14565;
    assign in14565_1 = {s13647[0]};
    assign in14565_2 = {s13648[0]};
    Full_Adder FA_14565(s14565, c14565, in14565_1, in14565_2, c13646);
    wire[0:0] s14566, in14566_1, in14566_2;
    wire c14566;
    assign in14566_1 = {c13648};
    assign in14566_2 = {c13649};
    Full_Adder FA_14566(s14566, c14566, in14566_1, in14566_2, c13647);
    wire[0:0] s14567, in14567_1, in14567_2;
    wire c14567;
    assign in14567_1 = {s13651[0]};
    assign in14567_2 = {s13652[0]};
    Full_Adder FA_14567(s14567, c14567, in14567_1, in14567_2, c13650);
    wire[0:0] s14568, in14568_1, in14568_2;
    wire c14568;
    assign in14568_1 = {c13652};
    assign in14568_2 = {c13653};
    Full_Adder FA_14568(s14568, c14568, in14568_1, in14568_2, c13651);
    wire[0:0] s14569, in14569_1, in14569_2;
    wire c14569;
    assign in14569_1 = {s13655[0]};
    assign in14569_2 = {s13656[0]};
    Full_Adder FA_14569(s14569, c14569, in14569_1, in14569_2, c13654);
    wire[0:0] s14570, in14570_1, in14570_2;
    wire c14570;
    assign in14570_1 = {c13656};
    assign in14570_2 = {c13657};
    Full_Adder FA_14570(s14570, c14570, in14570_1, in14570_2, c13655);
    wire[0:0] s14571, in14571_1, in14571_2;
    wire c14571;
    assign in14571_1 = {s13659[0]};
    assign in14571_2 = {s13660[0]};
    Full_Adder FA_14571(s14571, c14571, in14571_1, in14571_2, c13658);
    wire[0:0] s14572, in14572_1, in14572_2;
    wire c14572;
    assign in14572_1 = {c13660};
    assign in14572_2 = {c13661};
    Full_Adder FA_14572(s14572, c14572, in14572_1, in14572_2, c13659);
    wire[0:0] s14573, in14573_1, in14573_2;
    wire c14573;
    assign in14573_1 = {s13663[0]};
    assign in14573_2 = {s13664[0]};
    Full_Adder FA_14573(s14573, c14573, in14573_1, in14573_2, c13662);
    wire[0:0] s14574, in14574_1, in14574_2;
    wire c14574;
    assign in14574_1 = {c13664};
    assign in14574_2 = {c13665};
    Full_Adder FA_14574(s14574, c14574, in14574_1, in14574_2, c13663);
    wire[0:0] s14575, in14575_1, in14575_2;
    wire c14575;
    assign in14575_1 = {s13667[0]};
    assign in14575_2 = {s13668[0]};
    Full_Adder FA_14575(s14575, c14575, in14575_1, in14575_2, c13666);
    wire[0:0] s14576, in14576_1, in14576_2;
    wire c14576;
    assign in14576_1 = {c13668};
    assign in14576_2 = {c13669};
    Full_Adder FA_14576(s14576, c14576, in14576_1, in14576_2, c13667);
    wire[0:0] s14577, in14577_1, in14577_2;
    wire c14577;
    assign in14577_1 = {s13671[0]};
    assign in14577_2 = {s13672[0]};
    Full_Adder FA_14577(s14577, c14577, in14577_1, in14577_2, c13670);
    wire[0:0] s14578, in14578_1, in14578_2;
    wire c14578;
    assign in14578_1 = {c13672};
    assign in14578_2 = {c13673};
    Full_Adder FA_14578(s14578, c14578, in14578_1, in14578_2, c13671);
    wire[0:0] s14579, in14579_1, in14579_2;
    wire c14579;
    assign in14579_1 = {s13675[0]};
    assign in14579_2 = {s13676[0]};
    Full_Adder FA_14579(s14579, c14579, in14579_1, in14579_2, c13674);
    wire[0:0] s14580, in14580_1, in14580_2;
    wire c14580;
    assign in14580_1 = {c13676};
    assign in14580_2 = {c13677};
    Full_Adder FA_14580(s14580, c14580, in14580_1, in14580_2, c13675);
    wire[0:0] s14581, in14581_1, in14581_2;
    wire c14581;
    assign in14581_1 = {s13679[0]};
    assign in14581_2 = {s13680[0]};
    Full_Adder FA_14581(s14581, c14581, in14581_1, in14581_2, c13678);
    wire[0:0] s14582, in14582_1, in14582_2;
    wire c14582;
    assign in14582_1 = {c13680};
    assign in14582_2 = {c13681};
    Full_Adder FA_14582(s14582, c14582, in14582_1, in14582_2, c13679);
    wire[0:0] s14583, in14583_1, in14583_2;
    wire c14583;
    assign in14583_1 = {s13683[0]};
    assign in14583_2 = {s13684[0]};
    Full_Adder FA_14583(s14583, c14583, in14583_1, in14583_2, c13682);
    wire[0:0] s14584, in14584_1, in14584_2;
    wire c14584;
    assign in14584_1 = {c13684};
    assign in14584_2 = {c13685};
    Full_Adder FA_14584(s14584, c14584, in14584_1, in14584_2, c13683);
    wire[0:0] s14585, in14585_1, in14585_2;
    wire c14585;
    assign in14585_1 = {s13687[0]};
    assign in14585_2 = {s13688[0]};
    Full_Adder FA_14585(s14585, c14585, in14585_1, in14585_2, c13686);
    wire[0:0] s14586, in14586_1, in14586_2;
    wire c14586;
    assign in14586_1 = {c13688};
    assign in14586_2 = {c13689};
    Full_Adder FA_14586(s14586, c14586, in14586_1, in14586_2, c13687);
    wire[0:0] s14587, in14587_1, in14587_2;
    wire c14587;
    assign in14587_1 = {s13691[0]};
    assign in14587_2 = {s13692[0]};
    Full_Adder FA_14587(s14587, c14587, in14587_1, in14587_2, c13690);
    wire[0:0] s14588, in14588_1, in14588_2;
    wire c14588;
    assign in14588_1 = {c13692};
    assign in14588_2 = {c13693};
    Full_Adder FA_14588(s14588, c14588, in14588_1, in14588_2, c13691);
    wire[0:0] s14589, in14589_1, in14589_2;
    wire c14589;
    assign in14589_1 = {s13695[0]};
    assign in14589_2 = {s13696[0]};
    Full_Adder FA_14589(s14589, c14589, in14589_1, in14589_2, c13694);
    wire[0:0] s14590, in14590_1, in14590_2;
    wire c14590;
    assign in14590_1 = {c13696};
    assign in14590_2 = {c13697};
    Full_Adder FA_14590(s14590, c14590, in14590_1, in14590_2, c13695);
    wire[0:0] s14591, in14591_1, in14591_2;
    wire c14591;
    assign in14591_1 = {s13699[0]};
    assign in14591_2 = {s13700[0]};
    Full_Adder FA_14591(s14591, c14591, in14591_1, in14591_2, c13698);
    wire[0:0] s14592, in14592_1, in14592_2;
    wire c14592;
    assign in14592_1 = {c13700};
    assign in14592_2 = {c13701};
    Full_Adder FA_14592(s14592, c14592, in14592_1, in14592_2, c13699);
    wire[0:0] s14593, in14593_1, in14593_2;
    wire c14593;
    assign in14593_1 = {s13703[0]};
    assign in14593_2 = {s13704[0]};
    Full_Adder FA_14593(s14593, c14593, in14593_1, in14593_2, c13702);
    wire[0:0] s14594, in14594_1, in14594_2;
    wire c14594;
    assign in14594_1 = {c13704};
    assign in14594_2 = {c13705};
    Full_Adder FA_14594(s14594, c14594, in14594_1, in14594_2, c13703);
    wire[0:0] s14595, in14595_1, in14595_2;
    wire c14595;
    assign in14595_1 = {s13707[0]};
    assign in14595_2 = {s13708[0]};
    Full_Adder FA_14595(s14595, c14595, in14595_1, in14595_2, c13706);
    wire[0:0] s14596, in14596_1, in14596_2;
    wire c14596;
    assign in14596_1 = {c13708};
    assign in14596_2 = {c13709};
    Full_Adder FA_14596(s14596, c14596, in14596_1, in14596_2, c13707);
    wire[0:0] s14597, in14597_1, in14597_2;
    wire c14597;
    assign in14597_1 = {s13711[0]};
    assign in14597_2 = {s13712[0]};
    Full_Adder FA_14597(s14597, c14597, in14597_1, in14597_2, c13710);
    wire[0:0] s14598, in14598_1, in14598_2;
    wire c14598;
    assign in14598_1 = {c13712};
    assign in14598_2 = {c13713};
    Full_Adder FA_14598(s14598, c14598, in14598_1, in14598_2, c13711);
    wire[0:0] s14599, in14599_1, in14599_2;
    wire c14599;
    assign in14599_1 = {s13715[0]};
    assign in14599_2 = {s13716[0]};
    Full_Adder FA_14599(s14599, c14599, in14599_1, in14599_2, c13714);
    wire[0:0] s14600, in14600_1, in14600_2;
    wire c14600;
    assign in14600_1 = {c13716};
    assign in14600_2 = {c13717};
    Full_Adder FA_14600(s14600, c14600, in14600_1, in14600_2, c13715);
    wire[0:0] s14601, in14601_1, in14601_2;
    wire c14601;
    assign in14601_1 = {s13719[0]};
    assign in14601_2 = {s13720[0]};
    Full_Adder FA_14601(s14601, c14601, in14601_1, in14601_2, c13718);
    wire[0:0] s14602, in14602_1, in14602_2;
    wire c14602;
    assign in14602_1 = {c13720};
    assign in14602_2 = {c13721};
    Full_Adder FA_14602(s14602, c14602, in14602_1, in14602_2, c13719);
    wire[0:0] s14603, in14603_1, in14603_2;
    wire c14603;
    assign in14603_1 = {s13723[0]};
    assign in14603_2 = {s13724[0]};
    Full_Adder FA_14603(s14603, c14603, in14603_1, in14603_2, c13722);
    wire[0:0] s14604, in14604_1, in14604_2;
    wire c14604;
    assign in14604_1 = {c13724};
    assign in14604_2 = {c13725};
    Full_Adder FA_14604(s14604, c14604, in14604_1, in14604_2, c13723);
    wire[0:0] s14605, in14605_1, in14605_2;
    wire c14605;
    assign in14605_1 = {s13727[0]};
    assign in14605_2 = {s13728[0]};
    Full_Adder FA_14605(s14605, c14605, in14605_1, in14605_2, c13726);
    wire[0:0] s14606, in14606_1, in14606_2;
    wire c14606;
    assign in14606_1 = {c13728};
    assign in14606_2 = {c13729};
    Full_Adder FA_14606(s14606, c14606, in14606_1, in14606_2, c13727);
    wire[0:0] s14607, in14607_1, in14607_2;
    wire c14607;
    assign in14607_1 = {s13731[0]};
    assign in14607_2 = {s13732[0]};
    Full_Adder FA_14607(s14607, c14607, in14607_1, in14607_2, c13730);
    wire[0:0] s14608, in14608_1, in14608_2;
    wire c14608;
    assign in14608_1 = {c13732};
    assign in14608_2 = {c13733};
    Full_Adder FA_14608(s14608, c14608, in14608_1, in14608_2, c13731);
    wire[0:0] s14609, in14609_1, in14609_2;
    wire c14609;
    assign in14609_1 = {s13735[0]};
    assign in14609_2 = {s13736[0]};
    Full_Adder FA_14609(s14609, c14609, in14609_1, in14609_2, c13734);
    wire[0:0] s14610, in14610_1, in14610_2;
    wire c14610;
    assign in14610_1 = {c13736};
    assign in14610_2 = {c13737};
    Full_Adder FA_14610(s14610, c14610, in14610_1, in14610_2, c13735);
    wire[0:0] s14611, in14611_1, in14611_2;
    wire c14611;
    assign in14611_1 = {s13739[0]};
    assign in14611_2 = {s13740[0]};
    Full_Adder FA_14611(s14611, c14611, in14611_1, in14611_2, c13738);
    wire[0:0] s14612, in14612_1, in14612_2;
    wire c14612;
    assign in14612_1 = {c13740};
    assign in14612_2 = {c13741};
    Full_Adder FA_14612(s14612, c14612, in14612_1, in14612_2, c13739);
    wire[0:0] s14613, in14613_1, in14613_2;
    wire c14613;
    assign in14613_1 = {s13743[0]};
    assign in14613_2 = {s13744[0]};
    Full_Adder FA_14613(s14613, c14613, in14613_1, in14613_2, c13742);
    wire[0:0] s14614, in14614_1, in14614_2;
    wire c14614;
    assign in14614_1 = {c13744};
    assign in14614_2 = {c13745};
    Full_Adder FA_14614(s14614, c14614, in14614_1, in14614_2, c13743);
    wire[0:0] s14615, in14615_1, in14615_2;
    wire c14615;
    assign in14615_1 = {s13747[0]};
    assign in14615_2 = {s13748[0]};
    Full_Adder FA_14615(s14615, c14615, in14615_1, in14615_2, c13746);
    wire[0:0] s14616, in14616_1, in14616_2;
    wire c14616;
    assign in14616_1 = {c13748};
    assign in14616_2 = {c13749};
    Full_Adder FA_14616(s14616, c14616, in14616_1, in14616_2, c13747);
    wire[0:0] s14617, in14617_1, in14617_2;
    wire c14617;
    assign in14617_1 = {s13751[0]};
    assign in14617_2 = {s13752[0]};
    Full_Adder FA_14617(s14617, c14617, in14617_1, in14617_2, c13750);
    wire[0:0] s14618, in14618_1, in14618_2;
    wire c14618;
    assign in14618_1 = {c13752};
    assign in14618_2 = {c13753};
    Full_Adder FA_14618(s14618, c14618, in14618_1, in14618_2, c13751);
    wire[0:0] s14619, in14619_1, in14619_2;
    wire c14619;
    assign in14619_1 = {s13755[0]};
    assign in14619_2 = {s13756[0]};
    Full_Adder FA_14619(s14619, c14619, in14619_1, in14619_2, c13754);
    wire[0:0] s14620, in14620_1, in14620_2;
    wire c14620;
    assign in14620_1 = {c13756};
    assign in14620_2 = {c13757};
    Full_Adder FA_14620(s14620, c14620, in14620_1, in14620_2, c13755);
    wire[0:0] s14621, in14621_1, in14621_2;
    wire c14621;
    assign in14621_1 = {s13759[0]};
    assign in14621_2 = {s13760[0]};
    Full_Adder FA_14621(s14621, c14621, in14621_1, in14621_2, c13758);
    wire[0:0] s14622, in14622_1, in14622_2;
    wire c14622;
    assign in14622_1 = {c13760};
    assign in14622_2 = {c13761};
    Full_Adder FA_14622(s14622, c14622, in14622_1, in14622_2, c13759);
    wire[0:0] s14623, in14623_1, in14623_2;
    wire c14623;
    assign in14623_1 = {s13763[0]};
    assign in14623_2 = {s13764[0]};
    Full_Adder FA_14623(s14623, c14623, in14623_1, in14623_2, c13762);
    wire[0:0] s14624, in14624_1, in14624_2;
    wire c14624;
    assign in14624_1 = {c13764};
    assign in14624_2 = {c13765};
    Full_Adder FA_14624(s14624, c14624, in14624_1, in14624_2, c13763);
    wire[0:0] s14625, in14625_1, in14625_2;
    wire c14625;
    assign in14625_1 = {s13767[0]};
    assign in14625_2 = {s13768[0]};
    Full_Adder FA_14625(s14625, c14625, in14625_1, in14625_2, c13766);
    wire[0:0] s14626, in14626_1, in14626_2;
    wire c14626;
    assign in14626_1 = {c13768};
    assign in14626_2 = {c13769};
    Full_Adder FA_14626(s14626, c14626, in14626_1, in14626_2, c13767);
    wire[0:0] s14627, in14627_1, in14627_2;
    wire c14627;
    assign in14627_1 = {s13771[0]};
    assign in14627_2 = {s13772[0]};
    Full_Adder FA_14627(s14627, c14627, in14627_1, in14627_2, c13770);
    wire[0:0] s14628, in14628_1, in14628_2;
    wire c14628;
    assign in14628_1 = {c13772};
    assign in14628_2 = {c13773};
    Full_Adder FA_14628(s14628, c14628, in14628_1, in14628_2, c13771);
    wire[0:0] s14629, in14629_1, in14629_2;
    wire c14629;
    assign in14629_1 = {s13775[0]};
    assign in14629_2 = {s13776[0]};
    Full_Adder FA_14629(s14629, c14629, in14629_1, in14629_2, c13774);
    wire[0:0] s14630, in14630_1, in14630_2;
    wire c14630;
    assign in14630_1 = {c13776};
    assign in14630_2 = {c13777};
    Full_Adder FA_14630(s14630, c14630, in14630_1, in14630_2, c13775);
    wire[0:0] s14631, in14631_1, in14631_2;
    wire c14631;
    assign in14631_1 = {s13779[0]};
    assign in14631_2 = {s13780[0]};
    Full_Adder FA_14631(s14631, c14631, in14631_1, in14631_2, c13778);
    wire[0:0] s14632, in14632_1, in14632_2;
    wire c14632;
    assign in14632_1 = {c13780};
    assign in14632_2 = {c13781};
    Full_Adder FA_14632(s14632, c14632, in14632_1, in14632_2, c13779);
    wire[0:0] s14633, in14633_1, in14633_2;
    wire c14633;
    assign in14633_1 = {s13783[0]};
    assign in14633_2 = {s13784[0]};
    Full_Adder FA_14633(s14633, c14633, in14633_1, in14633_2, c13782);
    wire[0:0] s14634, in14634_1, in14634_2;
    wire c14634;
    assign in14634_1 = {c13784};
    assign in14634_2 = {c13785};
    Full_Adder FA_14634(s14634, c14634, in14634_1, in14634_2, c13783);
    wire[0:0] s14635, in14635_1, in14635_2;
    wire c14635;
    assign in14635_1 = {s13787[0]};
    assign in14635_2 = {s13788[0]};
    Full_Adder FA_14635(s14635, c14635, in14635_1, in14635_2, c13786);
    wire[0:0] s14636, in14636_1, in14636_2;
    wire c14636;
    assign in14636_1 = {c13788};
    assign in14636_2 = {c13789};
    Full_Adder FA_14636(s14636, c14636, in14636_1, in14636_2, c13787);
    wire[0:0] s14637, in14637_1, in14637_2;
    wire c14637;
    assign in14637_1 = {s13791[0]};
    assign in14637_2 = {s13792[0]};
    Full_Adder FA_14637(s14637, c14637, in14637_1, in14637_2, c13790);
    wire[0:0] s14638, in14638_1, in14638_2;
    wire c14638;
    assign in14638_1 = {c13792};
    assign in14638_2 = {c13793};
    Full_Adder FA_14638(s14638, c14638, in14638_1, in14638_2, c13791);
    wire[0:0] s14639, in14639_1, in14639_2;
    wire c14639;
    assign in14639_1 = {s13795[0]};
    assign in14639_2 = {s13796[0]};
    Full_Adder FA_14639(s14639, c14639, in14639_1, in14639_2, c13794);
    wire[0:0] s14640, in14640_1, in14640_2;
    wire c14640;
    assign in14640_1 = {c13796};
    assign in14640_2 = {c13797};
    Full_Adder FA_14640(s14640, c14640, in14640_1, in14640_2, c13795);
    wire[0:0] s14641, in14641_1, in14641_2;
    wire c14641;
    assign in14641_1 = {s13799[0]};
    assign in14641_2 = {s13800[0]};
    Full_Adder FA_14641(s14641, c14641, in14641_1, in14641_2, c13798);
    wire[0:0] s14642, in14642_1, in14642_2;
    wire c14642;
    assign in14642_1 = {c13800};
    assign in14642_2 = {c13801};
    Full_Adder FA_14642(s14642, c14642, in14642_1, in14642_2, c13799);
    wire[0:0] s14643, in14643_1, in14643_2;
    wire c14643;
    assign in14643_1 = {s13803[0]};
    assign in14643_2 = {s13804[0]};
    Full_Adder FA_14643(s14643, c14643, in14643_1, in14643_2, c13802);
    wire[0:0] s14644, in14644_1, in14644_2;
    wire c14644;
    assign in14644_1 = {c13804};
    assign in14644_2 = {c13805};
    Full_Adder FA_14644(s14644, c14644, in14644_1, in14644_2, c13803);
    wire[0:0] s14645, in14645_1, in14645_2;
    wire c14645;
    assign in14645_1 = {s13807[0]};
    assign in14645_2 = {s13808[0]};
    Full_Adder FA_14645(s14645, c14645, in14645_1, in14645_2, c13806);
    wire[0:0] s14646, in14646_1, in14646_2;
    wire c14646;
    assign in14646_1 = {c13808};
    assign in14646_2 = {c13809};
    Full_Adder FA_14646(s14646, c14646, in14646_1, in14646_2, c13807);
    wire[0:0] s14647, in14647_1, in14647_2;
    wire c14647;
    assign in14647_1 = {s13811[0]};
    assign in14647_2 = {s13812[0]};
    Full_Adder FA_14647(s14647, c14647, in14647_1, in14647_2, c13810);
    wire[0:0] s14648, in14648_1, in14648_2;
    wire c14648;
    assign in14648_1 = {c13812};
    assign in14648_2 = {c13813};
    Full_Adder FA_14648(s14648, c14648, in14648_1, in14648_2, c13811);
    wire[0:0] s14649, in14649_1, in14649_2;
    wire c14649;
    assign in14649_1 = {s13815[0]};
    assign in14649_2 = {s13816[0]};
    Full_Adder FA_14649(s14649, c14649, in14649_1, in14649_2, c13814);
    wire[0:0] s14650, in14650_1, in14650_2;
    wire c14650;
    assign in14650_1 = {c13816};
    assign in14650_2 = {c13817};
    Full_Adder FA_14650(s14650, c14650, in14650_1, in14650_2, c13815);
    wire[0:0] s14651, in14651_1, in14651_2;
    wire c14651;
    assign in14651_1 = {s13819[0]};
    assign in14651_2 = {s13820[0]};
    Full_Adder FA_14651(s14651, c14651, in14651_1, in14651_2, c13818);
    wire[0:0] s14652, in14652_1, in14652_2;
    wire c14652;
    assign in14652_1 = {c13820};
    assign in14652_2 = {c13821};
    Full_Adder FA_14652(s14652, c14652, in14652_1, in14652_2, c13819);
    wire[0:0] s14653, in14653_1, in14653_2;
    wire c14653;
    assign in14653_1 = {s13823[0]};
    assign in14653_2 = {s13824[0]};
    Full_Adder FA_14653(s14653, c14653, in14653_1, in14653_2, c13822);
    wire[0:0] s14654, in14654_1, in14654_2;
    wire c14654;
    assign in14654_1 = {c13824};
    assign in14654_2 = {c13825};
    Full_Adder FA_14654(s14654, c14654, in14654_1, in14654_2, c13823);
    wire[0:0] s14655, in14655_1, in14655_2;
    wire c14655;
    assign in14655_1 = {s13827[0]};
    assign in14655_2 = {s13828[0]};
    Full_Adder FA_14655(s14655, c14655, in14655_1, in14655_2, c13826);
    wire[0:0] s14656, in14656_1, in14656_2;
    wire c14656;
    assign in14656_1 = {c13828};
    assign in14656_2 = {c13829};
    Full_Adder FA_14656(s14656, c14656, in14656_1, in14656_2, c13827);
    wire[0:0] s14657, in14657_1, in14657_2;
    wire c14657;
    assign in14657_1 = {s13831[0]};
    assign in14657_2 = {s13832[0]};
    Full_Adder FA_14657(s14657, c14657, in14657_1, in14657_2, c13830);
    wire[0:0] s14658, in14658_1, in14658_2;
    wire c14658;
    assign in14658_1 = {c13832};
    assign in14658_2 = {c13833};
    Full_Adder FA_14658(s14658, c14658, in14658_1, in14658_2, c13831);
    wire[0:0] s14659, in14659_1, in14659_2;
    wire c14659;
    assign in14659_1 = {s13835[0]};
    assign in14659_2 = {s13836[0]};
    Full_Adder FA_14659(s14659, c14659, in14659_1, in14659_2, c13834);
    wire[0:0] s14660, in14660_1, in14660_2;
    wire c14660;
    assign in14660_1 = {c13836};
    assign in14660_2 = {c13837};
    Full_Adder FA_14660(s14660, c14660, in14660_1, in14660_2, c13835);
    wire[0:0] s14661, in14661_1, in14661_2;
    wire c14661;
    assign in14661_1 = {s13839[0]};
    assign in14661_2 = {s13840[0]};
    Full_Adder FA_14661(s14661, c14661, in14661_1, in14661_2, c13838);
    wire[0:0] s14662, in14662_1, in14662_2;
    wire c14662;
    assign in14662_1 = {c13840};
    assign in14662_2 = {c13841};
    Full_Adder FA_14662(s14662, c14662, in14662_1, in14662_2, c13839);
    wire[0:0] s14663, in14663_1, in14663_2;
    wire c14663;
    assign in14663_1 = {s13843[0]};
    assign in14663_2 = {s13844[0]};
    Full_Adder FA_14663(s14663, c14663, in14663_1, in14663_2, c13842);
    wire[0:0] s14664, in14664_1, in14664_2;
    wire c14664;
    assign in14664_1 = {c13844};
    assign in14664_2 = {c13845};
    Full_Adder FA_14664(s14664, c14664, in14664_1, in14664_2, c13843);
    wire[0:0] s14665, in14665_1, in14665_2;
    wire c14665;
    assign in14665_1 = {s13847[0]};
    assign in14665_2 = {s13848[0]};
    Full_Adder FA_14665(s14665, c14665, in14665_1, in14665_2, c13846);
    wire[0:0] s14666, in14666_1, in14666_2;
    wire c14666;
    assign in14666_1 = {c13848};
    assign in14666_2 = {c13849};
    Full_Adder FA_14666(s14666, c14666, in14666_1, in14666_2, c13847);
    wire[0:0] s14667, in14667_1, in14667_2;
    wire c14667;
    assign in14667_1 = {s13851[0]};
    assign in14667_2 = {s13852[0]};
    Full_Adder FA_14667(s14667, c14667, in14667_1, in14667_2, c13850);
    wire[0:0] s14668, in14668_1, in14668_2;
    wire c14668;
    assign in14668_1 = {c13852};
    assign in14668_2 = {c13853};
    Full_Adder FA_14668(s14668, c14668, in14668_1, in14668_2, c13851);
    wire[0:0] s14669, in14669_1, in14669_2;
    wire c14669;
    assign in14669_1 = {s13855[0]};
    assign in14669_2 = {s13856[0]};
    Full_Adder FA_14669(s14669, c14669, in14669_1, in14669_2, c13854);
    wire[0:0] s14670, in14670_1, in14670_2;
    wire c14670;
    assign in14670_1 = {c13856};
    assign in14670_2 = {c13857};
    Full_Adder FA_14670(s14670, c14670, in14670_1, in14670_2, c13855);
    wire[0:0] s14671, in14671_1, in14671_2;
    wire c14671;
    assign in14671_1 = {s13859[0]};
    assign in14671_2 = {s13860[0]};
    Full_Adder FA_14671(s14671, c14671, in14671_1, in14671_2, c13858);
    wire[0:0] s14672, in14672_1, in14672_2;
    wire c14672;
    assign in14672_1 = {c13860};
    assign in14672_2 = {c13861};
    Full_Adder FA_14672(s14672, c14672, in14672_1, in14672_2, c13859);
    wire[0:0] s14673, in14673_1, in14673_2;
    wire c14673;
    assign in14673_1 = {s13863[0]};
    assign in14673_2 = {s13864[0]};
    Full_Adder FA_14673(s14673, c14673, in14673_1, in14673_2, c13862);
    wire[0:0] s14674, in14674_1, in14674_2;
    wire c14674;
    assign in14674_1 = {c13864};
    assign in14674_2 = {c13865};
    Full_Adder FA_14674(s14674, c14674, in14674_1, in14674_2, c13863);
    wire[0:0] s14675, in14675_1, in14675_2;
    wire c14675;
    assign in14675_1 = {s13867[0]};
    assign in14675_2 = {s13868[0]};
    Full_Adder FA_14675(s14675, c14675, in14675_1, in14675_2, c13866);
    wire[0:0] s14676, in14676_1, in14676_2;
    wire c14676;
    assign in14676_1 = {c13868};
    assign in14676_2 = {c13869};
    Full_Adder FA_14676(s14676, c14676, in14676_1, in14676_2, c13867);
    wire[0:0] s14677, in14677_1, in14677_2;
    wire c14677;
    assign in14677_1 = {s13871[0]};
    assign in14677_2 = {s13872[0]};
    Full_Adder FA_14677(s14677, c14677, in14677_1, in14677_2, c13870);
    wire[0:0] s14678, in14678_1, in14678_2;
    wire c14678;
    assign in14678_1 = {c13872};
    assign in14678_2 = {c13873};
    Full_Adder FA_14678(s14678, c14678, in14678_1, in14678_2, c13871);
    wire[0:0] s14679, in14679_1, in14679_2;
    wire c14679;
    assign in14679_1 = {s13875[0]};
    assign in14679_2 = {s13876[0]};
    Full_Adder FA_14679(s14679, c14679, in14679_1, in14679_2, c13874);
    wire[0:0] s14680, in14680_1, in14680_2;
    wire c14680;
    assign in14680_1 = {c13876};
    assign in14680_2 = {c13877};
    Full_Adder FA_14680(s14680, c14680, in14680_1, in14680_2, c13875);
    wire[0:0] s14681, in14681_1, in14681_2;
    wire c14681;
    assign in14681_1 = {s13879[0]};
    assign in14681_2 = {s13880[0]};
    Full_Adder FA_14681(s14681, c14681, in14681_1, in14681_2, c13878);
    wire[0:0] s14682, in14682_1, in14682_2;
    wire c14682;
    assign in14682_1 = {c13880};
    assign in14682_2 = {c13881};
    Full_Adder FA_14682(s14682, c14682, in14682_1, in14682_2, c13879);
    wire[0:0] s14683, in14683_1, in14683_2;
    wire c14683;
    assign in14683_1 = {s13883[0]};
    assign in14683_2 = {s13884[0]};
    Full_Adder FA_14683(s14683, c14683, in14683_1, in14683_2, c13882);
    wire[0:0] s14684, in14684_1, in14684_2;
    wire c14684;
    assign in14684_1 = {c13884};
    assign in14684_2 = {c13885};
    Full_Adder FA_14684(s14684, c14684, in14684_1, in14684_2, c13883);
    wire[0:0] s14685, in14685_1, in14685_2;
    wire c14685;
    assign in14685_1 = {s13887[0]};
    assign in14685_2 = {s13888[0]};
    Full_Adder FA_14685(s14685, c14685, in14685_1, in14685_2, c13886);
    wire[0:0] s14686, in14686_1, in14686_2;
    wire c14686;
    assign in14686_1 = {c13888};
    assign in14686_2 = {c13889};
    Full_Adder FA_14686(s14686, c14686, in14686_1, in14686_2, c13887);
    wire[0:0] s14687, in14687_1, in14687_2;
    wire c14687;
    assign in14687_1 = {s13891[0]};
    assign in14687_2 = {s13892[0]};
    Full_Adder FA_14687(s14687, c14687, in14687_1, in14687_2, c13890);
    wire[0:0] s14688, in14688_1, in14688_2;
    wire c14688;
    assign in14688_1 = {c13892};
    assign in14688_2 = {c13893};
    Full_Adder FA_14688(s14688, c14688, in14688_1, in14688_2, c13891);
    wire[0:0] s14689, in14689_1, in14689_2;
    wire c14689;
    assign in14689_1 = {s13895[0]};
    assign in14689_2 = {s13896[0]};
    Full_Adder FA_14689(s14689, c14689, in14689_1, in14689_2, c13894);
    wire[0:0] s14690, in14690_1, in14690_2;
    wire c14690;
    assign in14690_1 = {c13896};
    assign in14690_2 = {c13897};
    Full_Adder FA_14690(s14690, c14690, in14690_1, in14690_2, c13895);
    wire[0:0] s14691, in14691_1, in14691_2;
    wire c14691;
    assign in14691_1 = {s13899[0]};
    assign in14691_2 = {s13900[0]};
    Full_Adder FA_14691(s14691, c14691, in14691_1, in14691_2, c13898);
    wire[0:0] s14692, in14692_1, in14692_2;
    wire c14692;
    assign in14692_1 = {c13900};
    assign in14692_2 = {c13901};
    Full_Adder FA_14692(s14692, c14692, in14692_1, in14692_2, c13899);
    wire[0:0] s14693, in14693_1, in14693_2;
    wire c14693;
    assign in14693_1 = {s13903[0]};
    assign in14693_2 = {s13904[0]};
    Full_Adder FA_14693(s14693, c14693, in14693_1, in14693_2, c13902);
    wire[0:0] s14694, in14694_1, in14694_2;
    wire c14694;
    assign in14694_1 = {c13904};
    assign in14694_2 = {c13905};
    Full_Adder FA_14694(s14694, c14694, in14694_1, in14694_2, c13903);
    wire[0:0] s14695, in14695_1, in14695_2;
    wire c14695;
    assign in14695_1 = {s13907[0]};
    assign in14695_2 = {s13908[0]};
    Full_Adder FA_14695(s14695, c14695, in14695_1, in14695_2, c13906);
    wire[0:0] s14696, in14696_1, in14696_2;
    wire c14696;
    assign in14696_1 = {c13908};
    assign in14696_2 = {c13909};
    Full_Adder FA_14696(s14696, c14696, in14696_1, in14696_2, c13907);
    wire[0:0] s14697, in14697_1, in14697_2;
    wire c14697;
    assign in14697_1 = {s13911[0]};
    assign in14697_2 = {s13912[0]};
    Full_Adder FA_14697(s14697, c14697, in14697_1, in14697_2, c13910);
    wire[0:0] s14698, in14698_1, in14698_2;
    wire c14698;
    assign in14698_1 = {c13912};
    assign in14698_2 = {c13913};
    Full_Adder FA_14698(s14698, c14698, in14698_1, in14698_2, c13911);
    wire[0:0] s14699, in14699_1, in14699_2;
    wire c14699;
    assign in14699_1 = {s13915[0]};
    assign in14699_2 = {s13916[0]};
    Full_Adder FA_14699(s14699, c14699, in14699_1, in14699_2, c13914);
    wire[0:0] s14700, in14700_1, in14700_2;
    wire c14700;
    assign in14700_1 = {c13916};
    assign in14700_2 = {c13917};
    Full_Adder FA_14700(s14700, c14700, in14700_1, in14700_2, c13915);
    wire[0:0] s14701, in14701_1, in14701_2;
    wire c14701;
    assign in14701_1 = {s13919[0]};
    assign in14701_2 = {s13920[0]};
    Full_Adder FA_14701(s14701, c14701, in14701_1, in14701_2, c13918);
    wire[0:0] s14702, in14702_1, in14702_2;
    wire c14702;
    assign in14702_1 = {c13920};
    assign in14702_2 = {c13921};
    Full_Adder FA_14702(s14702, c14702, in14702_1, in14702_2, c13919);
    wire[0:0] s14703, in14703_1, in14703_2;
    wire c14703;
    assign in14703_1 = {s13923[0]};
    assign in14703_2 = {s13924[0]};
    Full_Adder FA_14703(s14703, c14703, in14703_1, in14703_2, c13922);
    wire[0:0] s14704, in14704_1, in14704_2;
    wire c14704;
    assign in14704_1 = {c13924};
    assign in14704_2 = {c13925};
    Full_Adder FA_14704(s14704, c14704, in14704_1, in14704_2, c13923);
    wire[0:0] s14705, in14705_1, in14705_2;
    wire c14705;
    assign in14705_1 = {s13927[0]};
    assign in14705_2 = {s13928[0]};
    Full_Adder FA_14705(s14705, c14705, in14705_1, in14705_2, c13926);
    wire[0:0] s14706, in14706_1, in14706_2;
    wire c14706;
    assign in14706_1 = {c13928};
    assign in14706_2 = {c13929};
    Full_Adder FA_14706(s14706, c14706, in14706_1, in14706_2, c13927);
    wire[0:0] s14707, in14707_1, in14707_2;
    wire c14707;
    assign in14707_1 = {s13931[0]};
    assign in14707_2 = {s13932[0]};
    Full_Adder FA_14707(s14707, c14707, in14707_1, in14707_2, c13930);
    wire[0:0] s14708, in14708_1, in14708_2;
    wire c14708;
    assign in14708_1 = {c13932};
    assign in14708_2 = {c13933};
    Full_Adder FA_14708(s14708, c14708, in14708_1, in14708_2, c13931);
    wire[0:0] s14709, in14709_1, in14709_2;
    wire c14709;
    assign in14709_1 = {s13935[0]};
    assign in14709_2 = {s13936[0]};
    Full_Adder FA_14709(s14709, c14709, in14709_1, in14709_2, c13934);
    wire[0:0] s14710, in14710_1, in14710_2;
    wire c14710;
    assign in14710_1 = {c13936};
    assign in14710_2 = {c13937};
    Full_Adder FA_14710(s14710, c14710, in14710_1, in14710_2, c13935);
    wire[0:0] s14711, in14711_1, in14711_2;
    wire c14711;
    assign in14711_1 = {s13939[0]};
    assign in14711_2 = {s13940[0]};
    Full_Adder FA_14711(s14711, c14711, in14711_1, in14711_2, c13938);
    wire[0:0] s14712, in14712_1, in14712_2;
    wire c14712;
    assign in14712_1 = {c13940};
    assign in14712_2 = {c13941};
    Full_Adder FA_14712(s14712, c14712, in14712_1, in14712_2, c13939);
    wire[0:0] s14713, in14713_1, in14713_2;
    wire c14713;
    assign in14713_1 = {s13943[0]};
    assign in14713_2 = {s13944[0]};
    Full_Adder FA_14713(s14713, c14713, in14713_1, in14713_2, c13942);
    wire[0:0] s14714, in14714_1, in14714_2;
    wire c14714;
    assign in14714_1 = {c13944};
    assign in14714_2 = {c13945};
    Full_Adder FA_14714(s14714, c14714, in14714_1, in14714_2, c13943);
    wire[0:0] s14715, in14715_1, in14715_2;
    wire c14715;
    assign in14715_1 = {s13947[0]};
    assign in14715_2 = {s13948[0]};
    Full_Adder FA_14715(s14715, c14715, in14715_1, in14715_2, c13946);
    wire[0:0] s14716, in14716_1, in14716_2;
    wire c14716;
    assign in14716_1 = {c13948};
    assign in14716_2 = {c13949};
    Full_Adder FA_14716(s14716, c14716, in14716_1, in14716_2, c13947);
    wire[0:0] s14717, in14717_1, in14717_2;
    wire c14717;
    assign in14717_1 = {s13951[0]};
    assign in14717_2 = {s13952[0]};
    Full_Adder FA_14717(s14717, c14717, in14717_1, in14717_2, c13950);
    wire[0:0] s14718, in14718_1, in14718_2;
    wire c14718;
    assign in14718_1 = {c13952};
    assign in14718_2 = {c13953};
    Full_Adder FA_14718(s14718, c14718, in14718_1, in14718_2, c13951);
    wire[0:0] s14719, in14719_1, in14719_2;
    wire c14719;
    assign in14719_1 = {s13955[0]};
    assign in14719_2 = {s13956[0]};
    Full_Adder FA_14719(s14719, c14719, in14719_1, in14719_2, c13954);
    wire[0:0] s14720, in14720_1, in14720_2;
    wire c14720;
    assign in14720_1 = {c13956};
    assign in14720_2 = {c13957};
    Full_Adder FA_14720(s14720, c14720, in14720_1, in14720_2, c13955);
    wire[0:0] s14721, in14721_1, in14721_2;
    wire c14721;
    assign in14721_1 = {s13959[0]};
    assign in14721_2 = {s13960[0]};
    Full_Adder FA_14721(s14721, c14721, in14721_1, in14721_2, c13958);
    wire[0:0] s14722, in14722_1, in14722_2;
    wire c14722;
    assign in14722_1 = {c13960};
    assign in14722_2 = {c13961};
    Full_Adder FA_14722(s14722, c14722, in14722_1, in14722_2, c13959);
    wire[0:0] s14723, in14723_1, in14723_2;
    wire c14723;
    assign in14723_1 = {s13963[0]};
    assign in14723_2 = {s13964[0]};
    Full_Adder FA_14723(s14723, c14723, in14723_1, in14723_2, c13962);
    wire[0:0] s14724, in14724_1, in14724_2;
    wire c14724;
    assign in14724_1 = {c13964};
    assign in14724_2 = {c13965};
    Full_Adder FA_14724(s14724, c14724, in14724_1, in14724_2, c13963);
    wire[0:0] s14725, in14725_1, in14725_2;
    wire c14725;
    assign in14725_1 = {s13967[0]};
    assign in14725_2 = {s13968[0]};
    Full_Adder FA_14725(s14725, c14725, in14725_1, in14725_2, c13966);
    wire[0:0] s14726, in14726_1, in14726_2;
    wire c14726;
    assign in14726_1 = {c13968};
    assign in14726_2 = {c13969};
    Full_Adder FA_14726(s14726, c14726, in14726_1, in14726_2, c13967);
    wire[0:0] s14727, in14727_1, in14727_2;
    wire c14727;
    assign in14727_1 = {s13971[0]};
    assign in14727_2 = {s13972[0]};
    Full_Adder FA_14727(s14727, c14727, in14727_1, in14727_2, c13970);
    wire[0:0] s14728, in14728_1, in14728_2;
    wire c14728;
    assign in14728_1 = {c13972};
    assign in14728_2 = {c13973};
    Full_Adder FA_14728(s14728, c14728, in14728_1, in14728_2, c13971);
    wire[0:0] s14729, in14729_1, in14729_2;
    wire c14729;
    assign in14729_1 = {s13975[0]};
    assign in14729_2 = {s13976[0]};
    Full_Adder FA_14729(s14729, c14729, in14729_1, in14729_2, c13974);
    wire[0:0] s14730, in14730_1, in14730_2;
    wire c14730;
    assign in14730_1 = {c13976};
    assign in14730_2 = {c13977};
    Full_Adder FA_14730(s14730, c14730, in14730_1, in14730_2, c13975);
    wire[0:0] s14731, in14731_1, in14731_2;
    wire c14731;
    assign in14731_1 = {s13979[0]};
    assign in14731_2 = {s13980[0]};
    Full_Adder FA_14731(s14731, c14731, in14731_1, in14731_2, c13978);
    wire[0:0] s14732, in14732_1, in14732_2;
    wire c14732;
    assign in14732_1 = {c13980};
    assign in14732_2 = {c13981};
    Full_Adder FA_14732(s14732, c14732, in14732_1, in14732_2, c13979);
    wire[0:0] s14733, in14733_1, in14733_2;
    wire c14733;
    assign in14733_1 = {s13983[0]};
    assign in14733_2 = {s13984[0]};
    Full_Adder FA_14733(s14733, c14733, in14733_1, in14733_2, c13982);
    wire[0:0] s14734, in14734_1, in14734_2;
    wire c14734;
    assign in14734_1 = {c13984};
    assign in14734_2 = {c13985};
    Full_Adder FA_14734(s14734, c14734, in14734_1, in14734_2, c13983);
    wire[0:0] s14735, in14735_1, in14735_2;
    wire c14735;
    assign in14735_1 = {s13987[0]};
    assign in14735_2 = {s13988[0]};
    Full_Adder FA_14735(s14735, c14735, in14735_1, in14735_2, c13986);
    wire[0:0] s14736, in14736_1, in14736_2;
    wire c14736;
    assign in14736_1 = {c13988};
    assign in14736_2 = {c13989};
    Full_Adder FA_14736(s14736, c14736, in14736_1, in14736_2, c13987);
    wire[0:0] s14737, in14737_1, in14737_2;
    wire c14737;
    assign in14737_1 = {s13991[0]};
    assign in14737_2 = {s13992[0]};
    Full_Adder FA_14737(s14737, c14737, in14737_1, in14737_2, c13990);
    wire[0:0] s14738, in14738_1, in14738_2;
    wire c14738;
    assign in14738_1 = {c13992};
    assign in14738_2 = {c13993};
    Full_Adder FA_14738(s14738, c14738, in14738_1, in14738_2, c13991);
    wire[0:0] s14739, in14739_1, in14739_2;
    wire c14739;
    assign in14739_1 = {s13995[0]};
    assign in14739_2 = {s13996[0]};
    Full_Adder FA_14739(s14739, c14739, in14739_1, in14739_2, c13994);
    wire[0:0] s14740, in14740_1, in14740_2;
    wire c14740;
    assign in14740_1 = {c13996};
    assign in14740_2 = {c13997};
    Full_Adder FA_14740(s14740, c14740, in14740_1, in14740_2, c13995);
    wire[0:0] s14741, in14741_1, in14741_2;
    wire c14741;
    assign in14741_1 = {s13999[0]};
    assign in14741_2 = {s14000[0]};
    Full_Adder FA_14741(s14741, c14741, in14741_1, in14741_2, c13998);
    wire[0:0] s14742, in14742_1, in14742_2;
    wire c14742;
    assign in14742_1 = {c14000};
    assign in14742_2 = {c14001};
    Full_Adder FA_14742(s14742, c14742, in14742_1, in14742_2, c13999);
    wire[0:0] s14743, in14743_1, in14743_2;
    wire c14743;
    assign in14743_1 = {s14003[0]};
    assign in14743_2 = {s14004[0]};
    Full_Adder FA_14743(s14743, c14743, in14743_1, in14743_2, c14002);
    wire[0:0] s14744, in14744_1, in14744_2;
    wire c14744;
    assign in14744_1 = {c14004};
    assign in14744_2 = {c14005};
    Full_Adder FA_14744(s14744, c14744, in14744_1, in14744_2, c14003);
    wire[0:0] s14745, in14745_1, in14745_2;
    wire c14745;
    assign in14745_1 = {s14007[0]};
    assign in14745_2 = {s14008[0]};
    Full_Adder FA_14745(s14745, c14745, in14745_1, in14745_2, c14006);
    wire[0:0] s14746, in14746_1, in14746_2;
    wire c14746;
    assign in14746_1 = {c14008};
    assign in14746_2 = {c14009};
    Full_Adder FA_14746(s14746, c14746, in14746_1, in14746_2, c14007);
    wire[0:0] s14747, in14747_1, in14747_2;
    wire c14747;
    assign in14747_1 = {s14011[0]};
    assign in14747_2 = {s14012[0]};
    Full_Adder FA_14747(s14747, c14747, in14747_1, in14747_2, c14010);
    wire[0:0] s14748, in14748_1, in14748_2;
    wire c14748;
    assign in14748_1 = {c14012};
    assign in14748_2 = {c14013};
    Full_Adder FA_14748(s14748, c14748, in14748_1, in14748_2, c14011);
    wire[0:0] s14749, in14749_1, in14749_2;
    wire c14749;
    assign in14749_1 = {s14015[0]};
    assign in14749_2 = {s14016[0]};
    Full_Adder FA_14749(s14749, c14749, in14749_1, in14749_2, c14014);
    wire[0:0] s14750, in14750_1, in14750_2;
    wire c14750;
    assign in14750_1 = {c14016};
    assign in14750_2 = {c14017};
    Full_Adder FA_14750(s14750, c14750, in14750_1, in14750_2, c14015);
    wire[0:0] s14751, in14751_1, in14751_2;
    wire c14751;
    assign in14751_1 = {s14019[0]};
    assign in14751_2 = {s14020[0]};
    Full_Adder FA_14751(s14751, c14751, in14751_1, in14751_2, c14018);
    wire[0:0] s14752, in14752_1, in14752_2;
    wire c14752;
    assign in14752_1 = {c14020};
    assign in14752_2 = {c14021};
    Full_Adder FA_14752(s14752, c14752, in14752_1, in14752_2, c14019);
    wire[0:0] s14753, in14753_1, in14753_2;
    wire c14753;
    assign in14753_1 = {s14023[0]};
    assign in14753_2 = {s14024[0]};
    Full_Adder FA_14753(s14753, c14753, in14753_1, in14753_2, c14022);
    wire[0:0] s14754, in14754_1, in14754_2;
    wire c14754;
    assign in14754_1 = {c14024};
    assign in14754_2 = {c14025};
    Full_Adder FA_14754(s14754, c14754, in14754_1, in14754_2, c14023);
    wire[0:0] s14755, in14755_1, in14755_2;
    wire c14755;
    assign in14755_1 = {s14027[0]};
    assign in14755_2 = {s14028[0]};
    Full_Adder FA_14755(s14755, c14755, in14755_1, in14755_2, c14026);
    wire[0:0] s14756, in14756_1, in14756_2;
    wire c14756;
    assign in14756_1 = {c14028};
    assign in14756_2 = {c14029};
    Full_Adder FA_14756(s14756, c14756, in14756_1, in14756_2, c14027);
    wire[0:0] s14757, in14757_1, in14757_2;
    wire c14757;
    assign in14757_1 = {s14031[0]};
    assign in14757_2 = {s14032[0]};
    Full_Adder FA_14757(s14757, c14757, in14757_1, in14757_2, c14030);
    wire[0:0] s14758, in14758_1, in14758_2;
    wire c14758;
    assign in14758_1 = {c14032};
    assign in14758_2 = {c14033};
    Full_Adder FA_14758(s14758, c14758, in14758_1, in14758_2, c14031);
    wire[0:0] s14759, in14759_1, in14759_2;
    wire c14759;
    assign in14759_1 = {s14035[0]};
    assign in14759_2 = {s14036[0]};
    Full_Adder FA_14759(s14759, c14759, in14759_1, in14759_2, c14034);
    wire[0:0] s14760, in14760_1, in14760_2;
    wire c14760;
    assign in14760_1 = {c14036};
    assign in14760_2 = {c14037};
    Full_Adder FA_14760(s14760, c14760, in14760_1, in14760_2, c14035);
    wire[0:0] s14761, in14761_1, in14761_2;
    wire c14761;
    assign in14761_1 = {s14039[0]};
    assign in14761_2 = {s14040[0]};
    Full_Adder FA_14761(s14761, c14761, in14761_1, in14761_2, c14038);
    wire[0:0] s14762, in14762_1, in14762_2;
    wire c14762;
    assign in14762_1 = {c14040};
    assign in14762_2 = {c14041};
    Full_Adder FA_14762(s14762, c14762, in14762_1, in14762_2, c14039);
    wire[0:0] s14763, in14763_1, in14763_2;
    wire c14763;
    assign in14763_1 = {s14043[0]};
    assign in14763_2 = {s14044[0]};
    Full_Adder FA_14763(s14763, c14763, in14763_1, in14763_2, c14042);
    wire[0:0] s14764, in14764_1, in14764_2;
    wire c14764;
    assign in14764_1 = {c14044};
    assign in14764_2 = {c14045};
    Full_Adder FA_14764(s14764, c14764, in14764_1, in14764_2, c14043);
    wire[0:0] s14765, in14765_1, in14765_2;
    wire c14765;
    assign in14765_1 = {s14047[0]};
    assign in14765_2 = {s14048[0]};
    Full_Adder FA_14765(s14765, c14765, in14765_1, in14765_2, c14046);
    wire[0:0] s14766, in14766_1, in14766_2;
    wire c14766;
    assign in14766_1 = {c14048};
    assign in14766_2 = {c14049};
    Full_Adder FA_14766(s14766, c14766, in14766_1, in14766_2, c14047);
    wire[0:0] s14767, in14767_1, in14767_2;
    wire c14767;
    assign in14767_1 = {s14051[0]};
    assign in14767_2 = {s14052[0]};
    Full_Adder FA_14767(s14767, c14767, in14767_1, in14767_2, c14050);
    wire[0:0] s14768, in14768_1, in14768_2;
    wire c14768;
    assign in14768_1 = {c14052};
    assign in14768_2 = {c14053};
    Full_Adder FA_14768(s14768, c14768, in14768_1, in14768_2, c14051);
    wire[0:0] s14769, in14769_1, in14769_2;
    wire c14769;
    assign in14769_1 = {s14055[0]};
    assign in14769_2 = {s14056[0]};
    Full_Adder FA_14769(s14769, c14769, in14769_1, in14769_2, c14054);
    wire[0:0] s14770, in14770_1, in14770_2;
    wire c14770;
    assign in14770_1 = {c14056};
    assign in14770_2 = {c14057};
    Full_Adder FA_14770(s14770, c14770, in14770_1, in14770_2, c14055);
    wire[0:0] s14771, in14771_1, in14771_2;
    wire c14771;
    assign in14771_1 = {s14059[0]};
    assign in14771_2 = {s14060[0]};
    Full_Adder FA_14771(s14771, c14771, in14771_1, in14771_2, c14058);
    wire[0:0] s14772, in14772_1, in14772_2;
    wire c14772;
    assign in14772_1 = {c14060};
    assign in14772_2 = {c14061};
    Full_Adder FA_14772(s14772, c14772, in14772_1, in14772_2, c14059);
    wire[0:0] s14773, in14773_1, in14773_2;
    wire c14773;
    assign in14773_1 = {s14063[0]};
    assign in14773_2 = {s14064[0]};
    Full_Adder FA_14773(s14773, c14773, in14773_1, in14773_2, c14062);
    wire[0:0] s14774, in14774_1, in14774_2;
    wire c14774;
    assign in14774_1 = {c14064};
    assign in14774_2 = {c14065};
    Full_Adder FA_14774(s14774, c14774, in14774_1, in14774_2, c14063);
    wire[0:0] s14775, in14775_1, in14775_2;
    wire c14775;
    assign in14775_1 = {s14067[0]};
    assign in14775_2 = {s14068[0]};
    Full_Adder FA_14775(s14775, c14775, in14775_1, in14775_2, c14066);
    wire[0:0] s14776, in14776_1, in14776_2;
    wire c14776;
    assign in14776_1 = {c14068};
    assign in14776_2 = {c14069};
    Full_Adder FA_14776(s14776, c14776, in14776_1, in14776_2, c14067);
    wire[0:0] s14777, in14777_1, in14777_2;
    wire c14777;
    assign in14777_1 = {s14071[0]};
    assign in14777_2 = {s14072[0]};
    Full_Adder FA_14777(s14777, c14777, in14777_1, in14777_2, c14070);
    wire[0:0] s14778, in14778_1, in14778_2;
    wire c14778;
    assign in14778_1 = {c14072};
    assign in14778_2 = {c14073};
    Full_Adder FA_14778(s14778, c14778, in14778_1, in14778_2, c14071);
    wire[0:0] s14779, in14779_1, in14779_2;
    wire c14779;
    assign in14779_1 = {s14075[0]};
    assign in14779_2 = {s14076[0]};
    Full_Adder FA_14779(s14779, c14779, in14779_1, in14779_2, c14074);
    wire[0:0] s14780, in14780_1, in14780_2;
    wire c14780;
    assign in14780_1 = {c14076};
    assign in14780_2 = {c14077};
    Full_Adder FA_14780(s14780, c14780, in14780_1, in14780_2, c14075);
    wire[0:0] s14781, in14781_1, in14781_2;
    wire c14781;
    assign in14781_1 = {s14079[0]};
    assign in14781_2 = {s14080[0]};
    Full_Adder FA_14781(s14781, c14781, in14781_1, in14781_2, c14078);
    wire[0:0] s14782, in14782_1, in14782_2;
    wire c14782;
    assign in14782_1 = {c14080};
    assign in14782_2 = {c14081};
    Full_Adder FA_14782(s14782, c14782, in14782_1, in14782_2, c14079);
    wire[0:0] s14783, in14783_1, in14783_2;
    wire c14783;
    assign in14783_1 = {s14083[0]};
    assign in14783_2 = {s14084[0]};
    Full_Adder FA_14783(s14783, c14783, in14783_1, in14783_2, c14082);
    wire[0:0] s14784, in14784_1, in14784_2;
    wire c14784;
    assign in14784_1 = {c14084};
    assign in14784_2 = {c14085};
    Full_Adder FA_14784(s14784, c14784, in14784_1, in14784_2, c14083);
    wire[0:0] s14785, in14785_1, in14785_2;
    wire c14785;
    assign in14785_1 = {s14087[0]};
    assign in14785_2 = {s14088[0]};
    Full_Adder FA_14785(s14785, c14785, in14785_1, in14785_2, c14086);
    wire[0:0] s14786, in14786_1, in14786_2;
    wire c14786;
    assign in14786_1 = {c14088};
    assign in14786_2 = {c14089};
    Full_Adder FA_14786(s14786, c14786, in14786_1, in14786_2, c14087);
    wire[0:0] s14787, in14787_1, in14787_2;
    wire c14787;
    assign in14787_1 = {s14091[0]};
    assign in14787_2 = {s14092[0]};
    Full_Adder FA_14787(s14787, c14787, in14787_1, in14787_2, c14090);
    wire[0:0] s14788, in14788_1, in14788_2;
    wire c14788;
    assign in14788_1 = {c14092};
    assign in14788_2 = {c14093};
    Full_Adder FA_14788(s14788, c14788, in14788_1, in14788_2, c14091);
    wire[0:0] s14789, in14789_1, in14789_2;
    wire c14789;
    assign in14789_1 = {s14095[0]};
    assign in14789_2 = {s14096[0]};
    Full_Adder FA_14789(s14789, c14789, in14789_1, in14789_2, c14094);
    wire[0:0] s14790, in14790_1, in14790_2;
    wire c14790;
    assign in14790_1 = {c14096};
    assign in14790_2 = {c14097};
    Full_Adder FA_14790(s14790, c14790, in14790_1, in14790_2, c14095);
    wire[0:0] s14791, in14791_1, in14791_2;
    wire c14791;
    assign in14791_1 = {s14099[0]};
    assign in14791_2 = {s14100[0]};
    Full_Adder FA_14791(s14791, c14791, in14791_1, in14791_2, c14098);
    wire[0:0] s14792, in14792_1, in14792_2;
    wire c14792;
    assign in14792_1 = {c14100};
    assign in14792_2 = {c14101};
    Full_Adder FA_14792(s14792, c14792, in14792_1, in14792_2, c14099);
    wire[0:0] s14793, in14793_1, in14793_2;
    wire c14793;
    assign in14793_1 = {s14103[0]};
    assign in14793_2 = {s14104[0]};
    Full_Adder FA_14793(s14793, c14793, in14793_1, in14793_2, c14102);
    wire[0:0] s14794, in14794_1, in14794_2;
    wire c14794;
    assign in14794_1 = {c14104};
    assign in14794_2 = {c14105};
    Full_Adder FA_14794(s14794, c14794, in14794_1, in14794_2, c14103);
    wire[0:0] s14795, in14795_1, in14795_2;
    wire c14795;
    assign in14795_1 = {s14107[0]};
    assign in14795_2 = {s14108[0]};
    Full_Adder FA_14795(s14795, c14795, in14795_1, in14795_2, c14106);
    wire[0:0] s14796, in14796_1, in14796_2;
    wire c14796;
    assign in14796_1 = {c14108};
    assign in14796_2 = {c14109};
    Full_Adder FA_14796(s14796, c14796, in14796_1, in14796_2, c14107);
    wire[0:0] s14797, in14797_1, in14797_2;
    wire c14797;
    assign in14797_1 = {s14111[0]};
    assign in14797_2 = {s14112[0]};
    Full_Adder FA_14797(s14797, c14797, in14797_1, in14797_2, c14110);
    wire[0:0] s14798, in14798_1, in14798_2;
    wire c14798;
    assign in14798_1 = {c14112};
    assign in14798_2 = {c14113};
    Full_Adder FA_14798(s14798, c14798, in14798_1, in14798_2, c14111);
    wire[0:0] s14799, in14799_1, in14799_2;
    wire c14799;
    assign in14799_1 = {s14115[0]};
    assign in14799_2 = {s14116[0]};
    Full_Adder FA_14799(s14799, c14799, in14799_1, in14799_2, c14114);
    wire[0:0] s14800, in14800_1, in14800_2;
    wire c14800;
    assign in14800_1 = {c14116};
    assign in14800_2 = {c14117};
    Full_Adder FA_14800(s14800, c14800, in14800_1, in14800_2, c14115);
    wire[0:0] s14801, in14801_1, in14801_2;
    wire c14801;
    assign in14801_1 = {s14119[0]};
    assign in14801_2 = {s14120[0]};
    Full_Adder FA_14801(s14801, c14801, in14801_1, in14801_2, c14118);
    wire[0:0] s14802, in14802_1, in14802_2;
    wire c14802;
    assign in14802_1 = {c14120};
    assign in14802_2 = {c14121};
    Full_Adder FA_14802(s14802, c14802, in14802_1, in14802_2, c14119);
    wire[0:0] s14803, in14803_1, in14803_2;
    wire c14803;
    assign in14803_1 = {s14123[0]};
    assign in14803_2 = {s14124[0]};
    Full_Adder FA_14803(s14803, c14803, in14803_1, in14803_2, c14122);
    wire[0:0] s14804, in14804_1, in14804_2;
    wire c14804;
    assign in14804_1 = {c14124};
    assign in14804_2 = {c14125};
    Full_Adder FA_14804(s14804, c14804, in14804_1, in14804_2, c14123);
    wire[0:0] s14805, in14805_1, in14805_2;
    wire c14805;
    assign in14805_1 = {s14127[0]};
    assign in14805_2 = {s14128[0]};
    Full_Adder FA_14805(s14805, c14805, in14805_1, in14805_2, c14126);
    wire[0:0] s14806, in14806_1, in14806_2;
    wire c14806;
    assign in14806_1 = {c14128};
    assign in14806_2 = {c14129};
    Full_Adder FA_14806(s14806, c14806, in14806_1, in14806_2, c14127);
    wire[0:0] s14807, in14807_1, in14807_2;
    wire c14807;
    assign in14807_1 = {s14131[0]};
    assign in14807_2 = {s14132[0]};
    Full_Adder FA_14807(s14807, c14807, in14807_1, in14807_2, c14130);
    wire[0:0] s14808, in14808_1, in14808_2;
    wire c14808;
    assign in14808_1 = {c14132};
    assign in14808_2 = {c14133};
    Full_Adder FA_14808(s14808, c14808, in14808_1, in14808_2, c14131);
    wire[0:0] s14809, in14809_1, in14809_2;
    wire c14809;
    assign in14809_1 = {s14135[0]};
    assign in14809_2 = {s14136[0]};
    Full_Adder FA_14809(s14809, c14809, in14809_1, in14809_2, c14134);
    wire[0:0] s14810, in14810_1, in14810_2;
    wire c14810;
    assign in14810_1 = {c14136};
    assign in14810_2 = {c14137};
    Full_Adder FA_14810(s14810, c14810, in14810_1, in14810_2, c14135);
    wire[0:0] s14811, in14811_1, in14811_2;
    wire c14811;
    assign in14811_1 = {s14139[0]};
    assign in14811_2 = {s14140[0]};
    Full_Adder FA_14811(s14811, c14811, in14811_1, in14811_2, c14138);
    wire[0:0] s14812, in14812_1, in14812_2;
    wire c14812;
    assign in14812_1 = {c14140};
    assign in14812_2 = {c14141};
    Full_Adder FA_14812(s14812, c14812, in14812_1, in14812_2, c14139);
    wire[0:0] s14813, in14813_1, in14813_2;
    wire c14813;
    assign in14813_1 = {s14143[0]};
    assign in14813_2 = {s14144[0]};
    Full_Adder FA_14813(s14813, c14813, in14813_1, in14813_2, c14142);
    wire[0:0] s14814, in14814_1, in14814_2;
    wire c14814;
    assign in14814_1 = {c14144};
    assign in14814_2 = {c14145};
    Full_Adder FA_14814(s14814, c14814, in14814_1, in14814_2, c14143);
    wire[0:0] s14815, in14815_1, in14815_2;
    wire c14815;
    assign in14815_1 = {s14147[0]};
    assign in14815_2 = {s14148[0]};
    Full_Adder FA_14815(s14815, c14815, in14815_1, in14815_2, c14146);
    wire[0:0] s14816, in14816_1, in14816_2;
    wire c14816;
    assign in14816_1 = {c14148};
    assign in14816_2 = {c14149};
    Full_Adder FA_14816(s14816, c14816, in14816_1, in14816_2, c14147);
    wire[0:0] s14817, in14817_1, in14817_2;
    wire c14817;
    assign in14817_1 = {s14151[0]};
    assign in14817_2 = {s14152[0]};
    Full_Adder FA_14817(s14817, c14817, in14817_1, in14817_2, c14150);
    wire[0:0] s14818, in14818_1, in14818_2;
    wire c14818;
    assign in14818_1 = {c14152};
    assign in14818_2 = {c14153};
    Full_Adder FA_14818(s14818, c14818, in14818_1, in14818_2, c14151);
    wire[0:0] s14819, in14819_1, in14819_2;
    wire c14819;
    assign in14819_1 = {s14155[0]};
    assign in14819_2 = {s14156[0]};
    Full_Adder FA_14819(s14819, c14819, in14819_1, in14819_2, c14154);
    wire[0:0] s14820, in14820_1, in14820_2;
    wire c14820;
    assign in14820_1 = {c14156};
    assign in14820_2 = {c14157};
    Full_Adder FA_14820(s14820, c14820, in14820_1, in14820_2, c14155);
    wire[0:0] s14821, in14821_1, in14821_2;
    wire c14821;
    assign in14821_1 = {s14159[0]};
    assign in14821_2 = {s14160[0]};
    Full_Adder FA_14821(s14821, c14821, in14821_1, in14821_2, c14158);
    wire[0:0] s14822, in14822_1, in14822_2;
    wire c14822;
    assign in14822_1 = {c14160};
    assign in14822_2 = {c14161};
    Full_Adder FA_14822(s14822, c14822, in14822_1, in14822_2, c14159);
    wire[0:0] s14823, in14823_1, in14823_2;
    wire c14823;
    assign in14823_1 = {s14163[0]};
    assign in14823_2 = {s14164[0]};
    Full_Adder FA_14823(s14823, c14823, in14823_1, in14823_2, c14162);
    wire[0:0] s14824, in14824_1, in14824_2;
    wire c14824;
    assign in14824_1 = {c14164};
    assign in14824_2 = {c14165};
    Full_Adder FA_14824(s14824, c14824, in14824_1, in14824_2, c14163);
    wire[0:0] s14825, in14825_1, in14825_2;
    wire c14825;
    assign in14825_1 = {s14167[0]};
    assign in14825_2 = {s14168[0]};
    Full_Adder FA_14825(s14825, c14825, in14825_1, in14825_2, c14166);
    wire[0:0] s14826, in14826_1, in14826_2;
    wire c14826;
    assign in14826_1 = {c14168};
    assign in14826_2 = {c14169};
    Full_Adder FA_14826(s14826, c14826, in14826_1, in14826_2, c14167);
    wire[0:0] s14827, in14827_1, in14827_2;
    wire c14827;
    assign in14827_1 = {s14171[0]};
    assign in14827_2 = {s14172[0]};
    Full_Adder FA_14827(s14827, c14827, in14827_1, in14827_2, c14170);
    wire[0:0] s14828, in14828_1, in14828_2;
    wire c14828;
    assign in14828_1 = {c14172};
    assign in14828_2 = {c14173};
    Full_Adder FA_14828(s14828, c14828, in14828_1, in14828_2, c14171);
    wire[0:0] s14829, in14829_1, in14829_2;
    wire c14829;
    assign in14829_1 = {s14175[0]};
    assign in14829_2 = {s14176[0]};
    Full_Adder FA_14829(s14829, c14829, in14829_1, in14829_2, c14174);
    wire[0:0] s14830, in14830_1, in14830_2;
    wire c14830;
    assign in14830_1 = {c14176};
    assign in14830_2 = {c14177};
    Full_Adder FA_14830(s14830, c14830, in14830_1, in14830_2, c14175);
    wire[0:0] s14831, in14831_1, in14831_2;
    wire c14831;
    assign in14831_1 = {s14179[0]};
    assign in14831_2 = {s14180[0]};
    Full_Adder FA_14831(s14831, c14831, in14831_1, in14831_2, c14178);
    wire[0:0] s14832, in14832_1, in14832_2;
    wire c14832;
    assign in14832_1 = {c14180};
    assign in14832_2 = {c14181};
    Full_Adder FA_14832(s14832, c14832, in14832_1, in14832_2, c14179);
    wire[0:0] s14833, in14833_1, in14833_2;
    wire c14833;
    assign in14833_1 = {s14183[0]};
    assign in14833_2 = {s14184[0]};
    Full_Adder FA_14833(s14833, c14833, in14833_1, in14833_2, c14182);
    wire[0:0] s14834, in14834_1, in14834_2;
    wire c14834;
    assign in14834_1 = {c14184};
    assign in14834_2 = {c14185};
    Full_Adder FA_14834(s14834, c14834, in14834_1, in14834_2, c14183);
    wire[0:0] s14835, in14835_1, in14835_2;
    wire c14835;
    assign in14835_1 = {s14187[0]};
    assign in14835_2 = {s14188[0]};
    Full_Adder FA_14835(s14835, c14835, in14835_1, in14835_2, c14186);
    wire[0:0] s14836, in14836_1, in14836_2;
    wire c14836;
    assign in14836_1 = {c14188};
    assign in14836_2 = {c14189};
    Full_Adder FA_14836(s14836, c14836, in14836_1, in14836_2, c14187);
    wire[0:0] s14837, in14837_1, in14837_2;
    wire c14837;
    assign in14837_1 = {s14191[0]};
    assign in14837_2 = {s14192[0]};
    Full_Adder FA_14837(s14837, c14837, in14837_1, in14837_2, c14190);
    wire[0:0] s14838, in14838_1, in14838_2;
    wire c14838;
    assign in14838_1 = {c14192};
    assign in14838_2 = {c14193};
    Full_Adder FA_14838(s14838, c14838, in14838_1, in14838_2, c14191);
    wire[0:0] s14839, in14839_1, in14839_2;
    wire c14839;
    assign in14839_1 = {s14195[0]};
    assign in14839_2 = {s14196[0]};
    Full_Adder FA_14839(s14839, c14839, in14839_1, in14839_2, c14194);
    wire[0:0] s14840, in14840_1, in14840_2;
    wire c14840;
    assign in14840_1 = {c14196};
    assign in14840_2 = {c14197};
    Full_Adder FA_14840(s14840, c14840, in14840_1, in14840_2, c14195);
    wire[0:0] s14841, in14841_1, in14841_2;
    wire c14841;
    assign in14841_1 = {s14199[0]};
    assign in14841_2 = {s14200[0]};
    Full_Adder FA_14841(s14841, c14841, in14841_1, in14841_2, c14198);
    wire[0:0] s14842, in14842_1, in14842_2;
    wire c14842;
    assign in14842_1 = {c14200};
    assign in14842_2 = {c14201};
    Full_Adder FA_14842(s14842, c14842, in14842_1, in14842_2, c14199);
    wire[0:0] s14843, in14843_1, in14843_2;
    wire c14843;
    assign in14843_1 = {s14203[0]};
    assign in14843_2 = {s14204[0]};
    Full_Adder FA_14843(s14843, c14843, in14843_1, in14843_2, c14202);
    wire[0:0] s14844, in14844_1, in14844_2;
    wire c14844;
    assign in14844_1 = {c14204};
    assign in14844_2 = {c14205};
    Full_Adder FA_14844(s14844, c14844, in14844_1, in14844_2, c14203);
    wire[0:0] s14845, in14845_1, in14845_2;
    wire c14845;
    assign in14845_1 = {s14207[0]};
    assign in14845_2 = {s14208[0]};
    Full_Adder FA_14845(s14845, c14845, in14845_1, in14845_2, c14206);
    wire[0:0] s14846, in14846_1, in14846_2;
    wire c14846;
    assign in14846_1 = {c14208};
    assign in14846_2 = {c14209};
    Full_Adder FA_14846(s14846, c14846, in14846_1, in14846_2, c14207);
    wire[0:0] s14847, in14847_1, in14847_2;
    wire c14847;
    assign in14847_1 = {s14211[0]};
    assign in14847_2 = {s14212[0]};
    Full_Adder FA_14847(s14847, c14847, in14847_1, in14847_2, c14210);
    wire[0:0] s14848, in14848_1, in14848_2;
    wire c14848;
    assign in14848_1 = {c14212};
    assign in14848_2 = {c14213};
    Full_Adder FA_14848(s14848, c14848, in14848_1, in14848_2, c14211);
    wire[0:0] s14849, in14849_1, in14849_2;
    wire c14849;
    assign in14849_1 = {s14215[0]};
    assign in14849_2 = {s14216[0]};
    Full_Adder FA_14849(s14849, c14849, in14849_1, in14849_2, c14214);
    wire[0:0] s14850, in14850_1, in14850_2;
    wire c14850;
    assign in14850_1 = {c14216};
    assign in14850_2 = {c14217};
    Full_Adder FA_14850(s14850, c14850, in14850_1, in14850_2, c14215);
    wire[0:0] s14851, in14851_1, in14851_2;
    wire c14851;
    assign in14851_1 = {s14219[0]};
    assign in14851_2 = {s14220[0]};
    Full_Adder FA_14851(s14851, c14851, in14851_1, in14851_2, c14218);
    wire[0:0] s14852, in14852_1, in14852_2;
    wire c14852;
    assign in14852_1 = {c14220};
    assign in14852_2 = {c14221};
    Full_Adder FA_14852(s14852, c14852, in14852_1, in14852_2, c14219);
    wire[0:0] s14853, in14853_1, in14853_2;
    wire c14853;
    assign in14853_1 = {s14223[0]};
    assign in14853_2 = {s14224[0]};
    Full_Adder FA_14853(s14853, c14853, in14853_1, in14853_2, c14222);
    wire[0:0] s14854, in14854_1, in14854_2;
    wire c14854;
    assign in14854_1 = {c14224};
    assign in14854_2 = {c14225};
    Full_Adder FA_14854(s14854, c14854, in14854_1, in14854_2, c14223);
    wire[0:0] s14855, in14855_1, in14855_2;
    wire c14855;
    assign in14855_1 = {s14227[0]};
    assign in14855_2 = {s14228[0]};
    Full_Adder FA_14855(s14855, c14855, in14855_1, in14855_2, c14226);
    wire[0:0] s14856, in14856_1, in14856_2;
    wire c14856;
    assign in14856_1 = {c14228};
    assign in14856_2 = {c14229};
    Full_Adder FA_14856(s14856, c14856, in14856_1, in14856_2, c14227);
    wire[0:0] s14857, in14857_1, in14857_2;
    wire c14857;
    assign in14857_1 = {s14231[0]};
    assign in14857_2 = {s14232[0]};
    Full_Adder FA_14857(s14857, c14857, in14857_1, in14857_2, c14230);
    wire[0:0] s14858, in14858_1, in14858_2;
    wire c14858;
    assign in14858_1 = {c14232};
    assign in14858_2 = {c14233};
    Full_Adder FA_14858(s14858, c14858, in14858_1, in14858_2, c14231);
    wire[0:0] s14859, in14859_1, in14859_2;
    wire c14859;
    assign in14859_1 = {s14235[0]};
    assign in14859_2 = {s14236[0]};
    Full_Adder FA_14859(s14859, c14859, in14859_1, in14859_2, c14234);
    wire[0:0] s14860, in14860_1, in14860_2;
    wire c14860;
    assign in14860_1 = {c14236};
    assign in14860_2 = {c14237};
    Full_Adder FA_14860(s14860, c14860, in14860_1, in14860_2, c14235);
    wire[0:0] s14861, in14861_1, in14861_2;
    wire c14861;
    assign in14861_1 = {s14239[0]};
    assign in14861_2 = {s14240[0]};
    Full_Adder FA_14861(s14861, c14861, in14861_1, in14861_2, c14238);
    wire[0:0] s14862, in14862_1, in14862_2;
    wire c14862;
    assign in14862_1 = {c14240};
    assign in14862_2 = {c14241};
    Full_Adder FA_14862(s14862, c14862, in14862_1, in14862_2, c14239);
    wire[0:0] s14863, in14863_1, in14863_2;
    wire c14863;
    assign in14863_1 = {s14243[0]};
    assign in14863_2 = {s14244[0]};
    Full_Adder FA_14863(s14863, c14863, in14863_1, in14863_2, c14242);
    wire[0:0] s14864, in14864_1, in14864_2;
    wire c14864;
    assign in14864_1 = {c14244};
    assign in14864_2 = {c14245};
    Full_Adder FA_14864(s14864, c14864, in14864_1, in14864_2, c14243);
    wire[0:0] s14865, in14865_1, in14865_2;
    wire c14865;
    assign in14865_1 = {s14247[0]};
    assign in14865_2 = {s14248[0]};
    Full_Adder FA_14865(s14865, c14865, in14865_1, in14865_2, c14246);
    wire[0:0] s14866, in14866_1, in14866_2;
    wire c14866;
    assign in14866_1 = {c14248};
    assign in14866_2 = {c14249};
    Full_Adder FA_14866(s14866, c14866, in14866_1, in14866_2, c14247);
    wire[0:0] s14867, in14867_1, in14867_2;
    wire c14867;
    assign in14867_1 = {s14251[0]};
    assign in14867_2 = {s14252[0]};
    Full_Adder FA_14867(s14867, c14867, in14867_1, in14867_2, c14250);
    wire[0:0] s14868, in14868_1, in14868_2;
    wire c14868;
    assign in14868_1 = {c14252};
    assign in14868_2 = {c14253};
    Full_Adder FA_14868(s14868, c14868, in14868_1, in14868_2, c14251);
    wire[0:0] s14869, in14869_1, in14869_2;
    wire c14869;
    assign in14869_1 = {s14255[0]};
    assign in14869_2 = {s14256[0]};
    Full_Adder FA_14869(s14869, c14869, in14869_1, in14869_2, c14254);
    wire[0:0] s14870, in14870_1, in14870_2;
    wire c14870;
    assign in14870_1 = {c14256};
    assign in14870_2 = {c14257};
    Full_Adder FA_14870(s14870, c14870, in14870_1, in14870_2, c14255);
    wire[0:0] s14871, in14871_1, in14871_2;
    wire c14871;
    assign in14871_1 = {s14259[0]};
    assign in14871_2 = {s14260[0]};
    Full_Adder FA_14871(s14871, c14871, in14871_1, in14871_2, c14258);
    wire[0:0] s14872, in14872_1, in14872_2;
    wire c14872;
    assign in14872_1 = {c14260};
    assign in14872_2 = {c14261};
    Full_Adder FA_14872(s14872, c14872, in14872_1, in14872_2, c14259);
    wire[0:0] s14873, in14873_1, in14873_2;
    wire c14873;
    assign in14873_1 = {s14263[0]};
    assign in14873_2 = {s14264[0]};
    Full_Adder FA_14873(s14873, c14873, in14873_1, in14873_2, c14262);
    wire[0:0] s14874, in14874_1, in14874_2;
    wire c14874;
    assign in14874_1 = {c14264};
    assign in14874_2 = {c14265};
    Full_Adder FA_14874(s14874, c14874, in14874_1, in14874_2, c14263);
    wire[0:0] s14875, in14875_1, in14875_2;
    wire c14875;
    assign in14875_1 = {s14267[0]};
    assign in14875_2 = {s14268[0]};
    Full_Adder FA_14875(s14875, c14875, in14875_1, in14875_2, c14266);
    wire[0:0] s14876, in14876_1, in14876_2;
    wire c14876;
    assign in14876_1 = {c14268};
    assign in14876_2 = {c14269};
    Full_Adder FA_14876(s14876, c14876, in14876_1, in14876_2, c14267);
    wire[0:0] s14877, in14877_1, in14877_2;
    wire c14877;
    assign in14877_1 = {s14271[0]};
    assign in14877_2 = {s14272[0]};
    Full_Adder FA_14877(s14877, c14877, in14877_1, in14877_2, c14270);
    wire[0:0] s14878, in14878_1, in14878_2;
    wire c14878;
    assign in14878_1 = {c14272};
    assign in14878_2 = {c14273};
    Full_Adder FA_14878(s14878, c14878, in14878_1, in14878_2, c14271);
    wire[0:0] s14879, in14879_1, in14879_2;
    wire c14879;
    assign in14879_1 = {s14275[0]};
    assign in14879_2 = {s14276[0]};
    Full_Adder FA_14879(s14879, c14879, in14879_1, in14879_2, c14274);
    wire[0:0] s14880, in14880_1, in14880_2;
    wire c14880;
    assign in14880_1 = {c14276};
    assign in14880_2 = {c14277};
    Full_Adder FA_14880(s14880, c14880, in14880_1, in14880_2, c14275);
    wire[0:0] s14881, in14881_1, in14881_2;
    wire c14881;
    assign in14881_1 = {s14279[0]};
    assign in14881_2 = {s14280[0]};
    Full_Adder FA_14881(s14881, c14881, in14881_1, in14881_2, c14278);
    wire[0:0] s14882, in14882_1, in14882_2;
    wire c14882;
    assign in14882_1 = {c14280};
    assign in14882_2 = {c14281};
    Full_Adder FA_14882(s14882, c14882, in14882_1, in14882_2, c14279);
    wire[0:0] s14883, in14883_1, in14883_2;
    wire c14883;
    assign in14883_1 = {s14283[0]};
    assign in14883_2 = {s14284[0]};
    Full_Adder FA_14883(s14883, c14883, in14883_1, in14883_2, c14282);
    wire[0:0] s14884, in14884_1, in14884_2;
    wire c14884;
    assign in14884_1 = {c14284};
    assign in14884_2 = {c14285};
    Full_Adder FA_14884(s14884, c14884, in14884_1, in14884_2, c14283);
    wire[0:0] s14885, in14885_1, in14885_2;
    wire c14885;
    assign in14885_1 = {s14287[0]};
    assign in14885_2 = {s14288[0]};
    Full_Adder FA_14885(s14885, c14885, in14885_1, in14885_2, c14286);
    wire[0:0] s14886, in14886_1, in14886_2;
    wire c14886;
    assign in14886_1 = {c14288};
    assign in14886_2 = {c14289};
    Full_Adder FA_14886(s14886, c14886, in14886_1, in14886_2, c14287);
    wire[0:0] s14887, in14887_1, in14887_2;
    wire c14887;
    assign in14887_1 = {s14291[0]};
    assign in14887_2 = {s14292[0]};
    Full_Adder FA_14887(s14887, c14887, in14887_1, in14887_2, c14290);
    wire[0:0] s14888, in14888_1, in14888_2;
    wire c14888;
    assign in14888_1 = {c14292};
    assign in14888_2 = {c14293};
    Full_Adder FA_14888(s14888, c14888, in14888_1, in14888_2, c14291);
    wire[0:0] s14889, in14889_1, in14889_2;
    wire c14889;
    assign in14889_1 = {s14295[0]};
    assign in14889_2 = {s14296[0]};
    Full_Adder FA_14889(s14889, c14889, in14889_1, in14889_2, c14294);
    wire[0:0] s14890, in14890_1, in14890_2;
    wire c14890;
    assign in14890_1 = {c14296};
    assign in14890_2 = {c14297};
    Full_Adder FA_14890(s14890, c14890, in14890_1, in14890_2, c14295);
    wire[0:0] s14891, in14891_1, in14891_2;
    wire c14891;
    assign in14891_1 = {s14299[0]};
    assign in14891_2 = {s14300[0]};
    Full_Adder FA_14891(s14891, c14891, in14891_1, in14891_2, c14298);
    wire[0:0] s14892, in14892_1, in14892_2;
    wire c14892;
    assign in14892_1 = {c14300};
    assign in14892_2 = {c14301};
    Full_Adder FA_14892(s14892, c14892, in14892_1, in14892_2, c14299);
    wire[0:0] s14893, in14893_1, in14893_2;
    wire c14893;
    assign in14893_1 = {s14303[0]};
    assign in14893_2 = {s14304[0]};
    Full_Adder FA_14893(s14893, c14893, in14893_1, in14893_2, c14302);
    wire[0:0] s14894, in14894_1, in14894_2;
    wire c14894;
    assign in14894_1 = {c14304};
    assign in14894_2 = {c14305};
    Full_Adder FA_14894(s14894, c14894, in14894_1, in14894_2, c14303);
    wire[0:0] s14895, in14895_1, in14895_2;
    wire c14895;
    assign in14895_1 = {s14307[0]};
    assign in14895_2 = {s14308[0]};
    Full_Adder FA_14895(s14895, c14895, in14895_1, in14895_2, c14306);
    wire[0:0] s14896, in14896_1, in14896_2;
    wire c14896;
    assign in14896_1 = {c14308};
    assign in14896_2 = {c14309};
    Full_Adder FA_14896(s14896, c14896, in14896_1, in14896_2, c14307);
    wire[0:0] s14897, in14897_1, in14897_2;
    wire c14897;
    assign in14897_1 = {s14311[0]};
    assign in14897_2 = {s14312[0]};
    Full_Adder FA_14897(s14897, c14897, in14897_1, in14897_2, c14310);
    wire[0:0] s14898, in14898_1, in14898_2;
    wire c14898;
    assign in14898_1 = {c14312};
    assign in14898_2 = {c14313};
    Full_Adder FA_14898(s14898, c14898, in14898_1, in14898_2, c14311);
    wire[0:0] s14899, in14899_1, in14899_2;
    wire c14899;
    assign in14899_1 = {s14315[0]};
    assign in14899_2 = {s14316[0]};
    Full_Adder FA_14899(s14899, c14899, in14899_1, in14899_2, c14314);
    wire[0:0] s14900, in14900_1, in14900_2;
    wire c14900;
    assign in14900_1 = {c14316};
    assign in14900_2 = {c14317};
    Full_Adder FA_14900(s14900, c14900, in14900_1, in14900_2, c14315);
    wire[0:0] s14901, in14901_1, in14901_2;
    wire c14901;
    assign in14901_1 = {s14319[0]};
    assign in14901_2 = {s14320[0]};
    Full_Adder FA_14901(s14901, c14901, in14901_1, in14901_2, c14318);
    wire[0:0] s14902, in14902_1, in14902_2;
    wire c14902;
    assign in14902_1 = {c14320};
    assign in14902_2 = {c14321};
    Full_Adder FA_14902(s14902, c14902, in14902_1, in14902_2, c14319);
    wire[0:0] s14903, in14903_1, in14903_2;
    wire c14903;
    assign in14903_1 = {s14323[0]};
    assign in14903_2 = {s14324[0]};
    Full_Adder FA_14903(s14903, c14903, in14903_1, in14903_2, c14322);
    wire[0:0] s14904, in14904_1, in14904_2;
    wire c14904;
    assign in14904_1 = {c14324};
    assign in14904_2 = {c14325};
    Full_Adder FA_14904(s14904, c14904, in14904_1, in14904_2, c14323);
    wire[0:0] s14905, in14905_1, in14905_2;
    wire c14905;
    assign in14905_1 = {s14327[0]};
    assign in14905_2 = {s14328[0]};
    Full_Adder FA_14905(s14905, c14905, in14905_1, in14905_2, c14326);
    wire[0:0] s14906, in14906_1, in14906_2;
    wire c14906;
    assign in14906_1 = {c14328};
    assign in14906_2 = {c14329};
    Full_Adder FA_14906(s14906, c14906, in14906_1, in14906_2, c14327);
    wire[0:0] s14907, in14907_1, in14907_2;
    wire c14907;
    assign in14907_1 = {s14331[0]};
    assign in14907_2 = {s14332[0]};
    Full_Adder FA_14907(s14907, c14907, in14907_1, in14907_2, c14330);
    wire[0:0] s14908, in14908_1, in14908_2;
    wire c14908;
    assign in14908_1 = {c14332};
    assign in14908_2 = {c14333};
    Full_Adder FA_14908(s14908, c14908, in14908_1, in14908_2, c14331);
    wire[0:0] s14909, in14909_1, in14909_2;
    wire c14909;
    assign in14909_1 = {s14335[0]};
    assign in14909_2 = {s14336[0]};
    Full_Adder FA_14909(s14909, c14909, in14909_1, in14909_2, c14334);
    wire[0:0] s14910, in14910_1, in14910_2;
    wire c14910;
    assign in14910_1 = {c14336};
    assign in14910_2 = {c14337};
    Full_Adder FA_14910(s14910, c14910, in14910_1, in14910_2, c14335);
    wire[0:0] s14911, in14911_1, in14911_2;
    wire c14911;
    assign in14911_1 = {s14339[0]};
    assign in14911_2 = {s14340[0]};
    Full_Adder FA_14911(s14911, c14911, in14911_1, in14911_2, c14338);
    wire[0:0] s14912, in14912_1, in14912_2;
    wire c14912;
    assign in14912_1 = {c14340};
    assign in14912_2 = {c14341};
    Full_Adder FA_14912(s14912, c14912, in14912_1, in14912_2, c14339);
    wire[0:0] s14913, in14913_1, in14913_2;
    wire c14913;
    assign in14913_1 = {s14343[0]};
    assign in14913_2 = {s14344[0]};
    Full_Adder FA_14913(s14913, c14913, in14913_1, in14913_2, c14342);
    wire[0:0] s14914, in14914_1, in14914_2;
    wire c14914;
    assign in14914_1 = {c14344};
    assign in14914_2 = {c14345};
    Full_Adder FA_14914(s14914, c14914, in14914_1, in14914_2, c14343);
    wire[0:0] s14915, in14915_1, in14915_2;
    wire c14915;
    assign in14915_1 = {s14347[0]};
    assign in14915_2 = {s14348[0]};
    Full_Adder FA_14915(s14915, c14915, in14915_1, in14915_2, c14346);
    wire[0:0] s14916, in14916_1, in14916_2;
    wire c14916;
    assign in14916_1 = {c14348};
    assign in14916_2 = {c14349};
    Full_Adder FA_14916(s14916, c14916, in14916_1, in14916_2, c14347);
    wire[0:0] s14917, in14917_1, in14917_2;
    wire c14917;
    assign in14917_1 = {s14351[0]};
    assign in14917_2 = {s14352[0]};
    Full_Adder FA_14917(s14917, c14917, in14917_1, in14917_2, c14350);
    wire[0:0] s14918, in14918_1, in14918_2;
    wire c14918;
    assign in14918_1 = {c14352};
    assign in14918_2 = {c14353};
    Full_Adder FA_14918(s14918, c14918, in14918_1, in14918_2, c14351);
    wire[0:0] s14919, in14919_1, in14919_2;
    wire c14919;
    assign in14919_1 = {s14355[0]};
    assign in14919_2 = {s14356[0]};
    Full_Adder FA_14919(s14919, c14919, in14919_1, in14919_2, c14354);
    wire[0:0] s14920, in14920_1, in14920_2;
    wire c14920;
    assign in14920_1 = {c14356};
    assign in14920_2 = {c14357};
    Full_Adder FA_14920(s14920, c14920, in14920_1, in14920_2, c14355);
    wire[0:0] s14921, in14921_1, in14921_2;
    wire c14921;
    assign in14921_1 = {s14359[0]};
    assign in14921_2 = {s14360[0]};
    Full_Adder FA_14921(s14921, c14921, in14921_1, in14921_2, c14358);
    wire[0:0] s14922, in14922_1, in14922_2;
    wire c14922;
    assign in14922_1 = {c14360};
    assign in14922_2 = {c14361};
    Full_Adder FA_14922(s14922, c14922, in14922_1, in14922_2, c14359);
    wire[0:0] s14923, in14923_1, in14923_2;
    wire c14923;
    assign in14923_1 = {s14363[0]};
    assign in14923_2 = {s14364[0]};
    Full_Adder FA_14923(s14923, c14923, in14923_1, in14923_2, c14362);
    wire[0:0] s14924, in14924_1, in14924_2;
    wire c14924;
    assign in14924_1 = {c14364};
    assign in14924_2 = {c14365};
    Full_Adder FA_14924(s14924, c14924, in14924_1, in14924_2, c14363);
    wire[0:0] s14925, in14925_1, in14925_2;
    wire c14925;
    assign in14925_1 = {s14367[0]};
    assign in14925_2 = {s14368[0]};
    Full_Adder FA_14925(s14925, c14925, in14925_1, in14925_2, c14366);
    wire[0:0] s14926, in14926_1, in14926_2;
    wire c14926;
    assign in14926_1 = {c14368};
    assign in14926_2 = {c14369};
    Full_Adder FA_14926(s14926, c14926, in14926_1, in14926_2, c14367);
    wire[0:0] s14927, in14927_1, in14927_2;
    wire c14927;
    assign in14927_1 = {s14371[0]};
    assign in14927_2 = {s14372[0]};
    Full_Adder FA_14927(s14927, c14927, in14927_1, in14927_2, c14370);
    wire[0:0] s14928, in14928_1, in14928_2;
    wire c14928;
    assign in14928_1 = {c14372};
    assign in14928_2 = {c14373};
    Full_Adder FA_14928(s14928, c14928, in14928_1, in14928_2, c14371);
    wire[0:0] s14929, in14929_1, in14929_2;
    wire c14929;
    assign in14929_1 = {s14375[0]};
    assign in14929_2 = {s14376[0]};
    Full_Adder FA_14929(s14929, c14929, in14929_1, in14929_2, c14374);
    wire[0:0] s14930, in14930_1, in14930_2;
    wire c14930;
    assign in14930_1 = {c14376};
    assign in14930_2 = {c14377};
    Full_Adder FA_14930(s14930, c14930, in14930_1, in14930_2, c14375);
    wire[0:0] s14931, in14931_1, in14931_2;
    wire c14931;
    assign in14931_1 = {s14379[0]};
    assign in14931_2 = {s14380[0]};
    Full_Adder FA_14931(s14931, c14931, in14931_1, in14931_2, c14378);
    wire[0:0] s14932, in14932_1, in14932_2;
    wire c14932;
    assign in14932_1 = {c14380};
    assign in14932_2 = {c14381};
    Full_Adder FA_14932(s14932, c14932, in14932_1, in14932_2, c14379);
    wire[0:0] s14933, in14933_1, in14933_2;
    wire c14933;
    assign in14933_1 = {s14383[0]};
    assign in14933_2 = {s14384[0]};
    Full_Adder FA_14933(s14933, c14933, in14933_1, in14933_2, c14382);
    wire[0:0] s14934, in14934_1, in14934_2;
    wire c14934;
    assign in14934_1 = {c14384};
    assign in14934_2 = {c14385};
    Full_Adder FA_14934(s14934, c14934, in14934_1, in14934_2, c14383);
    wire[0:0] s14935, in14935_1, in14935_2;
    wire c14935;
    assign in14935_1 = {s14387[0]};
    assign in14935_2 = {s14388[0]};
    Full_Adder FA_14935(s14935, c14935, in14935_1, in14935_2, c14386);
    wire[0:0] s14936, in14936_1, in14936_2;
    wire c14936;
    assign in14936_1 = {c14388};
    assign in14936_2 = {c14389};
    Full_Adder FA_14936(s14936, c14936, in14936_1, in14936_2, c14387);
    wire[0:0] s14937, in14937_1, in14937_2;
    wire c14937;
    assign in14937_1 = {s14391[0]};
    assign in14937_2 = {s14392[0]};
    Full_Adder FA_14937(s14937, c14937, in14937_1, in14937_2, c14390);
    wire[0:0] s14938, in14938_1, in14938_2;
    wire c14938;
    assign in14938_1 = {c14392};
    assign in14938_2 = {c14393};
    Full_Adder FA_14938(s14938, c14938, in14938_1, in14938_2, c14391);
    wire[0:0] s14939, in14939_1, in14939_2;
    wire c14939;
    assign in14939_1 = {s14395[0]};
    assign in14939_2 = {s14396[0]};
    Full_Adder FA_14939(s14939, c14939, in14939_1, in14939_2, c14394);
    wire[0:0] s14940, in14940_1, in14940_2;
    wire c14940;
    assign in14940_1 = {c14396};
    assign in14940_2 = {c14397};
    Full_Adder FA_14940(s14940, c14940, in14940_1, in14940_2, c14395);
    wire[0:0] s14941, in14941_1, in14941_2;
    wire c14941;
    assign in14941_1 = {s14399[0]};
    assign in14941_2 = {s14400[0]};
    Full_Adder FA_14941(s14941, c14941, in14941_1, in14941_2, c14398);
    wire[0:0] s14942, in14942_1, in14942_2;
    wire c14942;
    assign in14942_1 = {c14400};
    assign in14942_2 = {c14401};
    Full_Adder FA_14942(s14942, c14942, in14942_1, in14942_2, c14399);
    wire[0:0] s14943, in14943_1, in14943_2;
    wire c14943;
    assign in14943_1 = {s14403[0]};
    assign in14943_2 = {s14404[0]};
    Full_Adder FA_14943(s14943, c14943, in14943_1, in14943_2, c14402);
    wire[0:0] s14944, in14944_1, in14944_2;
    wire c14944;
    assign in14944_1 = {c14404};
    assign in14944_2 = {c14405};
    Full_Adder FA_14944(s14944, c14944, in14944_1, in14944_2, c14403);
    wire[0:0] s14945, in14945_1, in14945_2;
    wire c14945;
    assign in14945_1 = {s14407[0]};
    assign in14945_2 = {s14408[0]};
    Full_Adder FA_14945(s14945, c14945, in14945_1, in14945_2, c14406);
    wire[0:0] s14946, in14946_1, in14946_2;
    wire c14946;
    assign in14946_1 = {c14408};
    assign in14946_2 = {c14409};
    Full_Adder FA_14946(s14946, c14946, in14946_1, in14946_2, c14407);
    wire[0:0] s14947, in14947_1, in14947_2;
    wire c14947;
    assign in14947_1 = {s14411[0]};
    assign in14947_2 = {s14412[0]};
    Full_Adder FA_14947(s14947, c14947, in14947_1, in14947_2, c14410);
    wire[0:0] s14948, in14948_1, in14948_2;
    wire c14948;
    assign in14948_1 = {c14412};
    assign in14948_2 = {c14413};
    Full_Adder FA_14948(s14948, c14948, in14948_1, in14948_2, c14411);
    wire[0:0] s14949, in14949_1, in14949_2;
    wire c14949;
    assign in14949_1 = {s14415[0]};
    assign in14949_2 = {s14416[0]};
    Full_Adder FA_14949(s14949, c14949, in14949_1, in14949_2, c14414);
    wire[0:0] s14950, in14950_1, in14950_2;
    wire c14950;
    assign in14950_1 = {c14416};
    assign in14950_2 = {c14417};
    Full_Adder FA_14950(s14950, c14950, in14950_1, in14950_2, c14415);
    wire[0:0] s14951, in14951_1, in14951_2;
    wire c14951;
    assign in14951_1 = {s14419[0]};
    assign in14951_2 = {s14420[0]};
    Full_Adder FA_14951(s14951, c14951, in14951_1, in14951_2, c14418);
    wire[0:0] s14952, in14952_1, in14952_2;
    wire c14952;
    assign in14952_1 = {c14420};
    assign in14952_2 = {c14421};
    Full_Adder FA_14952(s14952, c14952, in14952_1, in14952_2, c14419);
    wire[0:0] s14953, in14953_1, in14953_2;
    wire c14953;
    assign in14953_1 = {s14423[0]};
    assign in14953_2 = {s14424[0]};
    Full_Adder FA_14953(s14953, c14953, in14953_1, in14953_2, c14422);
    wire[0:0] s14954, in14954_1, in14954_2;
    wire c14954;
    assign in14954_1 = {c14424};
    assign in14954_2 = {c14425};
    Full_Adder FA_14954(s14954, c14954, in14954_1, in14954_2, c14423);
    wire[0:0] s14955, in14955_1, in14955_2;
    wire c14955;
    assign in14955_1 = {s14427[0]};
    assign in14955_2 = {s14428[0]};
    Full_Adder FA_14955(s14955, c14955, in14955_1, in14955_2, c14426);
    wire[0:0] s14956, in14956_1, in14956_2;
    wire c14956;
    assign in14956_1 = {c14428};
    assign in14956_2 = {c14429};
    Full_Adder FA_14956(s14956, c14956, in14956_1, in14956_2, c14427);
    wire[0:0] s14957, in14957_1, in14957_2;
    wire c14957;
    assign in14957_1 = {s14431[0]};
    assign in14957_2 = {s14432[0]};
    Full_Adder FA_14957(s14957, c14957, in14957_1, in14957_2, c14430);
    wire[0:0] s14958, in14958_1, in14958_2;
    wire c14958;
    assign in14958_1 = {c14432};
    assign in14958_2 = {c14433};
    Full_Adder FA_14958(s14958, c14958, in14958_1, in14958_2, c14431);
    wire[0:0] s14959, in14959_1, in14959_2;
    wire c14959;
    assign in14959_1 = {s14435[0]};
    assign in14959_2 = {s14436[0]};
    Full_Adder FA_14959(s14959, c14959, in14959_1, in14959_2, c14434);
    wire[0:0] s14960, in14960_1, in14960_2;
    wire c14960;
    assign in14960_1 = {c14436};
    assign in14960_2 = {c14437};
    Full_Adder FA_14960(s14960, c14960, in14960_1, in14960_2, c14435);
    wire[0:0] s14961, in14961_1, in14961_2;
    wire c14961;
    assign in14961_1 = {s14439[0]};
    assign in14961_2 = {s14440[0]};
    Full_Adder FA_14961(s14961, c14961, in14961_1, in14961_2, c14438);
    wire[0:0] s14962, in14962_1, in14962_2;
    wire c14962;
    assign in14962_1 = {c14440};
    assign in14962_2 = {c14441};
    Full_Adder FA_14962(s14962, c14962, in14962_1, in14962_2, c14439);
    wire[0:0] s14963, in14963_1, in14963_2;
    wire c14963;
    assign in14963_1 = {s14443[0]};
    assign in14963_2 = {s14444[0]};
    Full_Adder FA_14963(s14963, c14963, in14963_1, in14963_2, c14442);
    wire[0:0] s14964, in14964_1, in14964_2;
    wire c14964;
    assign in14964_1 = {c14444};
    assign in14964_2 = {c14445};
    Full_Adder FA_14964(s14964, c14964, in14964_1, in14964_2, c14443);
    wire[0:0] s14965, in14965_1, in14965_2;
    wire c14965;
    assign in14965_1 = {s14447[0]};
    assign in14965_2 = {s14448[0]};
    Full_Adder FA_14965(s14965, c14965, in14965_1, in14965_2, c14446);
    wire[0:0] s14966, in14966_1, in14966_2;
    wire c14966;
    assign in14966_1 = {c14448};
    assign in14966_2 = {c14449};
    Full_Adder FA_14966(s14966, c14966, in14966_1, in14966_2, c14447);
    wire[0:0] s14967, in14967_1, in14967_2;
    wire c14967;
    assign in14967_1 = {s14451[0]};
    assign in14967_2 = {s14452[0]};
    Full_Adder FA_14967(s14967, c14967, in14967_1, in14967_2, c14450);
    wire[0:0] s14968, in14968_1, in14968_2;
    wire c14968;
    assign in14968_1 = {c14452};
    assign in14968_2 = {c14453};
    Full_Adder FA_14968(s14968, c14968, in14968_1, in14968_2, c14451);
    wire[0:0] s14969, in14969_1, in14969_2;
    wire c14969;
    assign in14969_1 = {s14455[0]};
    assign in14969_2 = {s14456[0]};
    Full_Adder FA_14969(s14969, c14969, in14969_1, in14969_2, c14454);
    wire[0:0] s14970, in14970_1, in14970_2;
    wire c14970;
    assign in14970_1 = {c14456};
    assign in14970_2 = {c14457};
    Full_Adder FA_14970(s14970, c14970, in14970_1, in14970_2, c14455);
    wire[0:0] s14971, in14971_1, in14971_2;
    wire c14971;
    assign in14971_1 = {s14459[0]};
    assign in14971_2 = {s14460[0]};
    Full_Adder FA_14971(s14971, c14971, in14971_1, in14971_2, c14458);
    wire[0:0] s14972, in14972_1, in14972_2;
    wire c14972;
    assign in14972_1 = {c14460};
    assign in14972_2 = {c14461};
    Full_Adder FA_14972(s14972, c14972, in14972_1, in14972_2, c14459);
    wire[0:0] s14973, in14973_1, in14973_2;
    wire c14973;
    assign in14973_1 = {s14463[0]};
    assign in14973_2 = {s14464[0]};
    Full_Adder FA_14973(s14973, c14973, in14973_1, in14973_2, c14462);
    wire[0:0] s14974, in14974_1, in14974_2;
    wire c14974;
    assign in14974_1 = {c14464};
    assign in14974_2 = {c14465};
    Full_Adder FA_14974(s14974, c14974, in14974_1, in14974_2, c14463);
    wire[0:0] s14975, in14975_1, in14975_2;
    wire c14975;
    assign in14975_1 = {s14467[0]};
    assign in14975_2 = {s14468[0]};
    Full_Adder FA_14975(s14975, c14975, in14975_1, in14975_2, c14466);
    wire[0:0] s14976, in14976_1, in14976_2;
    wire c14976;
    assign in14976_1 = {c14468};
    assign in14976_2 = {c14469};
    Full_Adder FA_14976(s14976, c14976, in14976_1, in14976_2, c14467);
    wire[0:0] s14977, in14977_1, in14977_2;
    wire c14977;
    assign in14977_1 = {s14471[0]};
    assign in14977_2 = {s14472[0]};
    Full_Adder FA_14977(s14977, c14977, in14977_1, in14977_2, c14470);
    wire[0:0] s14978, in14978_1, in14978_2;
    wire c14978;
    assign in14978_1 = {c14472};
    assign in14978_2 = {c14473};
    Full_Adder FA_14978(s14978, c14978, in14978_1, in14978_2, c14471);
    wire[0:0] s14979, in14979_1, in14979_2;
    wire c14979;
    assign in14979_1 = {s14475[0]};
    assign in14979_2 = {s14476[0]};
    Full_Adder FA_14979(s14979, c14979, in14979_1, in14979_2, c14474);
    wire[0:0] s14980, in14980_1, in14980_2;
    wire c14980;
    assign in14980_1 = {c14476};
    assign in14980_2 = {c14477};
    Full_Adder FA_14980(s14980, c14980, in14980_1, in14980_2, c14475);
    wire[0:0] s14981, in14981_1, in14981_2;
    wire c14981;
    assign in14981_1 = {s14479[0]};
    assign in14981_2 = {s14480[0]};
    Full_Adder FA_14981(s14981, c14981, in14981_1, in14981_2, c14478);
    wire[0:0] s14982, in14982_1, in14982_2;
    wire c14982;
    assign in14982_1 = {c14480};
    assign in14982_2 = {c14481};
    Full_Adder FA_14982(s14982, c14982, in14982_1, in14982_2, c14479);
    wire[0:0] s14983, in14983_1, in14983_2;
    wire c14983;
    assign in14983_1 = {s14483[0]};
    assign in14983_2 = {s14484[0]};
    Full_Adder FA_14983(s14983, c14983, in14983_1, in14983_2, c14482);
    wire[0:0] s14984, in14984_1, in14984_2;
    wire c14984;
    assign in14984_1 = {c14484};
    assign in14984_2 = {c14485};
    Full_Adder FA_14984(s14984, c14984, in14984_1, in14984_2, c14483);
    wire[0:0] s14985, in14985_1, in14985_2;
    wire c14985;
    assign in14985_1 = {s14487[0]};
    assign in14985_2 = {s14488[0]};
    Full_Adder FA_14985(s14985, c14985, in14985_1, in14985_2, c14486);
    wire[0:0] s14986, in14986_1, in14986_2;
    wire c14986;
    assign in14986_1 = {c14488};
    assign in14986_2 = {c14489};
    Full_Adder FA_14986(s14986, c14986, in14986_1, in14986_2, c14487);
    wire[0:0] s14987, in14987_1, in14987_2;
    wire c14987;
    assign in14987_1 = {s14491[0]};
    assign in14987_2 = {s14492[0]};
    Full_Adder FA_14987(s14987, c14987, in14987_1, in14987_2, c14490);
    wire[0:0] s14988, in14988_1, in14988_2;
    wire c14988;
    assign in14988_1 = {c14492};
    assign in14988_2 = {c14493};
    Full_Adder FA_14988(s14988, c14988, in14988_1, in14988_2, c14491);
    wire[0:0] s14989, in14989_1, in14989_2;
    wire c14989;
    assign in14989_1 = {s14495[0]};
    assign in14989_2 = {s14496[0]};
    Full_Adder FA_14989(s14989, c14989, in14989_1, in14989_2, c14494);
    wire[0:0] s14990, in14990_1, in14990_2;
    wire c14990;
    assign in14990_1 = {c14496};
    assign in14990_2 = {c14497};
    Full_Adder FA_14990(s14990, c14990, in14990_1, in14990_2, c14495);
    wire[0:0] s14991, in14991_1, in14991_2;
    wire c14991;
    assign in14991_1 = {s14499[0]};
    assign in14991_2 = {s14500[0]};
    Full_Adder FA_14991(s14991, c14991, in14991_1, in14991_2, c14498);
    wire[0:0] s14992, in14992_1, in14992_2;
    wire c14992;
    assign in14992_1 = {c14500};
    assign in14992_2 = {c14501};
    Full_Adder FA_14992(s14992, c14992, in14992_1, in14992_2, c14499);
    wire[0:0] s14993, in14993_1, in14993_2;
    wire c14993;
    assign in14993_1 = {s14503[0]};
    assign in14993_2 = {s14504[0]};
    Full_Adder FA_14993(s14993, c14993, in14993_1, in14993_2, c14502);
    wire[0:0] s14994, in14994_1, in14994_2;
    wire c14994;
    assign in14994_1 = {c14504};
    assign in14994_2 = {c14505};
    Full_Adder FA_14994(s14994, c14994, in14994_1, in14994_2, c14503);
    wire[0:0] s14995, in14995_1, in14995_2;
    wire c14995;
    assign in14995_1 = {s14507[0]};
    assign in14995_2 = {s14508[0]};
    Full_Adder FA_14995(s14995, c14995, in14995_1, in14995_2, c14506);
    wire[0:0] s14996, in14996_1, in14996_2;
    wire c14996;
    assign in14996_1 = {c14508};
    assign in14996_2 = {c14509};
    Full_Adder FA_14996(s14996, c14996, in14996_1, in14996_2, c14507);
    wire[0:0] s14997, in14997_1, in14997_2;
    wire c14997;
    assign in14997_1 = {s14511[0]};
    assign in14997_2 = {s14512[0]};
    Full_Adder FA_14997(s14997, c14997, in14997_1, in14997_2, c14510);
    wire[0:0] s14998, in14998_1, in14998_2;
    wire c14998;
    assign in14998_1 = {c14511};
    assign in14998_2 = {c14512};
    Full_Adder FA_14998(s14998, c14998, in14998_1, in14998_2, pp127[118]);
    wire[0:0] s14999, in14999_1, in14999_2;
    wire c14999;
    assign in14999_1 = {c14514};
    assign in14999_2 = {s14515[0]};
    Full_Adder FA_14999(s14999, c14999, in14999_1, in14999_2, c14513);
    wire[0:0] s15000, in15000_1, in15000_2;
    wire c15000;
    assign in15000_1 = {pp126[120]};
    assign in15000_2 = {pp127[119]};
    Full_Adder FA_15000(s15000, c15000, in15000_1, in15000_2, pp125[121]);
    wire[0:0] s15001, in15001_1, in15001_2;
    wire c15001;
    assign in15001_1 = {c14516};
    assign in15001_2 = {c14517};
    Full_Adder FA_15001(s15001, c15001, in15001_1, in15001_2, c14515);
    wire[0:0] s15002, in15002_1, in15002_2;
    wire c15002;
    assign in15002_1 = {pp124[123]};
    assign in15002_2 = {pp125[122]};
    Full_Adder FA_15002(s15002, c15002, in15002_1, in15002_2, pp123[124]);
    wire[0:0] s15003, in15003_1, in15003_2;
    wire c15003;
    assign in15003_1 = {pp127[120]};
    assign in15003_2 = {c14518};
    Full_Adder FA_15003(s15003, c15003, in15003_1, in15003_2, pp126[121]);
    wire[0:0] s15004, in15004_1, in15004_2;
    wire c15004;
    assign in15004_1 = {pp122[126]};
    assign in15004_2 = {pp123[125]};
    Full_Adder FA_15004(s15004, c15004, in15004_1, in15004_2, pp121[127]);
    wire[0:0] s15005, in15005_1, in15005_2;
    wire c15005;
    assign in15005_1 = {pp125[123]};
    assign in15005_2 = {pp126[122]};
    Full_Adder FA_15005(s15005, c15005, in15005_1, in15005_2, pp124[124]);
    wire[0:0] s15006, in15006_1, in15006_2;
    wire c15006;
    assign in15006_1 = {pp123[126]};
    assign in15006_2 = {pp124[125]};
    Full_Adder FA_15006(s15006, c15006, in15006_1, in15006_2, pp122[127]);

    /*Stage 9*/
    wire[0:0] s15007, in15007_1, in15007_2;
    wire c15007;
    assign in15007_1 = {pp0[4]};
    assign in15007_2 = {pp1[3]};
    Half_Adder HA_15007(s15007, c15007, in15007_1, in15007_2);
    wire[0:0] s15008, in15008_1, in15008_2;
    wire c15008;
    assign in15008_1 = {pp1[4]};
    assign in15008_2 = {pp2[3]};
    Full_Adder FA_15008(s15008, c15008, in15008_1, in15008_2, pp0[5]);
    wire[0:0] s15009, in15009_1, in15009_2;
    wire c15009;
    assign in15009_1 = {pp3[2]};
    assign in15009_2 = {pp4[1]};
    Half_Adder HA_15009(s15009, c15009, in15009_1, in15009_2);
    wire[0:0] s15010, in15010_1, in15010_2;
    wire c15010;
    assign in15010_1 = {pp3[3]};
    assign in15010_2 = {pp4[2]};
    Full_Adder FA_15010(s15010, c15010, in15010_1, in15010_2, pp2[4]);
    wire[0:0] s15011, in15011_1, in15011_2;
    wire c15011;
    assign in15011_1 = {pp6[0]};
    assign in15011_2 = {s14521[0]};
    Full_Adder FA_15011(s15011, c15011, in15011_1, in15011_2, pp5[1]);
    wire[0:0] s15012, in15012_1, in15012_2;
    wire c15012;
    assign in15012_1 = {pp6[1]};
    assign in15012_2 = {pp7[0]};
    Full_Adder FA_15012(s15012, c15012, in15012_1, in15012_2, pp5[2]);
    wire[0:0] s15013, in15013_1, in15013_2;
    wire c15013;
    assign in15013_1 = {s14522[0]};
    assign in15013_2 = {s14523[0]};
    Full_Adder FA_15013(s15013, c15013, in15013_1, in15013_2, c14521);
    wire[0:0] s15014, in15014_1, in15014_2;
    wire c15014;
    assign in15014_1 = {s13573[0]};
    assign in15014_2 = {c14522};
    Full_Adder FA_15014(s15014, c15014, in15014_1, in15014_2, pp8[0]);
    wire[0:0] s15015, in15015_1, in15015_2;
    wire c15015;
    assign in15015_1 = {s14524[0]};
    assign in15015_2 = {s14525[0]};
    Full_Adder FA_15015(s15015, c15015, in15015_1, in15015_2, c14523);
    wire[0:0] s15016, in15016_1, in15016_2;
    wire c15016;
    assign in15016_1 = {s13575[0]};
    assign in15016_2 = {c14524};
    Full_Adder FA_15016(s15016, c15016, in15016_1, in15016_2, s13574[0]);
    wire[0:0] s15017, in15017_1, in15017_2;
    wire c15017;
    assign in15017_1 = {s14526[0]};
    assign in15017_2 = {s14527[0]};
    Full_Adder FA_15017(s15017, c15017, in15017_1, in15017_2, c14525);
    wire[0:0] s15018, in15018_1, in15018_2;
    wire c15018;
    assign in15018_1 = {s13578[0]};
    assign in15018_2 = {c14526};
    Full_Adder FA_15018(s15018, c15018, in15018_1, in15018_2, s13577[0]);
    wire[0:0] s15019, in15019_1, in15019_2;
    wire c15019;
    assign in15019_1 = {s14528[0]};
    assign in15019_2 = {s14529[0]};
    Full_Adder FA_15019(s15019, c15019, in15019_1, in15019_2, c14527);
    wire[0:0] s15020, in15020_1, in15020_2;
    wire c15020;
    assign in15020_1 = {s13582[0]};
    assign in15020_2 = {c14528};
    Full_Adder FA_15020(s15020, c15020, in15020_1, in15020_2, s13581[0]);
    wire[0:0] s15021, in15021_1, in15021_2;
    wire c15021;
    assign in15021_1 = {s14530[0]};
    assign in15021_2 = {s14531[0]};
    Full_Adder FA_15021(s15021, c15021, in15021_1, in15021_2, c14529);
    wire[0:0] s15022, in15022_1, in15022_2;
    wire c15022;
    assign in15022_1 = {s13586[0]};
    assign in15022_2 = {c14530};
    Full_Adder FA_15022(s15022, c15022, in15022_1, in15022_2, s13585[0]);
    wire[0:0] s15023, in15023_1, in15023_2;
    wire c15023;
    assign in15023_1 = {s14532[0]};
    assign in15023_2 = {s14533[0]};
    Full_Adder FA_15023(s15023, c15023, in15023_1, in15023_2, c14531);
    wire[0:0] s15024, in15024_1, in15024_2;
    wire c15024;
    assign in15024_1 = {s13590[0]};
    assign in15024_2 = {c14532};
    Full_Adder FA_15024(s15024, c15024, in15024_1, in15024_2, s13589[0]);
    wire[0:0] s15025, in15025_1, in15025_2;
    wire c15025;
    assign in15025_1 = {s14534[0]};
    assign in15025_2 = {s14535[0]};
    Full_Adder FA_15025(s15025, c15025, in15025_1, in15025_2, c14533);
    wire[0:0] s15026, in15026_1, in15026_2;
    wire c15026;
    assign in15026_1 = {s13594[0]};
    assign in15026_2 = {c14534};
    Full_Adder FA_15026(s15026, c15026, in15026_1, in15026_2, s13593[0]);
    wire[0:0] s15027, in15027_1, in15027_2;
    wire c15027;
    assign in15027_1 = {s14536[0]};
    assign in15027_2 = {s14537[0]};
    Full_Adder FA_15027(s15027, c15027, in15027_1, in15027_2, c14535);
    wire[0:0] s15028, in15028_1, in15028_2;
    wire c15028;
    assign in15028_1 = {s13598[0]};
    assign in15028_2 = {c14536};
    Full_Adder FA_15028(s15028, c15028, in15028_1, in15028_2, s13597[0]);
    wire[0:0] s15029, in15029_1, in15029_2;
    wire c15029;
    assign in15029_1 = {s14538[0]};
    assign in15029_2 = {s14539[0]};
    Full_Adder FA_15029(s15029, c15029, in15029_1, in15029_2, c14537);
    wire[0:0] s15030, in15030_1, in15030_2;
    wire c15030;
    assign in15030_1 = {s13602[0]};
    assign in15030_2 = {c14538};
    Full_Adder FA_15030(s15030, c15030, in15030_1, in15030_2, s13601[0]);
    wire[0:0] s15031, in15031_1, in15031_2;
    wire c15031;
    assign in15031_1 = {s14540[0]};
    assign in15031_2 = {s14541[0]};
    Full_Adder FA_15031(s15031, c15031, in15031_1, in15031_2, c14539);
    wire[0:0] s15032, in15032_1, in15032_2;
    wire c15032;
    assign in15032_1 = {s13606[0]};
    assign in15032_2 = {c14540};
    Full_Adder FA_15032(s15032, c15032, in15032_1, in15032_2, s13605[0]);
    wire[0:0] s15033, in15033_1, in15033_2;
    wire c15033;
    assign in15033_1 = {s14542[0]};
    assign in15033_2 = {s14543[0]};
    Full_Adder FA_15033(s15033, c15033, in15033_1, in15033_2, c14541);
    wire[0:0] s15034, in15034_1, in15034_2;
    wire c15034;
    assign in15034_1 = {s13610[0]};
    assign in15034_2 = {c14542};
    Full_Adder FA_15034(s15034, c15034, in15034_1, in15034_2, s13609[0]);
    wire[0:0] s15035, in15035_1, in15035_2;
    wire c15035;
    assign in15035_1 = {s14544[0]};
    assign in15035_2 = {s14545[0]};
    Full_Adder FA_15035(s15035, c15035, in15035_1, in15035_2, c14543);
    wire[0:0] s15036, in15036_1, in15036_2;
    wire c15036;
    assign in15036_1 = {s13614[0]};
    assign in15036_2 = {c14544};
    Full_Adder FA_15036(s15036, c15036, in15036_1, in15036_2, s13613[0]);
    wire[0:0] s15037, in15037_1, in15037_2;
    wire c15037;
    assign in15037_1 = {s14546[0]};
    assign in15037_2 = {s14547[0]};
    Full_Adder FA_15037(s15037, c15037, in15037_1, in15037_2, c14545);
    wire[0:0] s15038, in15038_1, in15038_2;
    wire c15038;
    assign in15038_1 = {s13618[0]};
    assign in15038_2 = {c14546};
    Full_Adder FA_15038(s15038, c15038, in15038_1, in15038_2, s13617[0]);
    wire[0:0] s15039, in15039_1, in15039_2;
    wire c15039;
    assign in15039_1 = {s14548[0]};
    assign in15039_2 = {s14549[0]};
    Full_Adder FA_15039(s15039, c15039, in15039_1, in15039_2, c14547);
    wire[0:0] s15040, in15040_1, in15040_2;
    wire c15040;
    assign in15040_1 = {s13622[0]};
    assign in15040_2 = {c14548};
    Full_Adder FA_15040(s15040, c15040, in15040_1, in15040_2, s13621[0]);
    wire[0:0] s15041, in15041_1, in15041_2;
    wire c15041;
    assign in15041_1 = {s14550[0]};
    assign in15041_2 = {s14551[0]};
    Full_Adder FA_15041(s15041, c15041, in15041_1, in15041_2, c14549);
    wire[0:0] s15042, in15042_1, in15042_2;
    wire c15042;
    assign in15042_1 = {s13626[0]};
    assign in15042_2 = {c14550};
    Full_Adder FA_15042(s15042, c15042, in15042_1, in15042_2, s13625[0]);
    wire[0:0] s15043, in15043_1, in15043_2;
    wire c15043;
    assign in15043_1 = {s14552[0]};
    assign in15043_2 = {s14553[0]};
    Full_Adder FA_15043(s15043, c15043, in15043_1, in15043_2, c14551);
    wire[0:0] s15044, in15044_1, in15044_2;
    wire c15044;
    assign in15044_1 = {s13630[0]};
    assign in15044_2 = {c14552};
    Full_Adder FA_15044(s15044, c15044, in15044_1, in15044_2, s13629[0]);
    wire[0:0] s15045, in15045_1, in15045_2;
    wire c15045;
    assign in15045_1 = {s14554[0]};
    assign in15045_2 = {s14555[0]};
    Full_Adder FA_15045(s15045, c15045, in15045_1, in15045_2, c14553);
    wire[0:0] s15046, in15046_1, in15046_2;
    wire c15046;
    assign in15046_1 = {s13634[0]};
    assign in15046_2 = {c14554};
    Full_Adder FA_15046(s15046, c15046, in15046_1, in15046_2, s13633[0]);
    wire[0:0] s15047, in15047_1, in15047_2;
    wire c15047;
    assign in15047_1 = {s14556[0]};
    assign in15047_2 = {s14557[0]};
    Full_Adder FA_15047(s15047, c15047, in15047_1, in15047_2, c14555);
    wire[0:0] s15048, in15048_1, in15048_2;
    wire c15048;
    assign in15048_1 = {s13638[0]};
    assign in15048_2 = {c14556};
    Full_Adder FA_15048(s15048, c15048, in15048_1, in15048_2, s13637[0]);
    wire[0:0] s15049, in15049_1, in15049_2;
    wire c15049;
    assign in15049_1 = {s14558[0]};
    assign in15049_2 = {s14559[0]};
    Full_Adder FA_15049(s15049, c15049, in15049_1, in15049_2, c14557);
    wire[0:0] s15050, in15050_1, in15050_2;
    wire c15050;
    assign in15050_1 = {s13642[0]};
    assign in15050_2 = {c14558};
    Full_Adder FA_15050(s15050, c15050, in15050_1, in15050_2, s13641[0]);
    wire[0:0] s15051, in15051_1, in15051_2;
    wire c15051;
    assign in15051_1 = {s14560[0]};
    assign in15051_2 = {s14561[0]};
    Full_Adder FA_15051(s15051, c15051, in15051_1, in15051_2, c14559);
    wire[0:0] s15052, in15052_1, in15052_2;
    wire c15052;
    assign in15052_1 = {s13646[0]};
    assign in15052_2 = {c14560};
    Full_Adder FA_15052(s15052, c15052, in15052_1, in15052_2, s13645[0]);
    wire[0:0] s15053, in15053_1, in15053_2;
    wire c15053;
    assign in15053_1 = {s14562[0]};
    assign in15053_2 = {s14563[0]};
    Full_Adder FA_15053(s15053, c15053, in15053_1, in15053_2, c14561);
    wire[0:0] s15054, in15054_1, in15054_2;
    wire c15054;
    assign in15054_1 = {s13650[0]};
    assign in15054_2 = {c14562};
    Full_Adder FA_15054(s15054, c15054, in15054_1, in15054_2, s13649[0]);
    wire[0:0] s15055, in15055_1, in15055_2;
    wire c15055;
    assign in15055_1 = {s14564[0]};
    assign in15055_2 = {s14565[0]};
    Full_Adder FA_15055(s15055, c15055, in15055_1, in15055_2, c14563);
    wire[0:0] s15056, in15056_1, in15056_2;
    wire c15056;
    assign in15056_1 = {s13654[0]};
    assign in15056_2 = {c14564};
    Full_Adder FA_15056(s15056, c15056, in15056_1, in15056_2, s13653[0]);
    wire[0:0] s15057, in15057_1, in15057_2;
    wire c15057;
    assign in15057_1 = {s14566[0]};
    assign in15057_2 = {s14567[0]};
    Full_Adder FA_15057(s15057, c15057, in15057_1, in15057_2, c14565);
    wire[0:0] s15058, in15058_1, in15058_2;
    wire c15058;
    assign in15058_1 = {s13658[0]};
    assign in15058_2 = {c14566};
    Full_Adder FA_15058(s15058, c15058, in15058_1, in15058_2, s13657[0]);
    wire[0:0] s15059, in15059_1, in15059_2;
    wire c15059;
    assign in15059_1 = {s14568[0]};
    assign in15059_2 = {s14569[0]};
    Full_Adder FA_15059(s15059, c15059, in15059_1, in15059_2, c14567);
    wire[0:0] s15060, in15060_1, in15060_2;
    wire c15060;
    assign in15060_1 = {s13662[0]};
    assign in15060_2 = {c14568};
    Full_Adder FA_15060(s15060, c15060, in15060_1, in15060_2, s13661[0]);
    wire[0:0] s15061, in15061_1, in15061_2;
    wire c15061;
    assign in15061_1 = {s14570[0]};
    assign in15061_2 = {s14571[0]};
    Full_Adder FA_15061(s15061, c15061, in15061_1, in15061_2, c14569);
    wire[0:0] s15062, in15062_1, in15062_2;
    wire c15062;
    assign in15062_1 = {s13666[0]};
    assign in15062_2 = {c14570};
    Full_Adder FA_15062(s15062, c15062, in15062_1, in15062_2, s13665[0]);
    wire[0:0] s15063, in15063_1, in15063_2;
    wire c15063;
    assign in15063_1 = {s14572[0]};
    assign in15063_2 = {s14573[0]};
    Full_Adder FA_15063(s15063, c15063, in15063_1, in15063_2, c14571);
    wire[0:0] s15064, in15064_1, in15064_2;
    wire c15064;
    assign in15064_1 = {s13670[0]};
    assign in15064_2 = {c14572};
    Full_Adder FA_15064(s15064, c15064, in15064_1, in15064_2, s13669[0]);
    wire[0:0] s15065, in15065_1, in15065_2;
    wire c15065;
    assign in15065_1 = {s14574[0]};
    assign in15065_2 = {s14575[0]};
    Full_Adder FA_15065(s15065, c15065, in15065_1, in15065_2, c14573);
    wire[0:0] s15066, in15066_1, in15066_2;
    wire c15066;
    assign in15066_1 = {s13674[0]};
    assign in15066_2 = {c14574};
    Full_Adder FA_15066(s15066, c15066, in15066_1, in15066_2, s13673[0]);
    wire[0:0] s15067, in15067_1, in15067_2;
    wire c15067;
    assign in15067_1 = {s14576[0]};
    assign in15067_2 = {s14577[0]};
    Full_Adder FA_15067(s15067, c15067, in15067_1, in15067_2, c14575);
    wire[0:0] s15068, in15068_1, in15068_2;
    wire c15068;
    assign in15068_1 = {s13678[0]};
    assign in15068_2 = {c14576};
    Full_Adder FA_15068(s15068, c15068, in15068_1, in15068_2, s13677[0]);
    wire[0:0] s15069, in15069_1, in15069_2;
    wire c15069;
    assign in15069_1 = {s14578[0]};
    assign in15069_2 = {s14579[0]};
    Full_Adder FA_15069(s15069, c15069, in15069_1, in15069_2, c14577);
    wire[0:0] s15070, in15070_1, in15070_2;
    wire c15070;
    assign in15070_1 = {s13682[0]};
    assign in15070_2 = {c14578};
    Full_Adder FA_15070(s15070, c15070, in15070_1, in15070_2, s13681[0]);
    wire[0:0] s15071, in15071_1, in15071_2;
    wire c15071;
    assign in15071_1 = {s14580[0]};
    assign in15071_2 = {s14581[0]};
    Full_Adder FA_15071(s15071, c15071, in15071_1, in15071_2, c14579);
    wire[0:0] s15072, in15072_1, in15072_2;
    wire c15072;
    assign in15072_1 = {s13686[0]};
    assign in15072_2 = {c14580};
    Full_Adder FA_15072(s15072, c15072, in15072_1, in15072_2, s13685[0]);
    wire[0:0] s15073, in15073_1, in15073_2;
    wire c15073;
    assign in15073_1 = {s14582[0]};
    assign in15073_2 = {s14583[0]};
    Full_Adder FA_15073(s15073, c15073, in15073_1, in15073_2, c14581);
    wire[0:0] s15074, in15074_1, in15074_2;
    wire c15074;
    assign in15074_1 = {s13690[0]};
    assign in15074_2 = {c14582};
    Full_Adder FA_15074(s15074, c15074, in15074_1, in15074_2, s13689[0]);
    wire[0:0] s15075, in15075_1, in15075_2;
    wire c15075;
    assign in15075_1 = {s14584[0]};
    assign in15075_2 = {s14585[0]};
    Full_Adder FA_15075(s15075, c15075, in15075_1, in15075_2, c14583);
    wire[0:0] s15076, in15076_1, in15076_2;
    wire c15076;
    assign in15076_1 = {s13694[0]};
    assign in15076_2 = {c14584};
    Full_Adder FA_15076(s15076, c15076, in15076_1, in15076_2, s13693[0]);
    wire[0:0] s15077, in15077_1, in15077_2;
    wire c15077;
    assign in15077_1 = {s14586[0]};
    assign in15077_2 = {s14587[0]};
    Full_Adder FA_15077(s15077, c15077, in15077_1, in15077_2, c14585);
    wire[0:0] s15078, in15078_1, in15078_2;
    wire c15078;
    assign in15078_1 = {s13698[0]};
    assign in15078_2 = {c14586};
    Full_Adder FA_15078(s15078, c15078, in15078_1, in15078_2, s13697[0]);
    wire[0:0] s15079, in15079_1, in15079_2;
    wire c15079;
    assign in15079_1 = {s14588[0]};
    assign in15079_2 = {s14589[0]};
    Full_Adder FA_15079(s15079, c15079, in15079_1, in15079_2, c14587);
    wire[0:0] s15080, in15080_1, in15080_2;
    wire c15080;
    assign in15080_1 = {s13702[0]};
    assign in15080_2 = {c14588};
    Full_Adder FA_15080(s15080, c15080, in15080_1, in15080_2, s13701[0]);
    wire[0:0] s15081, in15081_1, in15081_2;
    wire c15081;
    assign in15081_1 = {s14590[0]};
    assign in15081_2 = {s14591[0]};
    Full_Adder FA_15081(s15081, c15081, in15081_1, in15081_2, c14589);
    wire[0:0] s15082, in15082_1, in15082_2;
    wire c15082;
    assign in15082_1 = {s13706[0]};
    assign in15082_2 = {c14590};
    Full_Adder FA_15082(s15082, c15082, in15082_1, in15082_2, s13705[0]);
    wire[0:0] s15083, in15083_1, in15083_2;
    wire c15083;
    assign in15083_1 = {s14592[0]};
    assign in15083_2 = {s14593[0]};
    Full_Adder FA_15083(s15083, c15083, in15083_1, in15083_2, c14591);
    wire[0:0] s15084, in15084_1, in15084_2;
    wire c15084;
    assign in15084_1 = {s13710[0]};
    assign in15084_2 = {c14592};
    Full_Adder FA_15084(s15084, c15084, in15084_1, in15084_2, s13709[0]);
    wire[0:0] s15085, in15085_1, in15085_2;
    wire c15085;
    assign in15085_1 = {s14594[0]};
    assign in15085_2 = {s14595[0]};
    Full_Adder FA_15085(s15085, c15085, in15085_1, in15085_2, c14593);
    wire[0:0] s15086, in15086_1, in15086_2;
    wire c15086;
    assign in15086_1 = {s13714[0]};
    assign in15086_2 = {c14594};
    Full_Adder FA_15086(s15086, c15086, in15086_1, in15086_2, s13713[0]);
    wire[0:0] s15087, in15087_1, in15087_2;
    wire c15087;
    assign in15087_1 = {s14596[0]};
    assign in15087_2 = {s14597[0]};
    Full_Adder FA_15087(s15087, c15087, in15087_1, in15087_2, c14595);
    wire[0:0] s15088, in15088_1, in15088_2;
    wire c15088;
    assign in15088_1 = {s13718[0]};
    assign in15088_2 = {c14596};
    Full_Adder FA_15088(s15088, c15088, in15088_1, in15088_2, s13717[0]);
    wire[0:0] s15089, in15089_1, in15089_2;
    wire c15089;
    assign in15089_1 = {s14598[0]};
    assign in15089_2 = {s14599[0]};
    Full_Adder FA_15089(s15089, c15089, in15089_1, in15089_2, c14597);
    wire[0:0] s15090, in15090_1, in15090_2;
    wire c15090;
    assign in15090_1 = {s13722[0]};
    assign in15090_2 = {c14598};
    Full_Adder FA_15090(s15090, c15090, in15090_1, in15090_2, s13721[0]);
    wire[0:0] s15091, in15091_1, in15091_2;
    wire c15091;
    assign in15091_1 = {s14600[0]};
    assign in15091_2 = {s14601[0]};
    Full_Adder FA_15091(s15091, c15091, in15091_1, in15091_2, c14599);
    wire[0:0] s15092, in15092_1, in15092_2;
    wire c15092;
    assign in15092_1 = {s13726[0]};
    assign in15092_2 = {c14600};
    Full_Adder FA_15092(s15092, c15092, in15092_1, in15092_2, s13725[0]);
    wire[0:0] s15093, in15093_1, in15093_2;
    wire c15093;
    assign in15093_1 = {s14602[0]};
    assign in15093_2 = {s14603[0]};
    Full_Adder FA_15093(s15093, c15093, in15093_1, in15093_2, c14601);
    wire[0:0] s15094, in15094_1, in15094_2;
    wire c15094;
    assign in15094_1 = {s13730[0]};
    assign in15094_2 = {c14602};
    Full_Adder FA_15094(s15094, c15094, in15094_1, in15094_2, s13729[0]);
    wire[0:0] s15095, in15095_1, in15095_2;
    wire c15095;
    assign in15095_1 = {s14604[0]};
    assign in15095_2 = {s14605[0]};
    Full_Adder FA_15095(s15095, c15095, in15095_1, in15095_2, c14603);
    wire[0:0] s15096, in15096_1, in15096_2;
    wire c15096;
    assign in15096_1 = {s13734[0]};
    assign in15096_2 = {c14604};
    Full_Adder FA_15096(s15096, c15096, in15096_1, in15096_2, s13733[0]);
    wire[0:0] s15097, in15097_1, in15097_2;
    wire c15097;
    assign in15097_1 = {s14606[0]};
    assign in15097_2 = {s14607[0]};
    Full_Adder FA_15097(s15097, c15097, in15097_1, in15097_2, c14605);
    wire[0:0] s15098, in15098_1, in15098_2;
    wire c15098;
    assign in15098_1 = {s13738[0]};
    assign in15098_2 = {c14606};
    Full_Adder FA_15098(s15098, c15098, in15098_1, in15098_2, s13737[0]);
    wire[0:0] s15099, in15099_1, in15099_2;
    wire c15099;
    assign in15099_1 = {s14608[0]};
    assign in15099_2 = {s14609[0]};
    Full_Adder FA_15099(s15099, c15099, in15099_1, in15099_2, c14607);
    wire[0:0] s15100, in15100_1, in15100_2;
    wire c15100;
    assign in15100_1 = {s13742[0]};
    assign in15100_2 = {c14608};
    Full_Adder FA_15100(s15100, c15100, in15100_1, in15100_2, s13741[0]);
    wire[0:0] s15101, in15101_1, in15101_2;
    wire c15101;
    assign in15101_1 = {s14610[0]};
    assign in15101_2 = {s14611[0]};
    Full_Adder FA_15101(s15101, c15101, in15101_1, in15101_2, c14609);
    wire[0:0] s15102, in15102_1, in15102_2;
    wire c15102;
    assign in15102_1 = {s13746[0]};
    assign in15102_2 = {c14610};
    Full_Adder FA_15102(s15102, c15102, in15102_1, in15102_2, s13745[0]);
    wire[0:0] s15103, in15103_1, in15103_2;
    wire c15103;
    assign in15103_1 = {s14612[0]};
    assign in15103_2 = {s14613[0]};
    Full_Adder FA_15103(s15103, c15103, in15103_1, in15103_2, c14611);
    wire[0:0] s15104, in15104_1, in15104_2;
    wire c15104;
    assign in15104_1 = {s13750[0]};
    assign in15104_2 = {c14612};
    Full_Adder FA_15104(s15104, c15104, in15104_1, in15104_2, s13749[0]);
    wire[0:0] s15105, in15105_1, in15105_2;
    wire c15105;
    assign in15105_1 = {s14614[0]};
    assign in15105_2 = {s14615[0]};
    Full_Adder FA_15105(s15105, c15105, in15105_1, in15105_2, c14613);
    wire[0:0] s15106, in15106_1, in15106_2;
    wire c15106;
    assign in15106_1 = {s13754[0]};
    assign in15106_2 = {c14614};
    Full_Adder FA_15106(s15106, c15106, in15106_1, in15106_2, s13753[0]);
    wire[0:0] s15107, in15107_1, in15107_2;
    wire c15107;
    assign in15107_1 = {s14616[0]};
    assign in15107_2 = {s14617[0]};
    Full_Adder FA_15107(s15107, c15107, in15107_1, in15107_2, c14615);
    wire[0:0] s15108, in15108_1, in15108_2;
    wire c15108;
    assign in15108_1 = {s13758[0]};
    assign in15108_2 = {c14616};
    Full_Adder FA_15108(s15108, c15108, in15108_1, in15108_2, s13757[0]);
    wire[0:0] s15109, in15109_1, in15109_2;
    wire c15109;
    assign in15109_1 = {s14618[0]};
    assign in15109_2 = {s14619[0]};
    Full_Adder FA_15109(s15109, c15109, in15109_1, in15109_2, c14617);
    wire[0:0] s15110, in15110_1, in15110_2;
    wire c15110;
    assign in15110_1 = {s13762[0]};
    assign in15110_2 = {c14618};
    Full_Adder FA_15110(s15110, c15110, in15110_1, in15110_2, s13761[0]);
    wire[0:0] s15111, in15111_1, in15111_2;
    wire c15111;
    assign in15111_1 = {s14620[0]};
    assign in15111_2 = {s14621[0]};
    Full_Adder FA_15111(s15111, c15111, in15111_1, in15111_2, c14619);
    wire[0:0] s15112, in15112_1, in15112_2;
    wire c15112;
    assign in15112_1 = {s13766[0]};
    assign in15112_2 = {c14620};
    Full_Adder FA_15112(s15112, c15112, in15112_1, in15112_2, s13765[0]);
    wire[0:0] s15113, in15113_1, in15113_2;
    wire c15113;
    assign in15113_1 = {s14622[0]};
    assign in15113_2 = {s14623[0]};
    Full_Adder FA_15113(s15113, c15113, in15113_1, in15113_2, c14621);
    wire[0:0] s15114, in15114_1, in15114_2;
    wire c15114;
    assign in15114_1 = {s13770[0]};
    assign in15114_2 = {c14622};
    Full_Adder FA_15114(s15114, c15114, in15114_1, in15114_2, s13769[0]);
    wire[0:0] s15115, in15115_1, in15115_2;
    wire c15115;
    assign in15115_1 = {s14624[0]};
    assign in15115_2 = {s14625[0]};
    Full_Adder FA_15115(s15115, c15115, in15115_1, in15115_2, c14623);
    wire[0:0] s15116, in15116_1, in15116_2;
    wire c15116;
    assign in15116_1 = {s13774[0]};
    assign in15116_2 = {c14624};
    Full_Adder FA_15116(s15116, c15116, in15116_1, in15116_2, s13773[0]);
    wire[0:0] s15117, in15117_1, in15117_2;
    wire c15117;
    assign in15117_1 = {s14626[0]};
    assign in15117_2 = {s14627[0]};
    Full_Adder FA_15117(s15117, c15117, in15117_1, in15117_2, c14625);
    wire[0:0] s15118, in15118_1, in15118_2;
    wire c15118;
    assign in15118_1 = {s13778[0]};
    assign in15118_2 = {c14626};
    Full_Adder FA_15118(s15118, c15118, in15118_1, in15118_2, s13777[0]);
    wire[0:0] s15119, in15119_1, in15119_2;
    wire c15119;
    assign in15119_1 = {s14628[0]};
    assign in15119_2 = {s14629[0]};
    Full_Adder FA_15119(s15119, c15119, in15119_1, in15119_2, c14627);
    wire[0:0] s15120, in15120_1, in15120_2;
    wire c15120;
    assign in15120_1 = {s13782[0]};
    assign in15120_2 = {c14628};
    Full_Adder FA_15120(s15120, c15120, in15120_1, in15120_2, s13781[0]);
    wire[0:0] s15121, in15121_1, in15121_2;
    wire c15121;
    assign in15121_1 = {s14630[0]};
    assign in15121_2 = {s14631[0]};
    Full_Adder FA_15121(s15121, c15121, in15121_1, in15121_2, c14629);
    wire[0:0] s15122, in15122_1, in15122_2;
    wire c15122;
    assign in15122_1 = {s13786[0]};
    assign in15122_2 = {c14630};
    Full_Adder FA_15122(s15122, c15122, in15122_1, in15122_2, s13785[0]);
    wire[0:0] s15123, in15123_1, in15123_2;
    wire c15123;
    assign in15123_1 = {s14632[0]};
    assign in15123_2 = {s14633[0]};
    Full_Adder FA_15123(s15123, c15123, in15123_1, in15123_2, c14631);
    wire[0:0] s15124, in15124_1, in15124_2;
    wire c15124;
    assign in15124_1 = {s13790[0]};
    assign in15124_2 = {c14632};
    Full_Adder FA_15124(s15124, c15124, in15124_1, in15124_2, s13789[0]);
    wire[0:0] s15125, in15125_1, in15125_2;
    wire c15125;
    assign in15125_1 = {s14634[0]};
    assign in15125_2 = {s14635[0]};
    Full_Adder FA_15125(s15125, c15125, in15125_1, in15125_2, c14633);
    wire[0:0] s15126, in15126_1, in15126_2;
    wire c15126;
    assign in15126_1 = {s13794[0]};
    assign in15126_2 = {c14634};
    Full_Adder FA_15126(s15126, c15126, in15126_1, in15126_2, s13793[0]);
    wire[0:0] s15127, in15127_1, in15127_2;
    wire c15127;
    assign in15127_1 = {s14636[0]};
    assign in15127_2 = {s14637[0]};
    Full_Adder FA_15127(s15127, c15127, in15127_1, in15127_2, c14635);
    wire[0:0] s15128, in15128_1, in15128_2;
    wire c15128;
    assign in15128_1 = {s13798[0]};
    assign in15128_2 = {c14636};
    Full_Adder FA_15128(s15128, c15128, in15128_1, in15128_2, s13797[0]);
    wire[0:0] s15129, in15129_1, in15129_2;
    wire c15129;
    assign in15129_1 = {s14638[0]};
    assign in15129_2 = {s14639[0]};
    Full_Adder FA_15129(s15129, c15129, in15129_1, in15129_2, c14637);
    wire[0:0] s15130, in15130_1, in15130_2;
    wire c15130;
    assign in15130_1 = {s13802[0]};
    assign in15130_2 = {c14638};
    Full_Adder FA_15130(s15130, c15130, in15130_1, in15130_2, s13801[0]);
    wire[0:0] s15131, in15131_1, in15131_2;
    wire c15131;
    assign in15131_1 = {s14640[0]};
    assign in15131_2 = {s14641[0]};
    Full_Adder FA_15131(s15131, c15131, in15131_1, in15131_2, c14639);
    wire[0:0] s15132, in15132_1, in15132_2;
    wire c15132;
    assign in15132_1 = {s13806[0]};
    assign in15132_2 = {c14640};
    Full_Adder FA_15132(s15132, c15132, in15132_1, in15132_2, s13805[0]);
    wire[0:0] s15133, in15133_1, in15133_2;
    wire c15133;
    assign in15133_1 = {s14642[0]};
    assign in15133_2 = {s14643[0]};
    Full_Adder FA_15133(s15133, c15133, in15133_1, in15133_2, c14641);
    wire[0:0] s15134, in15134_1, in15134_2;
    wire c15134;
    assign in15134_1 = {s13810[0]};
    assign in15134_2 = {c14642};
    Full_Adder FA_15134(s15134, c15134, in15134_1, in15134_2, s13809[0]);
    wire[0:0] s15135, in15135_1, in15135_2;
    wire c15135;
    assign in15135_1 = {s14644[0]};
    assign in15135_2 = {s14645[0]};
    Full_Adder FA_15135(s15135, c15135, in15135_1, in15135_2, c14643);
    wire[0:0] s15136, in15136_1, in15136_2;
    wire c15136;
    assign in15136_1 = {s13814[0]};
    assign in15136_2 = {c14644};
    Full_Adder FA_15136(s15136, c15136, in15136_1, in15136_2, s13813[0]);
    wire[0:0] s15137, in15137_1, in15137_2;
    wire c15137;
    assign in15137_1 = {s14646[0]};
    assign in15137_2 = {s14647[0]};
    Full_Adder FA_15137(s15137, c15137, in15137_1, in15137_2, c14645);
    wire[0:0] s15138, in15138_1, in15138_2;
    wire c15138;
    assign in15138_1 = {s13818[0]};
    assign in15138_2 = {c14646};
    Full_Adder FA_15138(s15138, c15138, in15138_1, in15138_2, s13817[0]);
    wire[0:0] s15139, in15139_1, in15139_2;
    wire c15139;
    assign in15139_1 = {s14648[0]};
    assign in15139_2 = {s14649[0]};
    Full_Adder FA_15139(s15139, c15139, in15139_1, in15139_2, c14647);
    wire[0:0] s15140, in15140_1, in15140_2;
    wire c15140;
    assign in15140_1 = {s13822[0]};
    assign in15140_2 = {c14648};
    Full_Adder FA_15140(s15140, c15140, in15140_1, in15140_2, s13821[0]);
    wire[0:0] s15141, in15141_1, in15141_2;
    wire c15141;
    assign in15141_1 = {s14650[0]};
    assign in15141_2 = {s14651[0]};
    Full_Adder FA_15141(s15141, c15141, in15141_1, in15141_2, c14649);
    wire[0:0] s15142, in15142_1, in15142_2;
    wire c15142;
    assign in15142_1 = {s13826[0]};
    assign in15142_2 = {c14650};
    Full_Adder FA_15142(s15142, c15142, in15142_1, in15142_2, s13825[0]);
    wire[0:0] s15143, in15143_1, in15143_2;
    wire c15143;
    assign in15143_1 = {s14652[0]};
    assign in15143_2 = {s14653[0]};
    Full_Adder FA_15143(s15143, c15143, in15143_1, in15143_2, c14651);
    wire[0:0] s15144, in15144_1, in15144_2;
    wire c15144;
    assign in15144_1 = {s13830[0]};
    assign in15144_2 = {c14652};
    Full_Adder FA_15144(s15144, c15144, in15144_1, in15144_2, s13829[0]);
    wire[0:0] s15145, in15145_1, in15145_2;
    wire c15145;
    assign in15145_1 = {s14654[0]};
    assign in15145_2 = {s14655[0]};
    Full_Adder FA_15145(s15145, c15145, in15145_1, in15145_2, c14653);
    wire[0:0] s15146, in15146_1, in15146_2;
    wire c15146;
    assign in15146_1 = {s13834[0]};
    assign in15146_2 = {c14654};
    Full_Adder FA_15146(s15146, c15146, in15146_1, in15146_2, s13833[0]);
    wire[0:0] s15147, in15147_1, in15147_2;
    wire c15147;
    assign in15147_1 = {s14656[0]};
    assign in15147_2 = {s14657[0]};
    Full_Adder FA_15147(s15147, c15147, in15147_1, in15147_2, c14655);
    wire[0:0] s15148, in15148_1, in15148_2;
    wire c15148;
    assign in15148_1 = {s13838[0]};
    assign in15148_2 = {c14656};
    Full_Adder FA_15148(s15148, c15148, in15148_1, in15148_2, s13837[0]);
    wire[0:0] s15149, in15149_1, in15149_2;
    wire c15149;
    assign in15149_1 = {s14658[0]};
    assign in15149_2 = {s14659[0]};
    Full_Adder FA_15149(s15149, c15149, in15149_1, in15149_2, c14657);
    wire[0:0] s15150, in15150_1, in15150_2;
    wire c15150;
    assign in15150_1 = {s13842[0]};
    assign in15150_2 = {c14658};
    Full_Adder FA_15150(s15150, c15150, in15150_1, in15150_2, s13841[0]);
    wire[0:0] s15151, in15151_1, in15151_2;
    wire c15151;
    assign in15151_1 = {s14660[0]};
    assign in15151_2 = {s14661[0]};
    Full_Adder FA_15151(s15151, c15151, in15151_1, in15151_2, c14659);
    wire[0:0] s15152, in15152_1, in15152_2;
    wire c15152;
    assign in15152_1 = {s13846[0]};
    assign in15152_2 = {c14660};
    Full_Adder FA_15152(s15152, c15152, in15152_1, in15152_2, s13845[0]);
    wire[0:0] s15153, in15153_1, in15153_2;
    wire c15153;
    assign in15153_1 = {s14662[0]};
    assign in15153_2 = {s14663[0]};
    Full_Adder FA_15153(s15153, c15153, in15153_1, in15153_2, c14661);
    wire[0:0] s15154, in15154_1, in15154_2;
    wire c15154;
    assign in15154_1 = {s13850[0]};
    assign in15154_2 = {c14662};
    Full_Adder FA_15154(s15154, c15154, in15154_1, in15154_2, s13849[0]);
    wire[0:0] s15155, in15155_1, in15155_2;
    wire c15155;
    assign in15155_1 = {s14664[0]};
    assign in15155_2 = {s14665[0]};
    Full_Adder FA_15155(s15155, c15155, in15155_1, in15155_2, c14663);
    wire[0:0] s15156, in15156_1, in15156_2;
    wire c15156;
    assign in15156_1 = {s13854[0]};
    assign in15156_2 = {c14664};
    Full_Adder FA_15156(s15156, c15156, in15156_1, in15156_2, s13853[0]);
    wire[0:0] s15157, in15157_1, in15157_2;
    wire c15157;
    assign in15157_1 = {s14666[0]};
    assign in15157_2 = {s14667[0]};
    Full_Adder FA_15157(s15157, c15157, in15157_1, in15157_2, c14665);
    wire[0:0] s15158, in15158_1, in15158_2;
    wire c15158;
    assign in15158_1 = {s13858[0]};
    assign in15158_2 = {c14666};
    Full_Adder FA_15158(s15158, c15158, in15158_1, in15158_2, s13857[0]);
    wire[0:0] s15159, in15159_1, in15159_2;
    wire c15159;
    assign in15159_1 = {s14668[0]};
    assign in15159_2 = {s14669[0]};
    Full_Adder FA_15159(s15159, c15159, in15159_1, in15159_2, c14667);
    wire[0:0] s15160, in15160_1, in15160_2;
    wire c15160;
    assign in15160_1 = {s13862[0]};
    assign in15160_2 = {c14668};
    Full_Adder FA_15160(s15160, c15160, in15160_1, in15160_2, s13861[0]);
    wire[0:0] s15161, in15161_1, in15161_2;
    wire c15161;
    assign in15161_1 = {s14670[0]};
    assign in15161_2 = {s14671[0]};
    Full_Adder FA_15161(s15161, c15161, in15161_1, in15161_2, c14669);
    wire[0:0] s15162, in15162_1, in15162_2;
    wire c15162;
    assign in15162_1 = {s13866[0]};
    assign in15162_2 = {c14670};
    Full_Adder FA_15162(s15162, c15162, in15162_1, in15162_2, s13865[0]);
    wire[0:0] s15163, in15163_1, in15163_2;
    wire c15163;
    assign in15163_1 = {s14672[0]};
    assign in15163_2 = {s14673[0]};
    Full_Adder FA_15163(s15163, c15163, in15163_1, in15163_2, c14671);
    wire[0:0] s15164, in15164_1, in15164_2;
    wire c15164;
    assign in15164_1 = {s13870[0]};
    assign in15164_2 = {c14672};
    Full_Adder FA_15164(s15164, c15164, in15164_1, in15164_2, s13869[0]);
    wire[0:0] s15165, in15165_1, in15165_2;
    wire c15165;
    assign in15165_1 = {s14674[0]};
    assign in15165_2 = {s14675[0]};
    Full_Adder FA_15165(s15165, c15165, in15165_1, in15165_2, c14673);
    wire[0:0] s15166, in15166_1, in15166_2;
    wire c15166;
    assign in15166_1 = {s13874[0]};
    assign in15166_2 = {c14674};
    Full_Adder FA_15166(s15166, c15166, in15166_1, in15166_2, s13873[0]);
    wire[0:0] s15167, in15167_1, in15167_2;
    wire c15167;
    assign in15167_1 = {s14676[0]};
    assign in15167_2 = {s14677[0]};
    Full_Adder FA_15167(s15167, c15167, in15167_1, in15167_2, c14675);
    wire[0:0] s15168, in15168_1, in15168_2;
    wire c15168;
    assign in15168_1 = {s13878[0]};
    assign in15168_2 = {c14676};
    Full_Adder FA_15168(s15168, c15168, in15168_1, in15168_2, s13877[0]);
    wire[0:0] s15169, in15169_1, in15169_2;
    wire c15169;
    assign in15169_1 = {s14678[0]};
    assign in15169_2 = {s14679[0]};
    Full_Adder FA_15169(s15169, c15169, in15169_1, in15169_2, c14677);
    wire[0:0] s15170, in15170_1, in15170_2;
    wire c15170;
    assign in15170_1 = {s13882[0]};
    assign in15170_2 = {c14678};
    Full_Adder FA_15170(s15170, c15170, in15170_1, in15170_2, s13881[0]);
    wire[0:0] s15171, in15171_1, in15171_2;
    wire c15171;
    assign in15171_1 = {s14680[0]};
    assign in15171_2 = {s14681[0]};
    Full_Adder FA_15171(s15171, c15171, in15171_1, in15171_2, c14679);
    wire[0:0] s15172, in15172_1, in15172_2;
    wire c15172;
    assign in15172_1 = {s13886[0]};
    assign in15172_2 = {c14680};
    Full_Adder FA_15172(s15172, c15172, in15172_1, in15172_2, s13885[0]);
    wire[0:0] s15173, in15173_1, in15173_2;
    wire c15173;
    assign in15173_1 = {s14682[0]};
    assign in15173_2 = {s14683[0]};
    Full_Adder FA_15173(s15173, c15173, in15173_1, in15173_2, c14681);
    wire[0:0] s15174, in15174_1, in15174_2;
    wire c15174;
    assign in15174_1 = {s13890[0]};
    assign in15174_2 = {c14682};
    Full_Adder FA_15174(s15174, c15174, in15174_1, in15174_2, s13889[0]);
    wire[0:0] s15175, in15175_1, in15175_2;
    wire c15175;
    assign in15175_1 = {s14684[0]};
    assign in15175_2 = {s14685[0]};
    Full_Adder FA_15175(s15175, c15175, in15175_1, in15175_2, c14683);
    wire[0:0] s15176, in15176_1, in15176_2;
    wire c15176;
    assign in15176_1 = {s13894[0]};
    assign in15176_2 = {c14684};
    Full_Adder FA_15176(s15176, c15176, in15176_1, in15176_2, s13893[0]);
    wire[0:0] s15177, in15177_1, in15177_2;
    wire c15177;
    assign in15177_1 = {s14686[0]};
    assign in15177_2 = {s14687[0]};
    Full_Adder FA_15177(s15177, c15177, in15177_1, in15177_2, c14685);
    wire[0:0] s15178, in15178_1, in15178_2;
    wire c15178;
    assign in15178_1 = {s13898[0]};
    assign in15178_2 = {c14686};
    Full_Adder FA_15178(s15178, c15178, in15178_1, in15178_2, s13897[0]);
    wire[0:0] s15179, in15179_1, in15179_2;
    wire c15179;
    assign in15179_1 = {s14688[0]};
    assign in15179_2 = {s14689[0]};
    Full_Adder FA_15179(s15179, c15179, in15179_1, in15179_2, c14687);
    wire[0:0] s15180, in15180_1, in15180_2;
    wire c15180;
    assign in15180_1 = {s13902[0]};
    assign in15180_2 = {c14688};
    Full_Adder FA_15180(s15180, c15180, in15180_1, in15180_2, s13901[0]);
    wire[0:0] s15181, in15181_1, in15181_2;
    wire c15181;
    assign in15181_1 = {s14690[0]};
    assign in15181_2 = {s14691[0]};
    Full_Adder FA_15181(s15181, c15181, in15181_1, in15181_2, c14689);
    wire[0:0] s15182, in15182_1, in15182_2;
    wire c15182;
    assign in15182_1 = {s13906[0]};
    assign in15182_2 = {c14690};
    Full_Adder FA_15182(s15182, c15182, in15182_1, in15182_2, s13905[0]);
    wire[0:0] s15183, in15183_1, in15183_2;
    wire c15183;
    assign in15183_1 = {s14692[0]};
    assign in15183_2 = {s14693[0]};
    Full_Adder FA_15183(s15183, c15183, in15183_1, in15183_2, c14691);
    wire[0:0] s15184, in15184_1, in15184_2;
    wire c15184;
    assign in15184_1 = {s13910[0]};
    assign in15184_2 = {c14692};
    Full_Adder FA_15184(s15184, c15184, in15184_1, in15184_2, s13909[0]);
    wire[0:0] s15185, in15185_1, in15185_2;
    wire c15185;
    assign in15185_1 = {s14694[0]};
    assign in15185_2 = {s14695[0]};
    Full_Adder FA_15185(s15185, c15185, in15185_1, in15185_2, c14693);
    wire[0:0] s15186, in15186_1, in15186_2;
    wire c15186;
    assign in15186_1 = {s13914[0]};
    assign in15186_2 = {c14694};
    Full_Adder FA_15186(s15186, c15186, in15186_1, in15186_2, s13913[0]);
    wire[0:0] s15187, in15187_1, in15187_2;
    wire c15187;
    assign in15187_1 = {s14696[0]};
    assign in15187_2 = {s14697[0]};
    Full_Adder FA_15187(s15187, c15187, in15187_1, in15187_2, c14695);
    wire[0:0] s15188, in15188_1, in15188_2;
    wire c15188;
    assign in15188_1 = {s13918[0]};
    assign in15188_2 = {c14696};
    Full_Adder FA_15188(s15188, c15188, in15188_1, in15188_2, s13917[0]);
    wire[0:0] s15189, in15189_1, in15189_2;
    wire c15189;
    assign in15189_1 = {s14698[0]};
    assign in15189_2 = {s14699[0]};
    Full_Adder FA_15189(s15189, c15189, in15189_1, in15189_2, c14697);
    wire[0:0] s15190, in15190_1, in15190_2;
    wire c15190;
    assign in15190_1 = {s13922[0]};
    assign in15190_2 = {c14698};
    Full_Adder FA_15190(s15190, c15190, in15190_1, in15190_2, s13921[0]);
    wire[0:0] s15191, in15191_1, in15191_2;
    wire c15191;
    assign in15191_1 = {s14700[0]};
    assign in15191_2 = {s14701[0]};
    Full_Adder FA_15191(s15191, c15191, in15191_1, in15191_2, c14699);
    wire[0:0] s15192, in15192_1, in15192_2;
    wire c15192;
    assign in15192_1 = {s13926[0]};
    assign in15192_2 = {c14700};
    Full_Adder FA_15192(s15192, c15192, in15192_1, in15192_2, s13925[0]);
    wire[0:0] s15193, in15193_1, in15193_2;
    wire c15193;
    assign in15193_1 = {s14702[0]};
    assign in15193_2 = {s14703[0]};
    Full_Adder FA_15193(s15193, c15193, in15193_1, in15193_2, c14701);
    wire[0:0] s15194, in15194_1, in15194_2;
    wire c15194;
    assign in15194_1 = {s13930[0]};
    assign in15194_2 = {c14702};
    Full_Adder FA_15194(s15194, c15194, in15194_1, in15194_2, s13929[0]);
    wire[0:0] s15195, in15195_1, in15195_2;
    wire c15195;
    assign in15195_1 = {s14704[0]};
    assign in15195_2 = {s14705[0]};
    Full_Adder FA_15195(s15195, c15195, in15195_1, in15195_2, c14703);
    wire[0:0] s15196, in15196_1, in15196_2;
    wire c15196;
    assign in15196_1 = {s13934[0]};
    assign in15196_2 = {c14704};
    Full_Adder FA_15196(s15196, c15196, in15196_1, in15196_2, s13933[0]);
    wire[0:0] s15197, in15197_1, in15197_2;
    wire c15197;
    assign in15197_1 = {s14706[0]};
    assign in15197_2 = {s14707[0]};
    Full_Adder FA_15197(s15197, c15197, in15197_1, in15197_2, c14705);
    wire[0:0] s15198, in15198_1, in15198_2;
    wire c15198;
    assign in15198_1 = {s13938[0]};
    assign in15198_2 = {c14706};
    Full_Adder FA_15198(s15198, c15198, in15198_1, in15198_2, s13937[0]);
    wire[0:0] s15199, in15199_1, in15199_2;
    wire c15199;
    assign in15199_1 = {s14708[0]};
    assign in15199_2 = {s14709[0]};
    Full_Adder FA_15199(s15199, c15199, in15199_1, in15199_2, c14707);
    wire[0:0] s15200, in15200_1, in15200_2;
    wire c15200;
    assign in15200_1 = {s13942[0]};
    assign in15200_2 = {c14708};
    Full_Adder FA_15200(s15200, c15200, in15200_1, in15200_2, s13941[0]);
    wire[0:0] s15201, in15201_1, in15201_2;
    wire c15201;
    assign in15201_1 = {s14710[0]};
    assign in15201_2 = {s14711[0]};
    Full_Adder FA_15201(s15201, c15201, in15201_1, in15201_2, c14709);
    wire[0:0] s15202, in15202_1, in15202_2;
    wire c15202;
    assign in15202_1 = {s13946[0]};
    assign in15202_2 = {c14710};
    Full_Adder FA_15202(s15202, c15202, in15202_1, in15202_2, s13945[0]);
    wire[0:0] s15203, in15203_1, in15203_2;
    wire c15203;
    assign in15203_1 = {s14712[0]};
    assign in15203_2 = {s14713[0]};
    Full_Adder FA_15203(s15203, c15203, in15203_1, in15203_2, c14711);
    wire[0:0] s15204, in15204_1, in15204_2;
    wire c15204;
    assign in15204_1 = {s13950[0]};
    assign in15204_2 = {c14712};
    Full_Adder FA_15204(s15204, c15204, in15204_1, in15204_2, s13949[0]);
    wire[0:0] s15205, in15205_1, in15205_2;
    wire c15205;
    assign in15205_1 = {s14714[0]};
    assign in15205_2 = {s14715[0]};
    Full_Adder FA_15205(s15205, c15205, in15205_1, in15205_2, c14713);
    wire[0:0] s15206, in15206_1, in15206_2;
    wire c15206;
    assign in15206_1 = {s13954[0]};
    assign in15206_2 = {c14714};
    Full_Adder FA_15206(s15206, c15206, in15206_1, in15206_2, s13953[0]);
    wire[0:0] s15207, in15207_1, in15207_2;
    wire c15207;
    assign in15207_1 = {s14716[0]};
    assign in15207_2 = {s14717[0]};
    Full_Adder FA_15207(s15207, c15207, in15207_1, in15207_2, c14715);
    wire[0:0] s15208, in15208_1, in15208_2;
    wire c15208;
    assign in15208_1 = {s13958[0]};
    assign in15208_2 = {c14716};
    Full_Adder FA_15208(s15208, c15208, in15208_1, in15208_2, s13957[0]);
    wire[0:0] s15209, in15209_1, in15209_2;
    wire c15209;
    assign in15209_1 = {s14718[0]};
    assign in15209_2 = {s14719[0]};
    Full_Adder FA_15209(s15209, c15209, in15209_1, in15209_2, c14717);
    wire[0:0] s15210, in15210_1, in15210_2;
    wire c15210;
    assign in15210_1 = {s13962[0]};
    assign in15210_2 = {c14718};
    Full_Adder FA_15210(s15210, c15210, in15210_1, in15210_2, s13961[0]);
    wire[0:0] s15211, in15211_1, in15211_2;
    wire c15211;
    assign in15211_1 = {s14720[0]};
    assign in15211_2 = {s14721[0]};
    Full_Adder FA_15211(s15211, c15211, in15211_1, in15211_2, c14719);
    wire[0:0] s15212, in15212_1, in15212_2;
    wire c15212;
    assign in15212_1 = {s13966[0]};
    assign in15212_2 = {c14720};
    Full_Adder FA_15212(s15212, c15212, in15212_1, in15212_2, s13965[0]);
    wire[0:0] s15213, in15213_1, in15213_2;
    wire c15213;
    assign in15213_1 = {s14722[0]};
    assign in15213_2 = {s14723[0]};
    Full_Adder FA_15213(s15213, c15213, in15213_1, in15213_2, c14721);
    wire[0:0] s15214, in15214_1, in15214_2;
    wire c15214;
    assign in15214_1 = {s13970[0]};
    assign in15214_2 = {c14722};
    Full_Adder FA_15214(s15214, c15214, in15214_1, in15214_2, s13969[0]);
    wire[0:0] s15215, in15215_1, in15215_2;
    wire c15215;
    assign in15215_1 = {s14724[0]};
    assign in15215_2 = {s14725[0]};
    Full_Adder FA_15215(s15215, c15215, in15215_1, in15215_2, c14723);
    wire[0:0] s15216, in15216_1, in15216_2;
    wire c15216;
    assign in15216_1 = {s13974[0]};
    assign in15216_2 = {c14724};
    Full_Adder FA_15216(s15216, c15216, in15216_1, in15216_2, s13973[0]);
    wire[0:0] s15217, in15217_1, in15217_2;
    wire c15217;
    assign in15217_1 = {s14726[0]};
    assign in15217_2 = {s14727[0]};
    Full_Adder FA_15217(s15217, c15217, in15217_1, in15217_2, c14725);
    wire[0:0] s15218, in15218_1, in15218_2;
    wire c15218;
    assign in15218_1 = {s13978[0]};
    assign in15218_2 = {c14726};
    Full_Adder FA_15218(s15218, c15218, in15218_1, in15218_2, s13977[0]);
    wire[0:0] s15219, in15219_1, in15219_2;
    wire c15219;
    assign in15219_1 = {s14728[0]};
    assign in15219_2 = {s14729[0]};
    Full_Adder FA_15219(s15219, c15219, in15219_1, in15219_2, c14727);
    wire[0:0] s15220, in15220_1, in15220_2;
    wire c15220;
    assign in15220_1 = {s13982[0]};
    assign in15220_2 = {c14728};
    Full_Adder FA_15220(s15220, c15220, in15220_1, in15220_2, s13981[0]);
    wire[0:0] s15221, in15221_1, in15221_2;
    wire c15221;
    assign in15221_1 = {s14730[0]};
    assign in15221_2 = {s14731[0]};
    Full_Adder FA_15221(s15221, c15221, in15221_1, in15221_2, c14729);
    wire[0:0] s15222, in15222_1, in15222_2;
    wire c15222;
    assign in15222_1 = {s13986[0]};
    assign in15222_2 = {c14730};
    Full_Adder FA_15222(s15222, c15222, in15222_1, in15222_2, s13985[0]);
    wire[0:0] s15223, in15223_1, in15223_2;
    wire c15223;
    assign in15223_1 = {s14732[0]};
    assign in15223_2 = {s14733[0]};
    Full_Adder FA_15223(s15223, c15223, in15223_1, in15223_2, c14731);
    wire[0:0] s15224, in15224_1, in15224_2;
    wire c15224;
    assign in15224_1 = {s13990[0]};
    assign in15224_2 = {c14732};
    Full_Adder FA_15224(s15224, c15224, in15224_1, in15224_2, s13989[0]);
    wire[0:0] s15225, in15225_1, in15225_2;
    wire c15225;
    assign in15225_1 = {s14734[0]};
    assign in15225_2 = {s14735[0]};
    Full_Adder FA_15225(s15225, c15225, in15225_1, in15225_2, c14733);
    wire[0:0] s15226, in15226_1, in15226_2;
    wire c15226;
    assign in15226_1 = {s13994[0]};
    assign in15226_2 = {c14734};
    Full_Adder FA_15226(s15226, c15226, in15226_1, in15226_2, s13993[0]);
    wire[0:0] s15227, in15227_1, in15227_2;
    wire c15227;
    assign in15227_1 = {s14736[0]};
    assign in15227_2 = {s14737[0]};
    Full_Adder FA_15227(s15227, c15227, in15227_1, in15227_2, c14735);
    wire[0:0] s15228, in15228_1, in15228_2;
    wire c15228;
    assign in15228_1 = {s13998[0]};
    assign in15228_2 = {c14736};
    Full_Adder FA_15228(s15228, c15228, in15228_1, in15228_2, s13997[0]);
    wire[0:0] s15229, in15229_1, in15229_2;
    wire c15229;
    assign in15229_1 = {s14738[0]};
    assign in15229_2 = {s14739[0]};
    Full_Adder FA_15229(s15229, c15229, in15229_1, in15229_2, c14737);
    wire[0:0] s15230, in15230_1, in15230_2;
    wire c15230;
    assign in15230_1 = {s14002[0]};
    assign in15230_2 = {c14738};
    Full_Adder FA_15230(s15230, c15230, in15230_1, in15230_2, s14001[0]);
    wire[0:0] s15231, in15231_1, in15231_2;
    wire c15231;
    assign in15231_1 = {s14740[0]};
    assign in15231_2 = {s14741[0]};
    Full_Adder FA_15231(s15231, c15231, in15231_1, in15231_2, c14739);
    wire[0:0] s15232, in15232_1, in15232_2;
    wire c15232;
    assign in15232_1 = {s14006[0]};
    assign in15232_2 = {c14740};
    Full_Adder FA_15232(s15232, c15232, in15232_1, in15232_2, s14005[0]);
    wire[0:0] s15233, in15233_1, in15233_2;
    wire c15233;
    assign in15233_1 = {s14742[0]};
    assign in15233_2 = {s14743[0]};
    Full_Adder FA_15233(s15233, c15233, in15233_1, in15233_2, c14741);
    wire[0:0] s15234, in15234_1, in15234_2;
    wire c15234;
    assign in15234_1 = {s14010[0]};
    assign in15234_2 = {c14742};
    Full_Adder FA_15234(s15234, c15234, in15234_1, in15234_2, s14009[0]);
    wire[0:0] s15235, in15235_1, in15235_2;
    wire c15235;
    assign in15235_1 = {s14744[0]};
    assign in15235_2 = {s14745[0]};
    Full_Adder FA_15235(s15235, c15235, in15235_1, in15235_2, c14743);
    wire[0:0] s15236, in15236_1, in15236_2;
    wire c15236;
    assign in15236_1 = {s14014[0]};
    assign in15236_2 = {c14744};
    Full_Adder FA_15236(s15236, c15236, in15236_1, in15236_2, s14013[0]);
    wire[0:0] s15237, in15237_1, in15237_2;
    wire c15237;
    assign in15237_1 = {s14746[0]};
    assign in15237_2 = {s14747[0]};
    Full_Adder FA_15237(s15237, c15237, in15237_1, in15237_2, c14745);
    wire[0:0] s15238, in15238_1, in15238_2;
    wire c15238;
    assign in15238_1 = {s14018[0]};
    assign in15238_2 = {c14746};
    Full_Adder FA_15238(s15238, c15238, in15238_1, in15238_2, s14017[0]);
    wire[0:0] s15239, in15239_1, in15239_2;
    wire c15239;
    assign in15239_1 = {s14748[0]};
    assign in15239_2 = {s14749[0]};
    Full_Adder FA_15239(s15239, c15239, in15239_1, in15239_2, c14747);
    wire[0:0] s15240, in15240_1, in15240_2;
    wire c15240;
    assign in15240_1 = {s14022[0]};
    assign in15240_2 = {c14748};
    Full_Adder FA_15240(s15240, c15240, in15240_1, in15240_2, s14021[0]);
    wire[0:0] s15241, in15241_1, in15241_2;
    wire c15241;
    assign in15241_1 = {s14750[0]};
    assign in15241_2 = {s14751[0]};
    Full_Adder FA_15241(s15241, c15241, in15241_1, in15241_2, c14749);
    wire[0:0] s15242, in15242_1, in15242_2;
    wire c15242;
    assign in15242_1 = {s14026[0]};
    assign in15242_2 = {c14750};
    Full_Adder FA_15242(s15242, c15242, in15242_1, in15242_2, s14025[0]);
    wire[0:0] s15243, in15243_1, in15243_2;
    wire c15243;
    assign in15243_1 = {s14752[0]};
    assign in15243_2 = {s14753[0]};
    Full_Adder FA_15243(s15243, c15243, in15243_1, in15243_2, c14751);
    wire[0:0] s15244, in15244_1, in15244_2;
    wire c15244;
    assign in15244_1 = {s14030[0]};
    assign in15244_2 = {c14752};
    Full_Adder FA_15244(s15244, c15244, in15244_1, in15244_2, s14029[0]);
    wire[0:0] s15245, in15245_1, in15245_2;
    wire c15245;
    assign in15245_1 = {s14754[0]};
    assign in15245_2 = {s14755[0]};
    Full_Adder FA_15245(s15245, c15245, in15245_1, in15245_2, c14753);
    wire[0:0] s15246, in15246_1, in15246_2;
    wire c15246;
    assign in15246_1 = {s14034[0]};
    assign in15246_2 = {c14754};
    Full_Adder FA_15246(s15246, c15246, in15246_1, in15246_2, s14033[0]);
    wire[0:0] s15247, in15247_1, in15247_2;
    wire c15247;
    assign in15247_1 = {s14756[0]};
    assign in15247_2 = {s14757[0]};
    Full_Adder FA_15247(s15247, c15247, in15247_1, in15247_2, c14755);
    wire[0:0] s15248, in15248_1, in15248_2;
    wire c15248;
    assign in15248_1 = {s14038[0]};
    assign in15248_2 = {c14756};
    Full_Adder FA_15248(s15248, c15248, in15248_1, in15248_2, s14037[0]);
    wire[0:0] s15249, in15249_1, in15249_2;
    wire c15249;
    assign in15249_1 = {s14758[0]};
    assign in15249_2 = {s14759[0]};
    Full_Adder FA_15249(s15249, c15249, in15249_1, in15249_2, c14757);
    wire[0:0] s15250, in15250_1, in15250_2;
    wire c15250;
    assign in15250_1 = {s14042[0]};
    assign in15250_2 = {c14758};
    Full_Adder FA_15250(s15250, c15250, in15250_1, in15250_2, s14041[0]);
    wire[0:0] s15251, in15251_1, in15251_2;
    wire c15251;
    assign in15251_1 = {s14760[0]};
    assign in15251_2 = {s14761[0]};
    Full_Adder FA_15251(s15251, c15251, in15251_1, in15251_2, c14759);
    wire[0:0] s15252, in15252_1, in15252_2;
    wire c15252;
    assign in15252_1 = {s14046[0]};
    assign in15252_2 = {c14760};
    Full_Adder FA_15252(s15252, c15252, in15252_1, in15252_2, s14045[0]);
    wire[0:0] s15253, in15253_1, in15253_2;
    wire c15253;
    assign in15253_1 = {s14762[0]};
    assign in15253_2 = {s14763[0]};
    Full_Adder FA_15253(s15253, c15253, in15253_1, in15253_2, c14761);
    wire[0:0] s15254, in15254_1, in15254_2;
    wire c15254;
    assign in15254_1 = {s14050[0]};
    assign in15254_2 = {c14762};
    Full_Adder FA_15254(s15254, c15254, in15254_1, in15254_2, s14049[0]);
    wire[0:0] s15255, in15255_1, in15255_2;
    wire c15255;
    assign in15255_1 = {s14764[0]};
    assign in15255_2 = {s14765[0]};
    Full_Adder FA_15255(s15255, c15255, in15255_1, in15255_2, c14763);
    wire[0:0] s15256, in15256_1, in15256_2;
    wire c15256;
    assign in15256_1 = {s14054[0]};
    assign in15256_2 = {c14764};
    Full_Adder FA_15256(s15256, c15256, in15256_1, in15256_2, s14053[0]);
    wire[0:0] s15257, in15257_1, in15257_2;
    wire c15257;
    assign in15257_1 = {s14766[0]};
    assign in15257_2 = {s14767[0]};
    Full_Adder FA_15257(s15257, c15257, in15257_1, in15257_2, c14765);
    wire[0:0] s15258, in15258_1, in15258_2;
    wire c15258;
    assign in15258_1 = {s14058[0]};
    assign in15258_2 = {c14766};
    Full_Adder FA_15258(s15258, c15258, in15258_1, in15258_2, s14057[0]);
    wire[0:0] s15259, in15259_1, in15259_2;
    wire c15259;
    assign in15259_1 = {s14768[0]};
    assign in15259_2 = {s14769[0]};
    Full_Adder FA_15259(s15259, c15259, in15259_1, in15259_2, c14767);
    wire[0:0] s15260, in15260_1, in15260_2;
    wire c15260;
    assign in15260_1 = {s14062[0]};
    assign in15260_2 = {c14768};
    Full_Adder FA_15260(s15260, c15260, in15260_1, in15260_2, s14061[0]);
    wire[0:0] s15261, in15261_1, in15261_2;
    wire c15261;
    assign in15261_1 = {s14770[0]};
    assign in15261_2 = {s14771[0]};
    Full_Adder FA_15261(s15261, c15261, in15261_1, in15261_2, c14769);
    wire[0:0] s15262, in15262_1, in15262_2;
    wire c15262;
    assign in15262_1 = {s14066[0]};
    assign in15262_2 = {c14770};
    Full_Adder FA_15262(s15262, c15262, in15262_1, in15262_2, s14065[0]);
    wire[0:0] s15263, in15263_1, in15263_2;
    wire c15263;
    assign in15263_1 = {s14772[0]};
    assign in15263_2 = {s14773[0]};
    Full_Adder FA_15263(s15263, c15263, in15263_1, in15263_2, c14771);
    wire[0:0] s15264, in15264_1, in15264_2;
    wire c15264;
    assign in15264_1 = {s14070[0]};
    assign in15264_2 = {c14772};
    Full_Adder FA_15264(s15264, c15264, in15264_1, in15264_2, s14069[0]);
    wire[0:0] s15265, in15265_1, in15265_2;
    wire c15265;
    assign in15265_1 = {s14774[0]};
    assign in15265_2 = {s14775[0]};
    Full_Adder FA_15265(s15265, c15265, in15265_1, in15265_2, c14773);
    wire[0:0] s15266, in15266_1, in15266_2;
    wire c15266;
    assign in15266_1 = {s14074[0]};
    assign in15266_2 = {c14774};
    Full_Adder FA_15266(s15266, c15266, in15266_1, in15266_2, s14073[0]);
    wire[0:0] s15267, in15267_1, in15267_2;
    wire c15267;
    assign in15267_1 = {s14776[0]};
    assign in15267_2 = {s14777[0]};
    Full_Adder FA_15267(s15267, c15267, in15267_1, in15267_2, c14775);
    wire[0:0] s15268, in15268_1, in15268_2;
    wire c15268;
    assign in15268_1 = {s14078[0]};
    assign in15268_2 = {c14776};
    Full_Adder FA_15268(s15268, c15268, in15268_1, in15268_2, s14077[0]);
    wire[0:0] s15269, in15269_1, in15269_2;
    wire c15269;
    assign in15269_1 = {s14778[0]};
    assign in15269_2 = {s14779[0]};
    Full_Adder FA_15269(s15269, c15269, in15269_1, in15269_2, c14777);
    wire[0:0] s15270, in15270_1, in15270_2;
    wire c15270;
    assign in15270_1 = {s14082[0]};
    assign in15270_2 = {c14778};
    Full_Adder FA_15270(s15270, c15270, in15270_1, in15270_2, s14081[0]);
    wire[0:0] s15271, in15271_1, in15271_2;
    wire c15271;
    assign in15271_1 = {s14780[0]};
    assign in15271_2 = {s14781[0]};
    Full_Adder FA_15271(s15271, c15271, in15271_1, in15271_2, c14779);
    wire[0:0] s15272, in15272_1, in15272_2;
    wire c15272;
    assign in15272_1 = {s14086[0]};
    assign in15272_2 = {c14780};
    Full_Adder FA_15272(s15272, c15272, in15272_1, in15272_2, s14085[0]);
    wire[0:0] s15273, in15273_1, in15273_2;
    wire c15273;
    assign in15273_1 = {s14782[0]};
    assign in15273_2 = {s14783[0]};
    Full_Adder FA_15273(s15273, c15273, in15273_1, in15273_2, c14781);
    wire[0:0] s15274, in15274_1, in15274_2;
    wire c15274;
    assign in15274_1 = {s14090[0]};
    assign in15274_2 = {c14782};
    Full_Adder FA_15274(s15274, c15274, in15274_1, in15274_2, s14089[0]);
    wire[0:0] s15275, in15275_1, in15275_2;
    wire c15275;
    assign in15275_1 = {s14784[0]};
    assign in15275_2 = {s14785[0]};
    Full_Adder FA_15275(s15275, c15275, in15275_1, in15275_2, c14783);
    wire[0:0] s15276, in15276_1, in15276_2;
    wire c15276;
    assign in15276_1 = {s14094[0]};
    assign in15276_2 = {c14784};
    Full_Adder FA_15276(s15276, c15276, in15276_1, in15276_2, s14093[0]);
    wire[0:0] s15277, in15277_1, in15277_2;
    wire c15277;
    assign in15277_1 = {s14786[0]};
    assign in15277_2 = {s14787[0]};
    Full_Adder FA_15277(s15277, c15277, in15277_1, in15277_2, c14785);
    wire[0:0] s15278, in15278_1, in15278_2;
    wire c15278;
    assign in15278_1 = {s14098[0]};
    assign in15278_2 = {c14786};
    Full_Adder FA_15278(s15278, c15278, in15278_1, in15278_2, s14097[0]);
    wire[0:0] s15279, in15279_1, in15279_2;
    wire c15279;
    assign in15279_1 = {s14788[0]};
    assign in15279_2 = {s14789[0]};
    Full_Adder FA_15279(s15279, c15279, in15279_1, in15279_2, c14787);
    wire[0:0] s15280, in15280_1, in15280_2;
    wire c15280;
    assign in15280_1 = {s14102[0]};
    assign in15280_2 = {c14788};
    Full_Adder FA_15280(s15280, c15280, in15280_1, in15280_2, s14101[0]);
    wire[0:0] s15281, in15281_1, in15281_2;
    wire c15281;
    assign in15281_1 = {s14790[0]};
    assign in15281_2 = {s14791[0]};
    Full_Adder FA_15281(s15281, c15281, in15281_1, in15281_2, c14789);
    wire[0:0] s15282, in15282_1, in15282_2;
    wire c15282;
    assign in15282_1 = {s14106[0]};
    assign in15282_2 = {c14790};
    Full_Adder FA_15282(s15282, c15282, in15282_1, in15282_2, s14105[0]);
    wire[0:0] s15283, in15283_1, in15283_2;
    wire c15283;
    assign in15283_1 = {s14792[0]};
    assign in15283_2 = {s14793[0]};
    Full_Adder FA_15283(s15283, c15283, in15283_1, in15283_2, c14791);
    wire[0:0] s15284, in15284_1, in15284_2;
    wire c15284;
    assign in15284_1 = {s14110[0]};
    assign in15284_2 = {c14792};
    Full_Adder FA_15284(s15284, c15284, in15284_1, in15284_2, s14109[0]);
    wire[0:0] s15285, in15285_1, in15285_2;
    wire c15285;
    assign in15285_1 = {s14794[0]};
    assign in15285_2 = {s14795[0]};
    Full_Adder FA_15285(s15285, c15285, in15285_1, in15285_2, c14793);
    wire[0:0] s15286, in15286_1, in15286_2;
    wire c15286;
    assign in15286_1 = {s14114[0]};
    assign in15286_2 = {c14794};
    Full_Adder FA_15286(s15286, c15286, in15286_1, in15286_2, s14113[0]);
    wire[0:0] s15287, in15287_1, in15287_2;
    wire c15287;
    assign in15287_1 = {s14796[0]};
    assign in15287_2 = {s14797[0]};
    Full_Adder FA_15287(s15287, c15287, in15287_1, in15287_2, c14795);
    wire[0:0] s15288, in15288_1, in15288_2;
    wire c15288;
    assign in15288_1 = {s14118[0]};
    assign in15288_2 = {c14796};
    Full_Adder FA_15288(s15288, c15288, in15288_1, in15288_2, s14117[0]);
    wire[0:0] s15289, in15289_1, in15289_2;
    wire c15289;
    assign in15289_1 = {s14798[0]};
    assign in15289_2 = {s14799[0]};
    Full_Adder FA_15289(s15289, c15289, in15289_1, in15289_2, c14797);
    wire[0:0] s15290, in15290_1, in15290_2;
    wire c15290;
    assign in15290_1 = {s14122[0]};
    assign in15290_2 = {c14798};
    Full_Adder FA_15290(s15290, c15290, in15290_1, in15290_2, s14121[0]);
    wire[0:0] s15291, in15291_1, in15291_2;
    wire c15291;
    assign in15291_1 = {s14800[0]};
    assign in15291_2 = {s14801[0]};
    Full_Adder FA_15291(s15291, c15291, in15291_1, in15291_2, c14799);
    wire[0:0] s15292, in15292_1, in15292_2;
    wire c15292;
    assign in15292_1 = {s14126[0]};
    assign in15292_2 = {c14800};
    Full_Adder FA_15292(s15292, c15292, in15292_1, in15292_2, s14125[0]);
    wire[0:0] s15293, in15293_1, in15293_2;
    wire c15293;
    assign in15293_1 = {s14802[0]};
    assign in15293_2 = {s14803[0]};
    Full_Adder FA_15293(s15293, c15293, in15293_1, in15293_2, c14801);
    wire[0:0] s15294, in15294_1, in15294_2;
    wire c15294;
    assign in15294_1 = {s14130[0]};
    assign in15294_2 = {c14802};
    Full_Adder FA_15294(s15294, c15294, in15294_1, in15294_2, s14129[0]);
    wire[0:0] s15295, in15295_1, in15295_2;
    wire c15295;
    assign in15295_1 = {s14804[0]};
    assign in15295_2 = {s14805[0]};
    Full_Adder FA_15295(s15295, c15295, in15295_1, in15295_2, c14803);
    wire[0:0] s15296, in15296_1, in15296_2;
    wire c15296;
    assign in15296_1 = {s14134[0]};
    assign in15296_2 = {c14804};
    Full_Adder FA_15296(s15296, c15296, in15296_1, in15296_2, s14133[0]);
    wire[0:0] s15297, in15297_1, in15297_2;
    wire c15297;
    assign in15297_1 = {s14806[0]};
    assign in15297_2 = {s14807[0]};
    Full_Adder FA_15297(s15297, c15297, in15297_1, in15297_2, c14805);
    wire[0:0] s15298, in15298_1, in15298_2;
    wire c15298;
    assign in15298_1 = {s14138[0]};
    assign in15298_2 = {c14806};
    Full_Adder FA_15298(s15298, c15298, in15298_1, in15298_2, s14137[0]);
    wire[0:0] s15299, in15299_1, in15299_2;
    wire c15299;
    assign in15299_1 = {s14808[0]};
    assign in15299_2 = {s14809[0]};
    Full_Adder FA_15299(s15299, c15299, in15299_1, in15299_2, c14807);
    wire[0:0] s15300, in15300_1, in15300_2;
    wire c15300;
    assign in15300_1 = {s14142[0]};
    assign in15300_2 = {c14808};
    Full_Adder FA_15300(s15300, c15300, in15300_1, in15300_2, s14141[0]);
    wire[0:0] s15301, in15301_1, in15301_2;
    wire c15301;
    assign in15301_1 = {s14810[0]};
    assign in15301_2 = {s14811[0]};
    Full_Adder FA_15301(s15301, c15301, in15301_1, in15301_2, c14809);
    wire[0:0] s15302, in15302_1, in15302_2;
    wire c15302;
    assign in15302_1 = {s14146[0]};
    assign in15302_2 = {c14810};
    Full_Adder FA_15302(s15302, c15302, in15302_1, in15302_2, s14145[0]);
    wire[0:0] s15303, in15303_1, in15303_2;
    wire c15303;
    assign in15303_1 = {s14812[0]};
    assign in15303_2 = {s14813[0]};
    Full_Adder FA_15303(s15303, c15303, in15303_1, in15303_2, c14811);
    wire[0:0] s15304, in15304_1, in15304_2;
    wire c15304;
    assign in15304_1 = {s14150[0]};
    assign in15304_2 = {c14812};
    Full_Adder FA_15304(s15304, c15304, in15304_1, in15304_2, s14149[0]);
    wire[0:0] s15305, in15305_1, in15305_2;
    wire c15305;
    assign in15305_1 = {s14814[0]};
    assign in15305_2 = {s14815[0]};
    Full_Adder FA_15305(s15305, c15305, in15305_1, in15305_2, c14813);
    wire[0:0] s15306, in15306_1, in15306_2;
    wire c15306;
    assign in15306_1 = {s14154[0]};
    assign in15306_2 = {c14814};
    Full_Adder FA_15306(s15306, c15306, in15306_1, in15306_2, s14153[0]);
    wire[0:0] s15307, in15307_1, in15307_2;
    wire c15307;
    assign in15307_1 = {s14816[0]};
    assign in15307_2 = {s14817[0]};
    Full_Adder FA_15307(s15307, c15307, in15307_1, in15307_2, c14815);
    wire[0:0] s15308, in15308_1, in15308_2;
    wire c15308;
    assign in15308_1 = {s14158[0]};
    assign in15308_2 = {c14816};
    Full_Adder FA_15308(s15308, c15308, in15308_1, in15308_2, s14157[0]);
    wire[0:0] s15309, in15309_1, in15309_2;
    wire c15309;
    assign in15309_1 = {s14818[0]};
    assign in15309_2 = {s14819[0]};
    Full_Adder FA_15309(s15309, c15309, in15309_1, in15309_2, c14817);
    wire[0:0] s15310, in15310_1, in15310_2;
    wire c15310;
    assign in15310_1 = {s14162[0]};
    assign in15310_2 = {c14818};
    Full_Adder FA_15310(s15310, c15310, in15310_1, in15310_2, s14161[0]);
    wire[0:0] s15311, in15311_1, in15311_2;
    wire c15311;
    assign in15311_1 = {s14820[0]};
    assign in15311_2 = {s14821[0]};
    Full_Adder FA_15311(s15311, c15311, in15311_1, in15311_2, c14819);
    wire[0:0] s15312, in15312_1, in15312_2;
    wire c15312;
    assign in15312_1 = {s14166[0]};
    assign in15312_2 = {c14820};
    Full_Adder FA_15312(s15312, c15312, in15312_1, in15312_2, s14165[0]);
    wire[0:0] s15313, in15313_1, in15313_2;
    wire c15313;
    assign in15313_1 = {s14822[0]};
    assign in15313_2 = {s14823[0]};
    Full_Adder FA_15313(s15313, c15313, in15313_1, in15313_2, c14821);
    wire[0:0] s15314, in15314_1, in15314_2;
    wire c15314;
    assign in15314_1 = {s14170[0]};
    assign in15314_2 = {c14822};
    Full_Adder FA_15314(s15314, c15314, in15314_1, in15314_2, s14169[0]);
    wire[0:0] s15315, in15315_1, in15315_2;
    wire c15315;
    assign in15315_1 = {s14824[0]};
    assign in15315_2 = {s14825[0]};
    Full_Adder FA_15315(s15315, c15315, in15315_1, in15315_2, c14823);
    wire[0:0] s15316, in15316_1, in15316_2;
    wire c15316;
    assign in15316_1 = {s14174[0]};
    assign in15316_2 = {c14824};
    Full_Adder FA_15316(s15316, c15316, in15316_1, in15316_2, s14173[0]);
    wire[0:0] s15317, in15317_1, in15317_2;
    wire c15317;
    assign in15317_1 = {s14826[0]};
    assign in15317_2 = {s14827[0]};
    Full_Adder FA_15317(s15317, c15317, in15317_1, in15317_2, c14825);
    wire[0:0] s15318, in15318_1, in15318_2;
    wire c15318;
    assign in15318_1 = {s14178[0]};
    assign in15318_2 = {c14826};
    Full_Adder FA_15318(s15318, c15318, in15318_1, in15318_2, s14177[0]);
    wire[0:0] s15319, in15319_1, in15319_2;
    wire c15319;
    assign in15319_1 = {s14828[0]};
    assign in15319_2 = {s14829[0]};
    Full_Adder FA_15319(s15319, c15319, in15319_1, in15319_2, c14827);
    wire[0:0] s15320, in15320_1, in15320_2;
    wire c15320;
    assign in15320_1 = {s14182[0]};
    assign in15320_2 = {c14828};
    Full_Adder FA_15320(s15320, c15320, in15320_1, in15320_2, s14181[0]);
    wire[0:0] s15321, in15321_1, in15321_2;
    wire c15321;
    assign in15321_1 = {s14830[0]};
    assign in15321_2 = {s14831[0]};
    Full_Adder FA_15321(s15321, c15321, in15321_1, in15321_2, c14829);
    wire[0:0] s15322, in15322_1, in15322_2;
    wire c15322;
    assign in15322_1 = {s14186[0]};
    assign in15322_2 = {c14830};
    Full_Adder FA_15322(s15322, c15322, in15322_1, in15322_2, s14185[0]);
    wire[0:0] s15323, in15323_1, in15323_2;
    wire c15323;
    assign in15323_1 = {s14832[0]};
    assign in15323_2 = {s14833[0]};
    Full_Adder FA_15323(s15323, c15323, in15323_1, in15323_2, c14831);
    wire[0:0] s15324, in15324_1, in15324_2;
    wire c15324;
    assign in15324_1 = {s14190[0]};
    assign in15324_2 = {c14832};
    Full_Adder FA_15324(s15324, c15324, in15324_1, in15324_2, s14189[0]);
    wire[0:0] s15325, in15325_1, in15325_2;
    wire c15325;
    assign in15325_1 = {s14834[0]};
    assign in15325_2 = {s14835[0]};
    Full_Adder FA_15325(s15325, c15325, in15325_1, in15325_2, c14833);
    wire[0:0] s15326, in15326_1, in15326_2;
    wire c15326;
    assign in15326_1 = {s14194[0]};
    assign in15326_2 = {c14834};
    Full_Adder FA_15326(s15326, c15326, in15326_1, in15326_2, s14193[0]);
    wire[0:0] s15327, in15327_1, in15327_2;
    wire c15327;
    assign in15327_1 = {s14836[0]};
    assign in15327_2 = {s14837[0]};
    Full_Adder FA_15327(s15327, c15327, in15327_1, in15327_2, c14835);
    wire[0:0] s15328, in15328_1, in15328_2;
    wire c15328;
    assign in15328_1 = {s14198[0]};
    assign in15328_2 = {c14836};
    Full_Adder FA_15328(s15328, c15328, in15328_1, in15328_2, s14197[0]);
    wire[0:0] s15329, in15329_1, in15329_2;
    wire c15329;
    assign in15329_1 = {s14838[0]};
    assign in15329_2 = {s14839[0]};
    Full_Adder FA_15329(s15329, c15329, in15329_1, in15329_2, c14837);
    wire[0:0] s15330, in15330_1, in15330_2;
    wire c15330;
    assign in15330_1 = {s14202[0]};
    assign in15330_2 = {c14838};
    Full_Adder FA_15330(s15330, c15330, in15330_1, in15330_2, s14201[0]);
    wire[0:0] s15331, in15331_1, in15331_2;
    wire c15331;
    assign in15331_1 = {s14840[0]};
    assign in15331_2 = {s14841[0]};
    Full_Adder FA_15331(s15331, c15331, in15331_1, in15331_2, c14839);
    wire[0:0] s15332, in15332_1, in15332_2;
    wire c15332;
    assign in15332_1 = {s14206[0]};
    assign in15332_2 = {c14840};
    Full_Adder FA_15332(s15332, c15332, in15332_1, in15332_2, s14205[0]);
    wire[0:0] s15333, in15333_1, in15333_2;
    wire c15333;
    assign in15333_1 = {s14842[0]};
    assign in15333_2 = {s14843[0]};
    Full_Adder FA_15333(s15333, c15333, in15333_1, in15333_2, c14841);
    wire[0:0] s15334, in15334_1, in15334_2;
    wire c15334;
    assign in15334_1 = {s14210[0]};
    assign in15334_2 = {c14842};
    Full_Adder FA_15334(s15334, c15334, in15334_1, in15334_2, s14209[0]);
    wire[0:0] s15335, in15335_1, in15335_2;
    wire c15335;
    assign in15335_1 = {s14844[0]};
    assign in15335_2 = {s14845[0]};
    Full_Adder FA_15335(s15335, c15335, in15335_1, in15335_2, c14843);
    wire[0:0] s15336, in15336_1, in15336_2;
    wire c15336;
    assign in15336_1 = {s14214[0]};
    assign in15336_2 = {c14844};
    Full_Adder FA_15336(s15336, c15336, in15336_1, in15336_2, s14213[0]);
    wire[0:0] s15337, in15337_1, in15337_2;
    wire c15337;
    assign in15337_1 = {s14846[0]};
    assign in15337_2 = {s14847[0]};
    Full_Adder FA_15337(s15337, c15337, in15337_1, in15337_2, c14845);
    wire[0:0] s15338, in15338_1, in15338_2;
    wire c15338;
    assign in15338_1 = {s14218[0]};
    assign in15338_2 = {c14846};
    Full_Adder FA_15338(s15338, c15338, in15338_1, in15338_2, s14217[0]);
    wire[0:0] s15339, in15339_1, in15339_2;
    wire c15339;
    assign in15339_1 = {s14848[0]};
    assign in15339_2 = {s14849[0]};
    Full_Adder FA_15339(s15339, c15339, in15339_1, in15339_2, c14847);
    wire[0:0] s15340, in15340_1, in15340_2;
    wire c15340;
    assign in15340_1 = {s14222[0]};
    assign in15340_2 = {c14848};
    Full_Adder FA_15340(s15340, c15340, in15340_1, in15340_2, s14221[0]);
    wire[0:0] s15341, in15341_1, in15341_2;
    wire c15341;
    assign in15341_1 = {s14850[0]};
    assign in15341_2 = {s14851[0]};
    Full_Adder FA_15341(s15341, c15341, in15341_1, in15341_2, c14849);
    wire[0:0] s15342, in15342_1, in15342_2;
    wire c15342;
    assign in15342_1 = {s14226[0]};
    assign in15342_2 = {c14850};
    Full_Adder FA_15342(s15342, c15342, in15342_1, in15342_2, s14225[0]);
    wire[0:0] s15343, in15343_1, in15343_2;
    wire c15343;
    assign in15343_1 = {s14852[0]};
    assign in15343_2 = {s14853[0]};
    Full_Adder FA_15343(s15343, c15343, in15343_1, in15343_2, c14851);
    wire[0:0] s15344, in15344_1, in15344_2;
    wire c15344;
    assign in15344_1 = {s14230[0]};
    assign in15344_2 = {c14852};
    Full_Adder FA_15344(s15344, c15344, in15344_1, in15344_2, s14229[0]);
    wire[0:0] s15345, in15345_1, in15345_2;
    wire c15345;
    assign in15345_1 = {s14854[0]};
    assign in15345_2 = {s14855[0]};
    Full_Adder FA_15345(s15345, c15345, in15345_1, in15345_2, c14853);
    wire[0:0] s15346, in15346_1, in15346_2;
    wire c15346;
    assign in15346_1 = {s14234[0]};
    assign in15346_2 = {c14854};
    Full_Adder FA_15346(s15346, c15346, in15346_1, in15346_2, s14233[0]);
    wire[0:0] s15347, in15347_1, in15347_2;
    wire c15347;
    assign in15347_1 = {s14856[0]};
    assign in15347_2 = {s14857[0]};
    Full_Adder FA_15347(s15347, c15347, in15347_1, in15347_2, c14855);
    wire[0:0] s15348, in15348_1, in15348_2;
    wire c15348;
    assign in15348_1 = {s14238[0]};
    assign in15348_2 = {c14856};
    Full_Adder FA_15348(s15348, c15348, in15348_1, in15348_2, s14237[0]);
    wire[0:0] s15349, in15349_1, in15349_2;
    wire c15349;
    assign in15349_1 = {s14858[0]};
    assign in15349_2 = {s14859[0]};
    Full_Adder FA_15349(s15349, c15349, in15349_1, in15349_2, c14857);
    wire[0:0] s15350, in15350_1, in15350_2;
    wire c15350;
    assign in15350_1 = {s14242[0]};
    assign in15350_2 = {c14858};
    Full_Adder FA_15350(s15350, c15350, in15350_1, in15350_2, s14241[0]);
    wire[0:0] s15351, in15351_1, in15351_2;
    wire c15351;
    assign in15351_1 = {s14860[0]};
    assign in15351_2 = {s14861[0]};
    Full_Adder FA_15351(s15351, c15351, in15351_1, in15351_2, c14859);
    wire[0:0] s15352, in15352_1, in15352_2;
    wire c15352;
    assign in15352_1 = {s14246[0]};
    assign in15352_2 = {c14860};
    Full_Adder FA_15352(s15352, c15352, in15352_1, in15352_2, s14245[0]);
    wire[0:0] s15353, in15353_1, in15353_2;
    wire c15353;
    assign in15353_1 = {s14862[0]};
    assign in15353_2 = {s14863[0]};
    Full_Adder FA_15353(s15353, c15353, in15353_1, in15353_2, c14861);
    wire[0:0] s15354, in15354_1, in15354_2;
    wire c15354;
    assign in15354_1 = {s14250[0]};
    assign in15354_2 = {c14862};
    Full_Adder FA_15354(s15354, c15354, in15354_1, in15354_2, s14249[0]);
    wire[0:0] s15355, in15355_1, in15355_2;
    wire c15355;
    assign in15355_1 = {s14864[0]};
    assign in15355_2 = {s14865[0]};
    Full_Adder FA_15355(s15355, c15355, in15355_1, in15355_2, c14863);
    wire[0:0] s15356, in15356_1, in15356_2;
    wire c15356;
    assign in15356_1 = {s14254[0]};
    assign in15356_2 = {c14864};
    Full_Adder FA_15356(s15356, c15356, in15356_1, in15356_2, s14253[0]);
    wire[0:0] s15357, in15357_1, in15357_2;
    wire c15357;
    assign in15357_1 = {s14866[0]};
    assign in15357_2 = {s14867[0]};
    Full_Adder FA_15357(s15357, c15357, in15357_1, in15357_2, c14865);
    wire[0:0] s15358, in15358_1, in15358_2;
    wire c15358;
    assign in15358_1 = {s14258[0]};
    assign in15358_2 = {c14866};
    Full_Adder FA_15358(s15358, c15358, in15358_1, in15358_2, s14257[0]);
    wire[0:0] s15359, in15359_1, in15359_2;
    wire c15359;
    assign in15359_1 = {s14868[0]};
    assign in15359_2 = {s14869[0]};
    Full_Adder FA_15359(s15359, c15359, in15359_1, in15359_2, c14867);
    wire[0:0] s15360, in15360_1, in15360_2;
    wire c15360;
    assign in15360_1 = {s14262[0]};
    assign in15360_2 = {c14868};
    Full_Adder FA_15360(s15360, c15360, in15360_1, in15360_2, s14261[0]);
    wire[0:0] s15361, in15361_1, in15361_2;
    wire c15361;
    assign in15361_1 = {s14870[0]};
    assign in15361_2 = {s14871[0]};
    Full_Adder FA_15361(s15361, c15361, in15361_1, in15361_2, c14869);
    wire[0:0] s15362, in15362_1, in15362_2;
    wire c15362;
    assign in15362_1 = {s14266[0]};
    assign in15362_2 = {c14870};
    Full_Adder FA_15362(s15362, c15362, in15362_1, in15362_2, s14265[0]);
    wire[0:0] s15363, in15363_1, in15363_2;
    wire c15363;
    assign in15363_1 = {s14872[0]};
    assign in15363_2 = {s14873[0]};
    Full_Adder FA_15363(s15363, c15363, in15363_1, in15363_2, c14871);
    wire[0:0] s15364, in15364_1, in15364_2;
    wire c15364;
    assign in15364_1 = {s14270[0]};
    assign in15364_2 = {c14872};
    Full_Adder FA_15364(s15364, c15364, in15364_1, in15364_2, s14269[0]);
    wire[0:0] s15365, in15365_1, in15365_2;
    wire c15365;
    assign in15365_1 = {s14874[0]};
    assign in15365_2 = {s14875[0]};
    Full_Adder FA_15365(s15365, c15365, in15365_1, in15365_2, c14873);
    wire[0:0] s15366, in15366_1, in15366_2;
    wire c15366;
    assign in15366_1 = {s14274[0]};
    assign in15366_2 = {c14874};
    Full_Adder FA_15366(s15366, c15366, in15366_1, in15366_2, s14273[0]);
    wire[0:0] s15367, in15367_1, in15367_2;
    wire c15367;
    assign in15367_1 = {s14876[0]};
    assign in15367_2 = {s14877[0]};
    Full_Adder FA_15367(s15367, c15367, in15367_1, in15367_2, c14875);
    wire[0:0] s15368, in15368_1, in15368_2;
    wire c15368;
    assign in15368_1 = {s14278[0]};
    assign in15368_2 = {c14876};
    Full_Adder FA_15368(s15368, c15368, in15368_1, in15368_2, s14277[0]);
    wire[0:0] s15369, in15369_1, in15369_2;
    wire c15369;
    assign in15369_1 = {s14878[0]};
    assign in15369_2 = {s14879[0]};
    Full_Adder FA_15369(s15369, c15369, in15369_1, in15369_2, c14877);
    wire[0:0] s15370, in15370_1, in15370_2;
    wire c15370;
    assign in15370_1 = {s14282[0]};
    assign in15370_2 = {c14878};
    Full_Adder FA_15370(s15370, c15370, in15370_1, in15370_2, s14281[0]);
    wire[0:0] s15371, in15371_1, in15371_2;
    wire c15371;
    assign in15371_1 = {s14880[0]};
    assign in15371_2 = {s14881[0]};
    Full_Adder FA_15371(s15371, c15371, in15371_1, in15371_2, c14879);
    wire[0:0] s15372, in15372_1, in15372_2;
    wire c15372;
    assign in15372_1 = {s14286[0]};
    assign in15372_2 = {c14880};
    Full_Adder FA_15372(s15372, c15372, in15372_1, in15372_2, s14285[0]);
    wire[0:0] s15373, in15373_1, in15373_2;
    wire c15373;
    assign in15373_1 = {s14882[0]};
    assign in15373_2 = {s14883[0]};
    Full_Adder FA_15373(s15373, c15373, in15373_1, in15373_2, c14881);
    wire[0:0] s15374, in15374_1, in15374_2;
    wire c15374;
    assign in15374_1 = {s14290[0]};
    assign in15374_2 = {c14882};
    Full_Adder FA_15374(s15374, c15374, in15374_1, in15374_2, s14289[0]);
    wire[0:0] s15375, in15375_1, in15375_2;
    wire c15375;
    assign in15375_1 = {s14884[0]};
    assign in15375_2 = {s14885[0]};
    Full_Adder FA_15375(s15375, c15375, in15375_1, in15375_2, c14883);
    wire[0:0] s15376, in15376_1, in15376_2;
    wire c15376;
    assign in15376_1 = {s14294[0]};
    assign in15376_2 = {c14884};
    Full_Adder FA_15376(s15376, c15376, in15376_1, in15376_2, s14293[0]);
    wire[0:0] s15377, in15377_1, in15377_2;
    wire c15377;
    assign in15377_1 = {s14886[0]};
    assign in15377_2 = {s14887[0]};
    Full_Adder FA_15377(s15377, c15377, in15377_1, in15377_2, c14885);
    wire[0:0] s15378, in15378_1, in15378_2;
    wire c15378;
    assign in15378_1 = {s14298[0]};
    assign in15378_2 = {c14886};
    Full_Adder FA_15378(s15378, c15378, in15378_1, in15378_2, s14297[0]);
    wire[0:0] s15379, in15379_1, in15379_2;
    wire c15379;
    assign in15379_1 = {s14888[0]};
    assign in15379_2 = {s14889[0]};
    Full_Adder FA_15379(s15379, c15379, in15379_1, in15379_2, c14887);
    wire[0:0] s15380, in15380_1, in15380_2;
    wire c15380;
    assign in15380_1 = {s14302[0]};
    assign in15380_2 = {c14888};
    Full_Adder FA_15380(s15380, c15380, in15380_1, in15380_2, s14301[0]);
    wire[0:0] s15381, in15381_1, in15381_2;
    wire c15381;
    assign in15381_1 = {s14890[0]};
    assign in15381_2 = {s14891[0]};
    Full_Adder FA_15381(s15381, c15381, in15381_1, in15381_2, c14889);
    wire[0:0] s15382, in15382_1, in15382_2;
    wire c15382;
    assign in15382_1 = {s14306[0]};
    assign in15382_2 = {c14890};
    Full_Adder FA_15382(s15382, c15382, in15382_1, in15382_2, s14305[0]);
    wire[0:0] s15383, in15383_1, in15383_2;
    wire c15383;
    assign in15383_1 = {s14892[0]};
    assign in15383_2 = {s14893[0]};
    Full_Adder FA_15383(s15383, c15383, in15383_1, in15383_2, c14891);
    wire[0:0] s15384, in15384_1, in15384_2;
    wire c15384;
    assign in15384_1 = {s14310[0]};
    assign in15384_2 = {c14892};
    Full_Adder FA_15384(s15384, c15384, in15384_1, in15384_2, s14309[0]);
    wire[0:0] s15385, in15385_1, in15385_2;
    wire c15385;
    assign in15385_1 = {s14894[0]};
    assign in15385_2 = {s14895[0]};
    Full_Adder FA_15385(s15385, c15385, in15385_1, in15385_2, c14893);
    wire[0:0] s15386, in15386_1, in15386_2;
    wire c15386;
    assign in15386_1 = {s14314[0]};
    assign in15386_2 = {c14894};
    Full_Adder FA_15386(s15386, c15386, in15386_1, in15386_2, s14313[0]);
    wire[0:0] s15387, in15387_1, in15387_2;
    wire c15387;
    assign in15387_1 = {s14896[0]};
    assign in15387_2 = {s14897[0]};
    Full_Adder FA_15387(s15387, c15387, in15387_1, in15387_2, c14895);
    wire[0:0] s15388, in15388_1, in15388_2;
    wire c15388;
    assign in15388_1 = {s14318[0]};
    assign in15388_2 = {c14896};
    Full_Adder FA_15388(s15388, c15388, in15388_1, in15388_2, s14317[0]);
    wire[0:0] s15389, in15389_1, in15389_2;
    wire c15389;
    assign in15389_1 = {s14898[0]};
    assign in15389_2 = {s14899[0]};
    Full_Adder FA_15389(s15389, c15389, in15389_1, in15389_2, c14897);
    wire[0:0] s15390, in15390_1, in15390_2;
    wire c15390;
    assign in15390_1 = {s14322[0]};
    assign in15390_2 = {c14898};
    Full_Adder FA_15390(s15390, c15390, in15390_1, in15390_2, s14321[0]);
    wire[0:0] s15391, in15391_1, in15391_2;
    wire c15391;
    assign in15391_1 = {s14900[0]};
    assign in15391_2 = {s14901[0]};
    Full_Adder FA_15391(s15391, c15391, in15391_1, in15391_2, c14899);
    wire[0:0] s15392, in15392_1, in15392_2;
    wire c15392;
    assign in15392_1 = {s14326[0]};
    assign in15392_2 = {c14900};
    Full_Adder FA_15392(s15392, c15392, in15392_1, in15392_2, s14325[0]);
    wire[0:0] s15393, in15393_1, in15393_2;
    wire c15393;
    assign in15393_1 = {s14902[0]};
    assign in15393_2 = {s14903[0]};
    Full_Adder FA_15393(s15393, c15393, in15393_1, in15393_2, c14901);
    wire[0:0] s15394, in15394_1, in15394_2;
    wire c15394;
    assign in15394_1 = {s14330[0]};
    assign in15394_2 = {c14902};
    Full_Adder FA_15394(s15394, c15394, in15394_1, in15394_2, s14329[0]);
    wire[0:0] s15395, in15395_1, in15395_2;
    wire c15395;
    assign in15395_1 = {s14904[0]};
    assign in15395_2 = {s14905[0]};
    Full_Adder FA_15395(s15395, c15395, in15395_1, in15395_2, c14903);
    wire[0:0] s15396, in15396_1, in15396_2;
    wire c15396;
    assign in15396_1 = {s14334[0]};
    assign in15396_2 = {c14904};
    Full_Adder FA_15396(s15396, c15396, in15396_1, in15396_2, s14333[0]);
    wire[0:0] s15397, in15397_1, in15397_2;
    wire c15397;
    assign in15397_1 = {s14906[0]};
    assign in15397_2 = {s14907[0]};
    Full_Adder FA_15397(s15397, c15397, in15397_1, in15397_2, c14905);
    wire[0:0] s15398, in15398_1, in15398_2;
    wire c15398;
    assign in15398_1 = {s14338[0]};
    assign in15398_2 = {c14906};
    Full_Adder FA_15398(s15398, c15398, in15398_1, in15398_2, s14337[0]);
    wire[0:0] s15399, in15399_1, in15399_2;
    wire c15399;
    assign in15399_1 = {s14908[0]};
    assign in15399_2 = {s14909[0]};
    Full_Adder FA_15399(s15399, c15399, in15399_1, in15399_2, c14907);
    wire[0:0] s15400, in15400_1, in15400_2;
    wire c15400;
    assign in15400_1 = {s14342[0]};
    assign in15400_2 = {c14908};
    Full_Adder FA_15400(s15400, c15400, in15400_1, in15400_2, s14341[0]);
    wire[0:0] s15401, in15401_1, in15401_2;
    wire c15401;
    assign in15401_1 = {s14910[0]};
    assign in15401_2 = {s14911[0]};
    Full_Adder FA_15401(s15401, c15401, in15401_1, in15401_2, c14909);
    wire[0:0] s15402, in15402_1, in15402_2;
    wire c15402;
    assign in15402_1 = {s14346[0]};
    assign in15402_2 = {c14910};
    Full_Adder FA_15402(s15402, c15402, in15402_1, in15402_2, s14345[0]);
    wire[0:0] s15403, in15403_1, in15403_2;
    wire c15403;
    assign in15403_1 = {s14912[0]};
    assign in15403_2 = {s14913[0]};
    Full_Adder FA_15403(s15403, c15403, in15403_1, in15403_2, c14911);
    wire[0:0] s15404, in15404_1, in15404_2;
    wire c15404;
    assign in15404_1 = {s14350[0]};
    assign in15404_2 = {c14912};
    Full_Adder FA_15404(s15404, c15404, in15404_1, in15404_2, s14349[0]);
    wire[0:0] s15405, in15405_1, in15405_2;
    wire c15405;
    assign in15405_1 = {s14914[0]};
    assign in15405_2 = {s14915[0]};
    Full_Adder FA_15405(s15405, c15405, in15405_1, in15405_2, c14913);
    wire[0:0] s15406, in15406_1, in15406_2;
    wire c15406;
    assign in15406_1 = {s14354[0]};
    assign in15406_2 = {c14914};
    Full_Adder FA_15406(s15406, c15406, in15406_1, in15406_2, s14353[0]);
    wire[0:0] s15407, in15407_1, in15407_2;
    wire c15407;
    assign in15407_1 = {s14916[0]};
    assign in15407_2 = {s14917[0]};
    Full_Adder FA_15407(s15407, c15407, in15407_1, in15407_2, c14915);
    wire[0:0] s15408, in15408_1, in15408_2;
    wire c15408;
    assign in15408_1 = {s14358[0]};
    assign in15408_2 = {c14916};
    Full_Adder FA_15408(s15408, c15408, in15408_1, in15408_2, s14357[0]);
    wire[0:0] s15409, in15409_1, in15409_2;
    wire c15409;
    assign in15409_1 = {s14918[0]};
    assign in15409_2 = {s14919[0]};
    Full_Adder FA_15409(s15409, c15409, in15409_1, in15409_2, c14917);
    wire[0:0] s15410, in15410_1, in15410_2;
    wire c15410;
    assign in15410_1 = {s14362[0]};
    assign in15410_2 = {c14918};
    Full_Adder FA_15410(s15410, c15410, in15410_1, in15410_2, s14361[0]);
    wire[0:0] s15411, in15411_1, in15411_2;
    wire c15411;
    assign in15411_1 = {s14920[0]};
    assign in15411_2 = {s14921[0]};
    Full_Adder FA_15411(s15411, c15411, in15411_1, in15411_2, c14919);
    wire[0:0] s15412, in15412_1, in15412_2;
    wire c15412;
    assign in15412_1 = {s14366[0]};
    assign in15412_2 = {c14920};
    Full_Adder FA_15412(s15412, c15412, in15412_1, in15412_2, s14365[0]);
    wire[0:0] s15413, in15413_1, in15413_2;
    wire c15413;
    assign in15413_1 = {s14922[0]};
    assign in15413_2 = {s14923[0]};
    Full_Adder FA_15413(s15413, c15413, in15413_1, in15413_2, c14921);
    wire[0:0] s15414, in15414_1, in15414_2;
    wire c15414;
    assign in15414_1 = {s14370[0]};
    assign in15414_2 = {c14922};
    Full_Adder FA_15414(s15414, c15414, in15414_1, in15414_2, s14369[0]);
    wire[0:0] s15415, in15415_1, in15415_2;
    wire c15415;
    assign in15415_1 = {s14924[0]};
    assign in15415_2 = {s14925[0]};
    Full_Adder FA_15415(s15415, c15415, in15415_1, in15415_2, c14923);
    wire[0:0] s15416, in15416_1, in15416_2;
    wire c15416;
    assign in15416_1 = {s14374[0]};
    assign in15416_2 = {c14924};
    Full_Adder FA_15416(s15416, c15416, in15416_1, in15416_2, s14373[0]);
    wire[0:0] s15417, in15417_1, in15417_2;
    wire c15417;
    assign in15417_1 = {s14926[0]};
    assign in15417_2 = {s14927[0]};
    Full_Adder FA_15417(s15417, c15417, in15417_1, in15417_2, c14925);
    wire[0:0] s15418, in15418_1, in15418_2;
    wire c15418;
    assign in15418_1 = {s14378[0]};
    assign in15418_2 = {c14926};
    Full_Adder FA_15418(s15418, c15418, in15418_1, in15418_2, s14377[0]);
    wire[0:0] s15419, in15419_1, in15419_2;
    wire c15419;
    assign in15419_1 = {s14928[0]};
    assign in15419_2 = {s14929[0]};
    Full_Adder FA_15419(s15419, c15419, in15419_1, in15419_2, c14927);
    wire[0:0] s15420, in15420_1, in15420_2;
    wire c15420;
    assign in15420_1 = {s14382[0]};
    assign in15420_2 = {c14928};
    Full_Adder FA_15420(s15420, c15420, in15420_1, in15420_2, s14381[0]);
    wire[0:0] s15421, in15421_1, in15421_2;
    wire c15421;
    assign in15421_1 = {s14930[0]};
    assign in15421_2 = {s14931[0]};
    Full_Adder FA_15421(s15421, c15421, in15421_1, in15421_2, c14929);
    wire[0:0] s15422, in15422_1, in15422_2;
    wire c15422;
    assign in15422_1 = {s14386[0]};
    assign in15422_2 = {c14930};
    Full_Adder FA_15422(s15422, c15422, in15422_1, in15422_2, s14385[0]);
    wire[0:0] s15423, in15423_1, in15423_2;
    wire c15423;
    assign in15423_1 = {s14932[0]};
    assign in15423_2 = {s14933[0]};
    Full_Adder FA_15423(s15423, c15423, in15423_1, in15423_2, c14931);
    wire[0:0] s15424, in15424_1, in15424_2;
    wire c15424;
    assign in15424_1 = {s14390[0]};
    assign in15424_2 = {c14932};
    Full_Adder FA_15424(s15424, c15424, in15424_1, in15424_2, s14389[0]);
    wire[0:0] s15425, in15425_1, in15425_2;
    wire c15425;
    assign in15425_1 = {s14934[0]};
    assign in15425_2 = {s14935[0]};
    Full_Adder FA_15425(s15425, c15425, in15425_1, in15425_2, c14933);
    wire[0:0] s15426, in15426_1, in15426_2;
    wire c15426;
    assign in15426_1 = {s14394[0]};
    assign in15426_2 = {c14934};
    Full_Adder FA_15426(s15426, c15426, in15426_1, in15426_2, s14393[0]);
    wire[0:0] s15427, in15427_1, in15427_2;
    wire c15427;
    assign in15427_1 = {s14936[0]};
    assign in15427_2 = {s14937[0]};
    Full_Adder FA_15427(s15427, c15427, in15427_1, in15427_2, c14935);
    wire[0:0] s15428, in15428_1, in15428_2;
    wire c15428;
    assign in15428_1 = {s14398[0]};
    assign in15428_2 = {c14936};
    Full_Adder FA_15428(s15428, c15428, in15428_1, in15428_2, s14397[0]);
    wire[0:0] s15429, in15429_1, in15429_2;
    wire c15429;
    assign in15429_1 = {s14938[0]};
    assign in15429_2 = {s14939[0]};
    Full_Adder FA_15429(s15429, c15429, in15429_1, in15429_2, c14937);
    wire[0:0] s15430, in15430_1, in15430_2;
    wire c15430;
    assign in15430_1 = {s14402[0]};
    assign in15430_2 = {c14938};
    Full_Adder FA_15430(s15430, c15430, in15430_1, in15430_2, s14401[0]);
    wire[0:0] s15431, in15431_1, in15431_2;
    wire c15431;
    assign in15431_1 = {s14940[0]};
    assign in15431_2 = {s14941[0]};
    Full_Adder FA_15431(s15431, c15431, in15431_1, in15431_2, c14939);
    wire[0:0] s15432, in15432_1, in15432_2;
    wire c15432;
    assign in15432_1 = {s14406[0]};
    assign in15432_2 = {c14940};
    Full_Adder FA_15432(s15432, c15432, in15432_1, in15432_2, s14405[0]);
    wire[0:0] s15433, in15433_1, in15433_2;
    wire c15433;
    assign in15433_1 = {s14942[0]};
    assign in15433_2 = {s14943[0]};
    Full_Adder FA_15433(s15433, c15433, in15433_1, in15433_2, c14941);
    wire[0:0] s15434, in15434_1, in15434_2;
    wire c15434;
    assign in15434_1 = {s14410[0]};
    assign in15434_2 = {c14942};
    Full_Adder FA_15434(s15434, c15434, in15434_1, in15434_2, s14409[0]);
    wire[0:0] s15435, in15435_1, in15435_2;
    wire c15435;
    assign in15435_1 = {s14944[0]};
    assign in15435_2 = {s14945[0]};
    Full_Adder FA_15435(s15435, c15435, in15435_1, in15435_2, c14943);
    wire[0:0] s15436, in15436_1, in15436_2;
    wire c15436;
    assign in15436_1 = {s14414[0]};
    assign in15436_2 = {c14944};
    Full_Adder FA_15436(s15436, c15436, in15436_1, in15436_2, s14413[0]);
    wire[0:0] s15437, in15437_1, in15437_2;
    wire c15437;
    assign in15437_1 = {s14946[0]};
    assign in15437_2 = {s14947[0]};
    Full_Adder FA_15437(s15437, c15437, in15437_1, in15437_2, c14945);
    wire[0:0] s15438, in15438_1, in15438_2;
    wire c15438;
    assign in15438_1 = {s14418[0]};
    assign in15438_2 = {c14946};
    Full_Adder FA_15438(s15438, c15438, in15438_1, in15438_2, s14417[0]);
    wire[0:0] s15439, in15439_1, in15439_2;
    wire c15439;
    assign in15439_1 = {s14948[0]};
    assign in15439_2 = {s14949[0]};
    Full_Adder FA_15439(s15439, c15439, in15439_1, in15439_2, c14947);
    wire[0:0] s15440, in15440_1, in15440_2;
    wire c15440;
    assign in15440_1 = {s14422[0]};
    assign in15440_2 = {c14948};
    Full_Adder FA_15440(s15440, c15440, in15440_1, in15440_2, s14421[0]);
    wire[0:0] s15441, in15441_1, in15441_2;
    wire c15441;
    assign in15441_1 = {s14950[0]};
    assign in15441_2 = {s14951[0]};
    Full_Adder FA_15441(s15441, c15441, in15441_1, in15441_2, c14949);
    wire[0:0] s15442, in15442_1, in15442_2;
    wire c15442;
    assign in15442_1 = {s14426[0]};
    assign in15442_2 = {c14950};
    Full_Adder FA_15442(s15442, c15442, in15442_1, in15442_2, s14425[0]);
    wire[0:0] s15443, in15443_1, in15443_2;
    wire c15443;
    assign in15443_1 = {s14952[0]};
    assign in15443_2 = {s14953[0]};
    Full_Adder FA_15443(s15443, c15443, in15443_1, in15443_2, c14951);
    wire[0:0] s15444, in15444_1, in15444_2;
    wire c15444;
    assign in15444_1 = {s14430[0]};
    assign in15444_2 = {c14952};
    Full_Adder FA_15444(s15444, c15444, in15444_1, in15444_2, s14429[0]);
    wire[0:0] s15445, in15445_1, in15445_2;
    wire c15445;
    assign in15445_1 = {s14954[0]};
    assign in15445_2 = {s14955[0]};
    Full_Adder FA_15445(s15445, c15445, in15445_1, in15445_2, c14953);
    wire[0:0] s15446, in15446_1, in15446_2;
    wire c15446;
    assign in15446_1 = {s14434[0]};
    assign in15446_2 = {c14954};
    Full_Adder FA_15446(s15446, c15446, in15446_1, in15446_2, s14433[0]);
    wire[0:0] s15447, in15447_1, in15447_2;
    wire c15447;
    assign in15447_1 = {s14956[0]};
    assign in15447_2 = {s14957[0]};
    Full_Adder FA_15447(s15447, c15447, in15447_1, in15447_2, c14955);
    wire[0:0] s15448, in15448_1, in15448_2;
    wire c15448;
    assign in15448_1 = {s14438[0]};
    assign in15448_2 = {c14956};
    Full_Adder FA_15448(s15448, c15448, in15448_1, in15448_2, s14437[0]);
    wire[0:0] s15449, in15449_1, in15449_2;
    wire c15449;
    assign in15449_1 = {s14958[0]};
    assign in15449_2 = {s14959[0]};
    Full_Adder FA_15449(s15449, c15449, in15449_1, in15449_2, c14957);
    wire[0:0] s15450, in15450_1, in15450_2;
    wire c15450;
    assign in15450_1 = {s14442[0]};
    assign in15450_2 = {c14958};
    Full_Adder FA_15450(s15450, c15450, in15450_1, in15450_2, s14441[0]);
    wire[0:0] s15451, in15451_1, in15451_2;
    wire c15451;
    assign in15451_1 = {s14960[0]};
    assign in15451_2 = {s14961[0]};
    Full_Adder FA_15451(s15451, c15451, in15451_1, in15451_2, c14959);
    wire[0:0] s15452, in15452_1, in15452_2;
    wire c15452;
    assign in15452_1 = {s14446[0]};
    assign in15452_2 = {c14960};
    Full_Adder FA_15452(s15452, c15452, in15452_1, in15452_2, s14445[0]);
    wire[0:0] s15453, in15453_1, in15453_2;
    wire c15453;
    assign in15453_1 = {s14962[0]};
    assign in15453_2 = {s14963[0]};
    Full_Adder FA_15453(s15453, c15453, in15453_1, in15453_2, c14961);
    wire[0:0] s15454, in15454_1, in15454_2;
    wire c15454;
    assign in15454_1 = {s14450[0]};
    assign in15454_2 = {c14962};
    Full_Adder FA_15454(s15454, c15454, in15454_1, in15454_2, s14449[0]);
    wire[0:0] s15455, in15455_1, in15455_2;
    wire c15455;
    assign in15455_1 = {s14964[0]};
    assign in15455_2 = {s14965[0]};
    Full_Adder FA_15455(s15455, c15455, in15455_1, in15455_2, c14963);
    wire[0:0] s15456, in15456_1, in15456_2;
    wire c15456;
    assign in15456_1 = {s14454[0]};
    assign in15456_2 = {c14964};
    Full_Adder FA_15456(s15456, c15456, in15456_1, in15456_2, s14453[0]);
    wire[0:0] s15457, in15457_1, in15457_2;
    wire c15457;
    assign in15457_1 = {s14966[0]};
    assign in15457_2 = {s14967[0]};
    Full_Adder FA_15457(s15457, c15457, in15457_1, in15457_2, c14965);
    wire[0:0] s15458, in15458_1, in15458_2;
    wire c15458;
    assign in15458_1 = {s14458[0]};
    assign in15458_2 = {c14966};
    Full_Adder FA_15458(s15458, c15458, in15458_1, in15458_2, s14457[0]);
    wire[0:0] s15459, in15459_1, in15459_2;
    wire c15459;
    assign in15459_1 = {s14968[0]};
    assign in15459_2 = {s14969[0]};
    Full_Adder FA_15459(s15459, c15459, in15459_1, in15459_2, c14967);
    wire[0:0] s15460, in15460_1, in15460_2;
    wire c15460;
    assign in15460_1 = {s14462[0]};
    assign in15460_2 = {c14968};
    Full_Adder FA_15460(s15460, c15460, in15460_1, in15460_2, s14461[0]);
    wire[0:0] s15461, in15461_1, in15461_2;
    wire c15461;
    assign in15461_1 = {s14970[0]};
    assign in15461_2 = {s14971[0]};
    Full_Adder FA_15461(s15461, c15461, in15461_1, in15461_2, c14969);
    wire[0:0] s15462, in15462_1, in15462_2;
    wire c15462;
    assign in15462_1 = {s14466[0]};
    assign in15462_2 = {c14970};
    Full_Adder FA_15462(s15462, c15462, in15462_1, in15462_2, s14465[0]);
    wire[0:0] s15463, in15463_1, in15463_2;
    wire c15463;
    assign in15463_1 = {s14972[0]};
    assign in15463_2 = {s14973[0]};
    Full_Adder FA_15463(s15463, c15463, in15463_1, in15463_2, c14971);
    wire[0:0] s15464, in15464_1, in15464_2;
    wire c15464;
    assign in15464_1 = {s14470[0]};
    assign in15464_2 = {c14972};
    Full_Adder FA_15464(s15464, c15464, in15464_1, in15464_2, s14469[0]);
    wire[0:0] s15465, in15465_1, in15465_2;
    wire c15465;
    assign in15465_1 = {s14974[0]};
    assign in15465_2 = {s14975[0]};
    Full_Adder FA_15465(s15465, c15465, in15465_1, in15465_2, c14973);
    wire[0:0] s15466, in15466_1, in15466_2;
    wire c15466;
    assign in15466_1 = {s14474[0]};
    assign in15466_2 = {c14974};
    Full_Adder FA_15466(s15466, c15466, in15466_1, in15466_2, s14473[0]);
    wire[0:0] s15467, in15467_1, in15467_2;
    wire c15467;
    assign in15467_1 = {s14976[0]};
    assign in15467_2 = {s14977[0]};
    Full_Adder FA_15467(s15467, c15467, in15467_1, in15467_2, c14975);
    wire[0:0] s15468, in15468_1, in15468_2;
    wire c15468;
    assign in15468_1 = {s14478[0]};
    assign in15468_2 = {c14976};
    Full_Adder FA_15468(s15468, c15468, in15468_1, in15468_2, s14477[0]);
    wire[0:0] s15469, in15469_1, in15469_2;
    wire c15469;
    assign in15469_1 = {s14978[0]};
    assign in15469_2 = {s14979[0]};
    Full_Adder FA_15469(s15469, c15469, in15469_1, in15469_2, c14977);
    wire[0:0] s15470, in15470_1, in15470_2;
    wire c15470;
    assign in15470_1 = {s14482[0]};
    assign in15470_2 = {c14978};
    Full_Adder FA_15470(s15470, c15470, in15470_1, in15470_2, s14481[0]);
    wire[0:0] s15471, in15471_1, in15471_2;
    wire c15471;
    assign in15471_1 = {s14980[0]};
    assign in15471_2 = {s14981[0]};
    Full_Adder FA_15471(s15471, c15471, in15471_1, in15471_2, c14979);
    wire[0:0] s15472, in15472_1, in15472_2;
    wire c15472;
    assign in15472_1 = {s14486[0]};
    assign in15472_2 = {c14980};
    Full_Adder FA_15472(s15472, c15472, in15472_1, in15472_2, s14485[0]);
    wire[0:0] s15473, in15473_1, in15473_2;
    wire c15473;
    assign in15473_1 = {s14982[0]};
    assign in15473_2 = {s14983[0]};
    Full_Adder FA_15473(s15473, c15473, in15473_1, in15473_2, c14981);
    wire[0:0] s15474, in15474_1, in15474_2;
    wire c15474;
    assign in15474_1 = {s14490[0]};
    assign in15474_2 = {c14982};
    Full_Adder FA_15474(s15474, c15474, in15474_1, in15474_2, s14489[0]);
    wire[0:0] s15475, in15475_1, in15475_2;
    wire c15475;
    assign in15475_1 = {s14984[0]};
    assign in15475_2 = {s14985[0]};
    Full_Adder FA_15475(s15475, c15475, in15475_1, in15475_2, c14983);
    wire[0:0] s15476, in15476_1, in15476_2;
    wire c15476;
    assign in15476_1 = {s14494[0]};
    assign in15476_2 = {c14984};
    Full_Adder FA_15476(s15476, c15476, in15476_1, in15476_2, s14493[0]);
    wire[0:0] s15477, in15477_1, in15477_2;
    wire c15477;
    assign in15477_1 = {s14986[0]};
    assign in15477_2 = {s14987[0]};
    Full_Adder FA_15477(s15477, c15477, in15477_1, in15477_2, c14985);
    wire[0:0] s15478, in15478_1, in15478_2;
    wire c15478;
    assign in15478_1 = {s14498[0]};
    assign in15478_2 = {c14986};
    Full_Adder FA_15478(s15478, c15478, in15478_1, in15478_2, s14497[0]);
    wire[0:0] s15479, in15479_1, in15479_2;
    wire c15479;
    assign in15479_1 = {s14988[0]};
    assign in15479_2 = {s14989[0]};
    Full_Adder FA_15479(s15479, c15479, in15479_1, in15479_2, c14987);
    wire[0:0] s15480, in15480_1, in15480_2;
    wire c15480;
    assign in15480_1 = {s14502[0]};
    assign in15480_2 = {c14988};
    Full_Adder FA_15480(s15480, c15480, in15480_1, in15480_2, s14501[0]);
    wire[0:0] s15481, in15481_1, in15481_2;
    wire c15481;
    assign in15481_1 = {s14990[0]};
    assign in15481_2 = {s14991[0]};
    Full_Adder FA_15481(s15481, c15481, in15481_1, in15481_2, c14989);
    wire[0:0] s15482, in15482_1, in15482_2;
    wire c15482;
    assign in15482_1 = {s14506[0]};
    assign in15482_2 = {c14990};
    Full_Adder FA_15482(s15482, c15482, in15482_1, in15482_2, s14505[0]);
    wire[0:0] s15483, in15483_1, in15483_2;
    wire c15483;
    assign in15483_1 = {s14992[0]};
    assign in15483_2 = {s14993[0]};
    Full_Adder FA_15483(s15483, c15483, in15483_1, in15483_2, c14991);
    wire[0:0] s15484, in15484_1, in15484_2;
    wire c15484;
    assign in15484_1 = {s14510[0]};
    assign in15484_2 = {c14992};
    Full_Adder FA_15484(s15484, c15484, in15484_1, in15484_2, s14509[0]);
    wire[0:0] s15485, in15485_1, in15485_2;
    wire c15485;
    assign in15485_1 = {s14994[0]};
    assign in15485_2 = {s14995[0]};
    Full_Adder FA_15485(s15485, c15485, in15485_1, in15485_2, c14993);
    wire[0:0] s15486, in15486_1, in15486_2;
    wire c15486;
    assign in15486_1 = {s14514[0]};
    assign in15486_2 = {c14994};
    Full_Adder FA_15486(s15486, c15486, in15486_1, in15486_2, s14513[0]);
    wire[0:0] s15487, in15487_1, in15487_2;
    wire c15487;
    assign in15487_1 = {s14996[0]};
    assign in15487_2 = {s14997[0]};
    Full_Adder FA_15487(s15487, c15487, in15487_1, in15487_2, c14995);
    wire[0:0] s15488, in15488_1, in15488_2;
    wire c15488;
    assign in15488_1 = {s14517[0]};
    assign in15488_2 = {c14996};
    Full_Adder FA_15488(s15488, c15488, in15488_1, in15488_2, s14516[0]);
    wire[0:0] s15489, in15489_1, in15489_2;
    wire c15489;
    assign in15489_1 = {s14998[0]};
    assign in15489_2 = {s14999[0]};
    Full_Adder FA_15489(s15489, c15489, in15489_1, in15489_2, c14997);
    wire[0:0] s15490, in15490_1, in15490_2;
    wire c15490;
    assign in15490_1 = {s14519[0]};
    assign in15490_2 = {c14998};
    Full_Adder FA_15490(s15490, c15490, in15490_1, in15490_2, s14518[0]);
    wire[0:0] s15491, in15491_1, in15491_2;
    wire c15491;
    assign in15491_1 = {s15000[0]};
    assign in15491_2 = {s15001[0]};
    Full_Adder FA_15491(s15491, c15491, in15491_1, in15491_2, c14999);
    wire[0:0] s15492, in15492_1, in15492_2;
    wire c15492;
    assign in15492_1 = {s14520[0]};
    assign in15492_2 = {c15000};
    Full_Adder FA_15492(s15492, c15492, in15492_1, in15492_2, c14519);
    wire[0:0] s15493, in15493_1, in15493_2;
    wire c15493;
    assign in15493_1 = {s15002[0]};
    assign in15493_2 = {s15003[0]};
    Full_Adder FA_15493(s15493, c15493, in15493_1, in15493_2, c15001);
    wire[0:0] s15494, in15494_1, in15494_2;
    wire c15494;
    assign in15494_1 = {c14520};
    assign in15494_2 = {c15002};
    Full_Adder FA_15494(s15494, c15494, in15494_1, in15494_2, pp127[121]);
    wire[0:0] s15495, in15495_1, in15495_2;
    wire c15495;
    assign in15495_1 = {s15004[0]};
    assign in15495_2 = {s15005[0]};
    Full_Adder FA_15495(s15495, c15495, in15495_1, in15495_2, c15003);
    wire[0:0] s15496, in15496_1, in15496_2;
    wire c15496;
    assign in15496_1 = {pp126[123]};
    assign in15496_2 = {pp127[122]};
    Full_Adder FA_15496(s15496, c15496, in15496_1, in15496_2, pp125[124]);
    wire[0:0] s15497, in15497_1, in15497_2;
    wire c15497;
    assign in15497_1 = {c15005};
    assign in15497_2 = {s15006[0]};
    Full_Adder FA_15497(s15497, c15497, in15497_1, in15497_2, c15004);
    wire[0:0] s15498, in15498_1, in15498_2;
    wire c15498;
    assign in15498_1 = {pp124[126]};
    assign in15498_2 = {pp125[125]};
    Full_Adder FA_15498(s15498, c15498, in15498_1, in15498_2, pp123[127]);
    wire[0:0] s15499, in15499_1, in15499_2;
    wire c15499;
    assign in15499_1 = {pp127[123]};
    assign in15499_2 = {c15006};
    Full_Adder FA_15499(s15499, c15499, in15499_1, in15499_2, pp126[124]);
    wire[0:0] s15500, in15500_1, in15500_2;
    wire c15500;
    assign in15500_1 = {pp125[126]};
    assign in15500_2 = {pp126[125]};
    Full_Adder FA_15500(s15500, c15500, in15500_1, in15500_2, pp124[127]);

    /*Stage 10*/
    wire[0:0] s15501, in15501_1, in15501_2;
    wire c15501;
    assign in15501_1 = {pp0[3]};
    assign in15501_2 = {pp1[2]};
    Half_Adder HA_15501(s15501, c15501, in15501_1, in15501_2);
    wire[0:0] s15502, in15502_1, in15502_2;
    wire c15502;
    assign in15502_1 = {pp3[1]};
    assign in15502_2 = {pp4[0]};
    Full_Adder FA_15502(s15502, c15502, in15502_1, in15502_2, pp2[2]);
    wire[0:0] s15503, in15503_1, in15503_2;
    wire c15503;
    assign in15503_1 = {c15007};
    assign in15503_2 = {s15008[0]};
    Full_Adder FA_15503(s15503, c15503, in15503_1, in15503_2, pp5[0]);
    wire[0:0] s15504, in15504_1, in15504_2;
    wire c15504;
    assign in15504_1 = {c15009};
    assign in15504_2 = {s15010[0]};
    Full_Adder FA_15504(s15504, c15504, in15504_1, in15504_2, c15008);
    wire[0:0] s15505, in15505_1, in15505_2;
    wire c15505;
    assign in15505_1 = {c15011};
    assign in15505_2 = {s15012[0]};
    Full_Adder FA_15505(s15505, c15505, in15505_1, in15505_2, c15010);
    wire[0:0] s15506, in15506_1, in15506_2;
    wire c15506;
    assign in15506_1 = {c15013};
    assign in15506_2 = {s15014[0]};
    Full_Adder FA_15506(s15506, c15506, in15506_1, in15506_2, c15012);
    wire[0:0] s15507, in15507_1, in15507_2;
    wire c15507;
    assign in15507_1 = {c15015};
    assign in15507_2 = {s15016[0]};
    Full_Adder FA_15507(s15507, c15507, in15507_1, in15507_2, c15014);
    wire[0:0] s15508, in15508_1, in15508_2;
    wire c15508;
    assign in15508_1 = {c15017};
    assign in15508_2 = {s15018[0]};
    Full_Adder FA_15508(s15508, c15508, in15508_1, in15508_2, c15016);
    wire[0:0] s15509, in15509_1, in15509_2;
    wire c15509;
    assign in15509_1 = {c15019};
    assign in15509_2 = {s15020[0]};
    Full_Adder FA_15509(s15509, c15509, in15509_1, in15509_2, c15018);
    wire[0:0] s15510, in15510_1, in15510_2;
    wire c15510;
    assign in15510_1 = {c15021};
    assign in15510_2 = {s15022[0]};
    Full_Adder FA_15510(s15510, c15510, in15510_1, in15510_2, c15020);
    wire[0:0] s15511, in15511_1, in15511_2;
    wire c15511;
    assign in15511_1 = {c15023};
    assign in15511_2 = {s15024[0]};
    Full_Adder FA_15511(s15511, c15511, in15511_1, in15511_2, c15022);
    wire[0:0] s15512, in15512_1, in15512_2;
    wire c15512;
    assign in15512_1 = {c15025};
    assign in15512_2 = {s15026[0]};
    Full_Adder FA_15512(s15512, c15512, in15512_1, in15512_2, c15024);
    wire[0:0] s15513, in15513_1, in15513_2;
    wire c15513;
    assign in15513_1 = {c15027};
    assign in15513_2 = {s15028[0]};
    Full_Adder FA_15513(s15513, c15513, in15513_1, in15513_2, c15026);
    wire[0:0] s15514, in15514_1, in15514_2;
    wire c15514;
    assign in15514_1 = {c15029};
    assign in15514_2 = {s15030[0]};
    Full_Adder FA_15514(s15514, c15514, in15514_1, in15514_2, c15028);
    wire[0:0] s15515, in15515_1, in15515_2;
    wire c15515;
    assign in15515_1 = {c15031};
    assign in15515_2 = {s15032[0]};
    Full_Adder FA_15515(s15515, c15515, in15515_1, in15515_2, c15030);
    wire[0:0] s15516, in15516_1, in15516_2;
    wire c15516;
    assign in15516_1 = {c15033};
    assign in15516_2 = {s15034[0]};
    Full_Adder FA_15516(s15516, c15516, in15516_1, in15516_2, c15032);
    wire[0:0] s15517, in15517_1, in15517_2;
    wire c15517;
    assign in15517_1 = {c15035};
    assign in15517_2 = {s15036[0]};
    Full_Adder FA_15517(s15517, c15517, in15517_1, in15517_2, c15034);
    wire[0:0] s15518, in15518_1, in15518_2;
    wire c15518;
    assign in15518_1 = {c15037};
    assign in15518_2 = {s15038[0]};
    Full_Adder FA_15518(s15518, c15518, in15518_1, in15518_2, c15036);
    wire[0:0] s15519, in15519_1, in15519_2;
    wire c15519;
    assign in15519_1 = {c15039};
    assign in15519_2 = {s15040[0]};
    Full_Adder FA_15519(s15519, c15519, in15519_1, in15519_2, c15038);
    wire[0:0] s15520, in15520_1, in15520_2;
    wire c15520;
    assign in15520_1 = {c15041};
    assign in15520_2 = {s15042[0]};
    Full_Adder FA_15520(s15520, c15520, in15520_1, in15520_2, c15040);
    wire[0:0] s15521, in15521_1, in15521_2;
    wire c15521;
    assign in15521_1 = {c15043};
    assign in15521_2 = {s15044[0]};
    Full_Adder FA_15521(s15521, c15521, in15521_1, in15521_2, c15042);
    wire[0:0] s15522, in15522_1, in15522_2;
    wire c15522;
    assign in15522_1 = {c15045};
    assign in15522_2 = {s15046[0]};
    Full_Adder FA_15522(s15522, c15522, in15522_1, in15522_2, c15044);
    wire[0:0] s15523, in15523_1, in15523_2;
    wire c15523;
    assign in15523_1 = {c15047};
    assign in15523_2 = {s15048[0]};
    Full_Adder FA_15523(s15523, c15523, in15523_1, in15523_2, c15046);
    wire[0:0] s15524, in15524_1, in15524_2;
    wire c15524;
    assign in15524_1 = {c15049};
    assign in15524_2 = {s15050[0]};
    Full_Adder FA_15524(s15524, c15524, in15524_1, in15524_2, c15048);
    wire[0:0] s15525, in15525_1, in15525_2;
    wire c15525;
    assign in15525_1 = {c15051};
    assign in15525_2 = {s15052[0]};
    Full_Adder FA_15525(s15525, c15525, in15525_1, in15525_2, c15050);
    wire[0:0] s15526, in15526_1, in15526_2;
    wire c15526;
    assign in15526_1 = {c15053};
    assign in15526_2 = {s15054[0]};
    Full_Adder FA_15526(s15526, c15526, in15526_1, in15526_2, c15052);
    wire[0:0] s15527, in15527_1, in15527_2;
    wire c15527;
    assign in15527_1 = {c15055};
    assign in15527_2 = {s15056[0]};
    Full_Adder FA_15527(s15527, c15527, in15527_1, in15527_2, c15054);
    wire[0:0] s15528, in15528_1, in15528_2;
    wire c15528;
    assign in15528_1 = {c15057};
    assign in15528_2 = {s15058[0]};
    Full_Adder FA_15528(s15528, c15528, in15528_1, in15528_2, c15056);
    wire[0:0] s15529, in15529_1, in15529_2;
    wire c15529;
    assign in15529_1 = {c15059};
    assign in15529_2 = {s15060[0]};
    Full_Adder FA_15529(s15529, c15529, in15529_1, in15529_2, c15058);
    wire[0:0] s15530, in15530_1, in15530_2;
    wire c15530;
    assign in15530_1 = {c15061};
    assign in15530_2 = {s15062[0]};
    Full_Adder FA_15530(s15530, c15530, in15530_1, in15530_2, c15060);
    wire[0:0] s15531, in15531_1, in15531_2;
    wire c15531;
    assign in15531_1 = {c15063};
    assign in15531_2 = {s15064[0]};
    Full_Adder FA_15531(s15531, c15531, in15531_1, in15531_2, c15062);
    wire[0:0] s15532, in15532_1, in15532_2;
    wire c15532;
    assign in15532_1 = {c15065};
    assign in15532_2 = {s15066[0]};
    Full_Adder FA_15532(s15532, c15532, in15532_1, in15532_2, c15064);
    wire[0:0] s15533, in15533_1, in15533_2;
    wire c15533;
    assign in15533_1 = {c15067};
    assign in15533_2 = {s15068[0]};
    Full_Adder FA_15533(s15533, c15533, in15533_1, in15533_2, c15066);
    wire[0:0] s15534, in15534_1, in15534_2;
    wire c15534;
    assign in15534_1 = {c15069};
    assign in15534_2 = {s15070[0]};
    Full_Adder FA_15534(s15534, c15534, in15534_1, in15534_2, c15068);
    wire[0:0] s15535, in15535_1, in15535_2;
    wire c15535;
    assign in15535_1 = {c15071};
    assign in15535_2 = {s15072[0]};
    Full_Adder FA_15535(s15535, c15535, in15535_1, in15535_2, c15070);
    wire[0:0] s15536, in15536_1, in15536_2;
    wire c15536;
    assign in15536_1 = {c15073};
    assign in15536_2 = {s15074[0]};
    Full_Adder FA_15536(s15536, c15536, in15536_1, in15536_2, c15072);
    wire[0:0] s15537, in15537_1, in15537_2;
    wire c15537;
    assign in15537_1 = {c15075};
    assign in15537_2 = {s15076[0]};
    Full_Adder FA_15537(s15537, c15537, in15537_1, in15537_2, c15074);
    wire[0:0] s15538, in15538_1, in15538_2;
    wire c15538;
    assign in15538_1 = {c15077};
    assign in15538_2 = {s15078[0]};
    Full_Adder FA_15538(s15538, c15538, in15538_1, in15538_2, c15076);
    wire[0:0] s15539, in15539_1, in15539_2;
    wire c15539;
    assign in15539_1 = {c15079};
    assign in15539_2 = {s15080[0]};
    Full_Adder FA_15539(s15539, c15539, in15539_1, in15539_2, c15078);
    wire[0:0] s15540, in15540_1, in15540_2;
    wire c15540;
    assign in15540_1 = {c15081};
    assign in15540_2 = {s15082[0]};
    Full_Adder FA_15540(s15540, c15540, in15540_1, in15540_2, c15080);
    wire[0:0] s15541, in15541_1, in15541_2;
    wire c15541;
    assign in15541_1 = {c15083};
    assign in15541_2 = {s15084[0]};
    Full_Adder FA_15541(s15541, c15541, in15541_1, in15541_2, c15082);
    wire[0:0] s15542, in15542_1, in15542_2;
    wire c15542;
    assign in15542_1 = {c15085};
    assign in15542_2 = {s15086[0]};
    Full_Adder FA_15542(s15542, c15542, in15542_1, in15542_2, c15084);
    wire[0:0] s15543, in15543_1, in15543_2;
    wire c15543;
    assign in15543_1 = {c15087};
    assign in15543_2 = {s15088[0]};
    Full_Adder FA_15543(s15543, c15543, in15543_1, in15543_2, c15086);
    wire[0:0] s15544, in15544_1, in15544_2;
    wire c15544;
    assign in15544_1 = {c15089};
    assign in15544_2 = {s15090[0]};
    Full_Adder FA_15544(s15544, c15544, in15544_1, in15544_2, c15088);
    wire[0:0] s15545, in15545_1, in15545_2;
    wire c15545;
    assign in15545_1 = {c15091};
    assign in15545_2 = {s15092[0]};
    Full_Adder FA_15545(s15545, c15545, in15545_1, in15545_2, c15090);
    wire[0:0] s15546, in15546_1, in15546_2;
    wire c15546;
    assign in15546_1 = {c15093};
    assign in15546_2 = {s15094[0]};
    Full_Adder FA_15546(s15546, c15546, in15546_1, in15546_2, c15092);
    wire[0:0] s15547, in15547_1, in15547_2;
    wire c15547;
    assign in15547_1 = {c15095};
    assign in15547_2 = {s15096[0]};
    Full_Adder FA_15547(s15547, c15547, in15547_1, in15547_2, c15094);
    wire[0:0] s15548, in15548_1, in15548_2;
    wire c15548;
    assign in15548_1 = {c15097};
    assign in15548_2 = {s15098[0]};
    Full_Adder FA_15548(s15548, c15548, in15548_1, in15548_2, c15096);
    wire[0:0] s15549, in15549_1, in15549_2;
    wire c15549;
    assign in15549_1 = {c15099};
    assign in15549_2 = {s15100[0]};
    Full_Adder FA_15549(s15549, c15549, in15549_1, in15549_2, c15098);
    wire[0:0] s15550, in15550_1, in15550_2;
    wire c15550;
    assign in15550_1 = {c15101};
    assign in15550_2 = {s15102[0]};
    Full_Adder FA_15550(s15550, c15550, in15550_1, in15550_2, c15100);
    wire[0:0] s15551, in15551_1, in15551_2;
    wire c15551;
    assign in15551_1 = {c15103};
    assign in15551_2 = {s15104[0]};
    Full_Adder FA_15551(s15551, c15551, in15551_1, in15551_2, c15102);
    wire[0:0] s15552, in15552_1, in15552_2;
    wire c15552;
    assign in15552_1 = {c15105};
    assign in15552_2 = {s15106[0]};
    Full_Adder FA_15552(s15552, c15552, in15552_1, in15552_2, c15104);
    wire[0:0] s15553, in15553_1, in15553_2;
    wire c15553;
    assign in15553_1 = {c15107};
    assign in15553_2 = {s15108[0]};
    Full_Adder FA_15553(s15553, c15553, in15553_1, in15553_2, c15106);
    wire[0:0] s15554, in15554_1, in15554_2;
    wire c15554;
    assign in15554_1 = {c15109};
    assign in15554_2 = {s15110[0]};
    Full_Adder FA_15554(s15554, c15554, in15554_1, in15554_2, c15108);
    wire[0:0] s15555, in15555_1, in15555_2;
    wire c15555;
    assign in15555_1 = {c15111};
    assign in15555_2 = {s15112[0]};
    Full_Adder FA_15555(s15555, c15555, in15555_1, in15555_2, c15110);
    wire[0:0] s15556, in15556_1, in15556_2;
    wire c15556;
    assign in15556_1 = {c15113};
    assign in15556_2 = {s15114[0]};
    Full_Adder FA_15556(s15556, c15556, in15556_1, in15556_2, c15112);
    wire[0:0] s15557, in15557_1, in15557_2;
    wire c15557;
    assign in15557_1 = {c15115};
    assign in15557_2 = {s15116[0]};
    Full_Adder FA_15557(s15557, c15557, in15557_1, in15557_2, c15114);
    wire[0:0] s15558, in15558_1, in15558_2;
    wire c15558;
    assign in15558_1 = {c15117};
    assign in15558_2 = {s15118[0]};
    Full_Adder FA_15558(s15558, c15558, in15558_1, in15558_2, c15116);
    wire[0:0] s15559, in15559_1, in15559_2;
    wire c15559;
    assign in15559_1 = {c15119};
    assign in15559_2 = {s15120[0]};
    Full_Adder FA_15559(s15559, c15559, in15559_1, in15559_2, c15118);
    wire[0:0] s15560, in15560_1, in15560_2;
    wire c15560;
    assign in15560_1 = {c15121};
    assign in15560_2 = {s15122[0]};
    Full_Adder FA_15560(s15560, c15560, in15560_1, in15560_2, c15120);
    wire[0:0] s15561, in15561_1, in15561_2;
    wire c15561;
    assign in15561_1 = {c15123};
    assign in15561_2 = {s15124[0]};
    Full_Adder FA_15561(s15561, c15561, in15561_1, in15561_2, c15122);
    wire[0:0] s15562, in15562_1, in15562_2;
    wire c15562;
    assign in15562_1 = {c15125};
    assign in15562_2 = {s15126[0]};
    Full_Adder FA_15562(s15562, c15562, in15562_1, in15562_2, c15124);
    wire[0:0] s15563, in15563_1, in15563_2;
    wire c15563;
    assign in15563_1 = {c15127};
    assign in15563_2 = {s15128[0]};
    Full_Adder FA_15563(s15563, c15563, in15563_1, in15563_2, c15126);
    wire[0:0] s15564, in15564_1, in15564_2;
    wire c15564;
    assign in15564_1 = {c15129};
    assign in15564_2 = {s15130[0]};
    Full_Adder FA_15564(s15564, c15564, in15564_1, in15564_2, c15128);
    wire[0:0] s15565, in15565_1, in15565_2;
    wire c15565;
    assign in15565_1 = {c15131};
    assign in15565_2 = {s15132[0]};
    Full_Adder FA_15565(s15565, c15565, in15565_1, in15565_2, c15130);
    wire[0:0] s15566, in15566_1, in15566_2;
    wire c15566;
    assign in15566_1 = {c15133};
    assign in15566_2 = {s15134[0]};
    Full_Adder FA_15566(s15566, c15566, in15566_1, in15566_2, c15132);
    wire[0:0] s15567, in15567_1, in15567_2;
    wire c15567;
    assign in15567_1 = {c15135};
    assign in15567_2 = {s15136[0]};
    Full_Adder FA_15567(s15567, c15567, in15567_1, in15567_2, c15134);
    wire[0:0] s15568, in15568_1, in15568_2;
    wire c15568;
    assign in15568_1 = {c15137};
    assign in15568_2 = {s15138[0]};
    Full_Adder FA_15568(s15568, c15568, in15568_1, in15568_2, c15136);
    wire[0:0] s15569, in15569_1, in15569_2;
    wire c15569;
    assign in15569_1 = {c15139};
    assign in15569_2 = {s15140[0]};
    Full_Adder FA_15569(s15569, c15569, in15569_1, in15569_2, c15138);
    wire[0:0] s15570, in15570_1, in15570_2;
    wire c15570;
    assign in15570_1 = {c15141};
    assign in15570_2 = {s15142[0]};
    Full_Adder FA_15570(s15570, c15570, in15570_1, in15570_2, c15140);
    wire[0:0] s15571, in15571_1, in15571_2;
    wire c15571;
    assign in15571_1 = {c15143};
    assign in15571_2 = {s15144[0]};
    Full_Adder FA_15571(s15571, c15571, in15571_1, in15571_2, c15142);
    wire[0:0] s15572, in15572_1, in15572_2;
    wire c15572;
    assign in15572_1 = {c15145};
    assign in15572_2 = {s15146[0]};
    Full_Adder FA_15572(s15572, c15572, in15572_1, in15572_2, c15144);
    wire[0:0] s15573, in15573_1, in15573_2;
    wire c15573;
    assign in15573_1 = {c15147};
    assign in15573_2 = {s15148[0]};
    Full_Adder FA_15573(s15573, c15573, in15573_1, in15573_2, c15146);
    wire[0:0] s15574, in15574_1, in15574_2;
    wire c15574;
    assign in15574_1 = {c15149};
    assign in15574_2 = {s15150[0]};
    Full_Adder FA_15574(s15574, c15574, in15574_1, in15574_2, c15148);
    wire[0:0] s15575, in15575_1, in15575_2;
    wire c15575;
    assign in15575_1 = {c15151};
    assign in15575_2 = {s15152[0]};
    Full_Adder FA_15575(s15575, c15575, in15575_1, in15575_2, c15150);
    wire[0:0] s15576, in15576_1, in15576_2;
    wire c15576;
    assign in15576_1 = {c15153};
    assign in15576_2 = {s15154[0]};
    Full_Adder FA_15576(s15576, c15576, in15576_1, in15576_2, c15152);
    wire[0:0] s15577, in15577_1, in15577_2;
    wire c15577;
    assign in15577_1 = {c15155};
    assign in15577_2 = {s15156[0]};
    Full_Adder FA_15577(s15577, c15577, in15577_1, in15577_2, c15154);
    wire[0:0] s15578, in15578_1, in15578_2;
    wire c15578;
    assign in15578_1 = {c15157};
    assign in15578_2 = {s15158[0]};
    Full_Adder FA_15578(s15578, c15578, in15578_1, in15578_2, c15156);
    wire[0:0] s15579, in15579_1, in15579_2;
    wire c15579;
    assign in15579_1 = {c15159};
    assign in15579_2 = {s15160[0]};
    Full_Adder FA_15579(s15579, c15579, in15579_1, in15579_2, c15158);
    wire[0:0] s15580, in15580_1, in15580_2;
    wire c15580;
    assign in15580_1 = {c15161};
    assign in15580_2 = {s15162[0]};
    Full_Adder FA_15580(s15580, c15580, in15580_1, in15580_2, c15160);
    wire[0:0] s15581, in15581_1, in15581_2;
    wire c15581;
    assign in15581_1 = {c15163};
    assign in15581_2 = {s15164[0]};
    Full_Adder FA_15581(s15581, c15581, in15581_1, in15581_2, c15162);
    wire[0:0] s15582, in15582_1, in15582_2;
    wire c15582;
    assign in15582_1 = {c15165};
    assign in15582_2 = {s15166[0]};
    Full_Adder FA_15582(s15582, c15582, in15582_1, in15582_2, c15164);
    wire[0:0] s15583, in15583_1, in15583_2;
    wire c15583;
    assign in15583_1 = {c15167};
    assign in15583_2 = {s15168[0]};
    Full_Adder FA_15583(s15583, c15583, in15583_1, in15583_2, c15166);
    wire[0:0] s15584, in15584_1, in15584_2;
    wire c15584;
    assign in15584_1 = {c15169};
    assign in15584_2 = {s15170[0]};
    Full_Adder FA_15584(s15584, c15584, in15584_1, in15584_2, c15168);
    wire[0:0] s15585, in15585_1, in15585_2;
    wire c15585;
    assign in15585_1 = {c15171};
    assign in15585_2 = {s15172[0]};
    Full_Adder FA_15585(s15585, c15585, in15585_1, in15585_2, c15170);
    wire[0:0] s15586, in15586_1, in15586_2;
    wire c15586;
    assign in15586_1 = {c15173};
    assign in15586_2 = {s15174[0]};
    Full_Adder FA_15586(s15586, c15586, in15586_1, in15586_2, c15172);
    wire[0:0] s15587, in15587_1, in15587_2;
    wire c15587;
    assign in15587_1 = {c15175};
    assign in15587_2 = {s15176[0]};
    Full_Adder FA_15587(s15587, c15587, in15587_1, in15587_2, c15174);
    wire[0:0] s15588, in15588_1, in15588_2;
    wire c15588;
    assign in15588_1 = {c15177};
    assign in15588_2 = {s15178[0]};
    Full_Adder FA_15588(s15588, c15588, in15588_1, in15588_2, c15176);
    wire[0:0] s15589, in15589_1, in15589_2;
    wire c15589;
    assign in15589_1 = {c15179};
    assign in15589_2 = {s15180[0]};
    Full_Adder FA_15589(s15589, c15589, in15589_1, in15589_2, c15178);
    wire[0:0] s15590, in15590_1, in15590_2;
    wire c15590;
    assign in15590_1 = {c15181};
    assign in15590_2 = {s15182[0]};
    Full_Adder FA_15590(s15590, c15590, in15590_1, in15590_2, c15180);
    wire[0:0] s15591, in15591_1, in15591_2;
    wire c15591;
    assign in15591_1 = {c15183};
    assign in15591_2 = {s15184[0]};
    Full_Adder FA_15591(s15591, c15591, in15591_1, in15591_2, c15182);
    wire[0:0] s15592, in15592_1, in15592_2;
    wire c15592;
    assign in15592_1 = {c15185};
    assign in15592_2 = {s15186[0]};
    Full_Adder FA_15592(s15592, c15592, in15592_1, in15592_2, c15184);
    wire[0:0] s15593, in15593_1, in15593_2;
    wire c15593;
    assign in15593_1 = {c15187};
    assign in15593_2 = {s15188[0]};
    Full_Adder FA_15593(s15593, c15593, in15593_1, in15593_2, c15186);
    wire[0:0] s15594, in15594_1, in15594_2;
    wire c15594;
    assign in15594_1 = {c15189};
    assign in15594_2 = {s15190[0]};
    Full_Adder FA_15594(s15594, c15594, in15594_1, in15594_2, c15188);
    wire[0:0] s15595, in15595_1, in15595_2;
    wire c15595;
    assign in15595_1 = {c15191};
    assign in15595_2 = {s15192[0]};
    Full_Adder FA_15595(s15595, c15595, in15595_1, in15595_2, c15190);
    wire[0:0] s15596, in15596_1, in15596_2;
    wire c15596;
    assign in15596_1 = {c15193};
    assign in15596_2 = {s15194[0]};
    Full_Adder FA_15596(s15596, c15596, in15596_1, in15596_2, c15192);
    wire[0:0] s15597, in15597_1, in15597_2;
    wire c15597;
    assign in15597_1 = {c15195};
    assign in15597_2 = {s15196[0]};
    Full_Adder FA_15597(s15597, c15597, in15597_1, in15597_2, c15194);
    wire[0:0] s15598, in15598_1, in15598_2;
    wire c15598;
    assign in15598_1 = {c15197};
    assign in15598_2 = {s15198[0]};
    Full_Adder FA_15598(s15598, c15598, in15598_1, in15598_2, c15196);
    wire[0:0] s15599, in15599_1, in15599_2;
    wire c15599;
    assign in15599_1 = {c15199};
    assign in15599_2 = {s15200[0]};
    Full_Adder FA_15599(s15599, c15599, in15599_1, in15599_2, c15198);
    wire[0:0] s15600, in15600_1, in15600_2;
    wire c15600;
    assign in15600_1 = {c15201};
    assign in15600_2 = {s15202[0]};
    Full_Adder FA_15600(s15600, c15600, in15600_1, in15600_2, c15200);
    wire[0:0] s15601, in15601_1, in15601_2;
    wire c15601;
    assign in15601_1 = {c15203};
    assign in15601_2 = {s15204[0]};
    Full_Adder FA_15601(s15601, c15601, in15601_1, in15601_2, c15202);
    wire[0:0] s15602, in15602_1, in15602_2;
    wire c15602;
    assign in15602_1 = {c15205};
    assign in15602_2 = {s15206[0]};
    Full_Adder FA_15602(s15602, c15602, in15602_1, in15602_2, c15204);
    wire[0:0] s15603, in15603_1, in15603_2;
    wire c15603;
    assign in15603_1 = {c15207};
    assign in15603_2 = {s15208[0]};
    Full_Adder FA_15603(s15603, c15603, in15603_1, in15603_2, c15206);
    wire[0:0] s15604, in15604_1, in15604_2;
    wire c15604;
    assign in15604_1 = {c15209};
    assign in15604_2 = {s15210[0]};
    Full_Adder FA_15604(s15604, c15604, in15604_1, in15604_2, c15208);
    wire[0:0] s15605, in15605_1, in15605_2;
    wire c15605;
    assign in15605_1 = {c15211};
    assign in15605_2 = {s15212[0]};
    Full_Adder FA_15605(s15605, c15605, in15605_1, in15605_2, c15210);
    wire[0:0] s15606, in15606_1, in15606_2;
    wire c15606;
    assign in15606_1 = {c15213};
    assign in15606_2 = {s15214[0]};
    Full_Adder FA_15606(s15606, c15606, in15606_1, in15606_2, c15212);
    wire[0:0] s15607, in15607_1, in15607_2;
    wire c15607;
    assign in15607_1 = {c15215};
    assign in15607_2 = {s15216[0]};
    Full_Adder FA_15607(s15607, c15607, in15607_1, in15607_2, c15214);
    wire[0:0] s15608, in15608_1, in15608_2;
    wire c15608;
    assign in15608_1 = {c15217};
    assign in15608_2 = {s15218[0]};
    Full_Adder FA_15608(s15608, c15608, in15608_1, in15608_2, c15216);
    wire[0:0] s15609, in15609_1, in15609_2;
    wire c15609;
    assign in15609_1 = {c15219};
    assign in15609_2 = {s15220[0]};
    Full_Adder FA_15609(s15609, c15609, in15609_1, in15609_2, c15218);
    wire[0:0] s15610, in15610_1, in15610_2;
    wire c15610;
    assign in15610_1 = {c15221};
    assign in15610_2 = {s15222[0]};
    Full_Adder FA_15610(s15610, c15610, in15610_1, in15610_2, c15220);
    wire[0:0] s15611, in15611_1, in15611_2;
    wire c15611;
    assign in15611_1 = {c15223};
    assign in15611_2 = {s15224[0]};
    Full_Adder FA_15611(s15611, c15611, in15611_1, in15611_2, c15222);
    wire[0:0] s15612, in15612_1, in15612_2;
    wire c15612;
    assign in15612_1 = {c15225};
    assign in15612_2 = {s15226[0]};
    Full_Adder FA_15612(s15612, c15612, in15612_1, in15612_2, c15224);
    wire[0:0] s15613, in15613_1, in15613_2;
    wire c15613;
    assign in15613_1 = {c15227};
    assign in15613_2 = {s15228[0]};
    Full_Adder FA_15613(s15613, c15613, in15613_1, in15613_2, c15226);
    wire[0:0] s15614, in15614_1, in15614_2;
    wire c15614;
    assign in15614_1 = {c15229};
    assign in15614_2 = {s15230[0]};
    Full_Adder FA_15614(s15614, c15614, in15614_1, in15614_2, c15228);
    wire[0:0] s15615, in15615_1, in15615_2;
    wire c15615;
    assign in15615_1 = {c15231};
    assign in15615_2 = {s15232[0]};
    Full_Adder FA_15615(s15615, c15615, in15615_1, in15615_2, c15230);
    wire[0:0] s15616, in15616_1, in15616_2;
    wire c15616;
    assign in15616_1 = {c15233};
    assign in15616_2 = {s15234[0]};
    Full_Adder FA_15616(s15616, c15616, in15616_1, in15616_2, c15232);
    wire[0:0] s15617, in15617_1, in15617_2;
    wire c15617;
    assign in15617_1 = {c15235};
    assign in15617_2 = {s15236[0]};
    Full_Adder FA_15617(s15617, c15617, in15617_1, in15617_2, c15234);
    wire[0:0] s15618, in15618_1, in15618_2;
    wire c15618;
    assign in15618_1 = {c15237};
    assign in15618_2 = {s15238[0]};
    Full_Adder FA_15618(s15618, c15618, in15618_1, in15618_2, c15236);
    wire[0:0] s15619, in15619_1, in15619_2;
    wire c15619;
    assign in15619_1 = {c15239};
    assign in15619_2 = {s15240[0]};
    Full_Adder FA_15619(s15619, c15619, in15619_1, in15619_2, c15238);
    wire[0:0] s15620, in15620_1, in15620_2;
    wire c15620;
    assign in15620_1 = {c15241};
    assign in15620_2 = {s15242[0]};
    Full_Adder FA_15620(s15620, c15620, in15620_1, in15620_2, c15240);
    wire[0:0] s15621, in15621_1, in15621_2;
    wire c15621;
    assign in15621_1 = {c15243};
    assign in15621_2 = {s15244[0]};
    Full_Adder FA_15621(s15621, c15621, in15621_1, in15621_2, c15242);
    wire[0:0] s15622, in15622_1, in15622_2;
    wire c15622;
    assign in15622_1 = {c15245};
    assign in15622_2 = {s15246[0]};
    Full_Adder FA_15622(s15622, c15622, in15622_1, in15622_2, c15244);
    wire[0:0] s15623, in15623_1, in15623_2;
    wire c15623;
    assign in15623_1 = {c15247};
    assign in15623_2 = {s15248[0]};
    Full_Adder FA_15623(s15623, c15623, in15623_1, in15623_2, c15246);
    wire[0:0] s15624, in15624_1, in15624_2;
    wire c15624;
    assign in15624_1 = {c15249};
    assign in15624_2 = {s15250[0]};
    Full_Adder FA_15624(s15624, c15624, in15624_1, in15624_2, c15248);
    wire[0:0] s15625, in15625_1, in15625_2;
    wire c15625;
    assign in15625_1 = {c15251};
    assign in15625_2 = {s15252[0]};
    Full_Adder FA_15625(s15625, c15625, in15625_1, in15625_2, c15250);
    wire[0:0] s15626, in15626_1, in15626_2;
    wire c15626;
    assign in15626_1 = {c15253};
    assign in15626_2 = {s15254[0]};
    Full_Adder FA_15626(s15626, c15626, in15626_1, in15626_2, c15252);
    wire[0:0] s15627, in15627_1, in15627_2;
    wire c15627;
    assign in15627_1 = {c15255};
    assign in15627_2 = {s15256[0]};
    Full_Adder FA_15627(s15627, c15627, in15627_1, in15627_2, c15254);
    wire[0:0] s15628, in15628_1, in15628_2;
    wire c15628;
    assign in15628_1 = {c15257};
    assign in15628_2 = {s15258[0]};
    Full_Adder FA_15628(s15628, c15628, in15628_1, in15628_2, c15256);
    wire[0:0] s15629, in15629_1, in15629_2;
    wire c15629;
    assign in15629_1 = {c15259};
    assign in15629_2 = {s15260[0]};
    Full_Adder FA_15629(s15629, c15629, in15629_1, in15629_2, c15258);
    wire[0:0] s15630, in15630_1, in15630_2;
    wire c15630;
    assign in15630_1 = {c15261};
    assign in15630_2 = {s15262[0]};
    Full_Adder FA_15630(s15630, c15630, in15630_1, in15630_2, c15260);
    wire[0:0] s15631, in15631_1, in15631_2;
    wire c15631;
    assign in15631_1 = {c15263};
    assign in15631_2 = {s15264[0]};
    Full_Adder FA_15631(s15631, c15631, in15631_1, in15631_2, c15262);
    wire[0:0] s15632, in15632_1, in15632_2;
    wire c15632;
    assign in15632_1 = {c15265};
    assign in15632_2 = {s15266[0]};
    Full_Adder FA_15632(s15632, c15632, in15632_1, in15632_2, c15264);
    wire[0:0] s15633, in15633_1, in15633_2;
    wire c15633;
    assign in15633_1 = {c15267};
    assign in15633_2 = {s15268[0]};
    Full_Adder FA_15633(s15633, c15633, in15633_1, in15633_2, c15266);
    wire[0:0] s15634, in15634_1, in15634_2;
    wire c15634;
    assign in15634_1 = {c15269};
    assign in15634_2 = {s15270[0]};
    Full_Adder FA_15634(s15634, c15634, in15634_1, in15634_2, c15268);
    wire[0:0] s15635, in15635_1, in15635_2;
    wire c15635;
    assign in15635_1 = {c15271};
    assign in15635_2 = {s15272[0]};
    Full_Adder FA_15635(s15635, c15635, in15635_1, in15635_2, c15270);
    wire[0:0] s15636, in15636_1, in15636_2;
    wire c15636;
    assign in15636_1 = {c15273};
    assign in15636_2 = {s15274[0]};
    Full_Adder FA_15636(s15636, c15636, in15636_1, in15636_2, c15272);
    wire[0:0] s15637, in15637_1, in15637_2;
    wire c15637;
    assign in15637_1 = {c15275};
    assign in15637_2 = {s15276[0]};
    Full_Adder FA_15637(s15637, c15637, in15637_1, in15637_2, c15274);
    wire[0:0] s15638, in15638_1, in15638_2;
    wire c15638;
    assign in15638_1 = {c15277};
    assign in15638_2 = {s15278[0]};
    Full_Adder FA_15638(s15638, c15638, in15638_1, in15638_2, c15276);
    wire[0:0] s15639, in15639_1, in15639_2;
    wire c15639;
    assign in15639_1 = {c15279};
    assign in15639_2 = {s15280[0]};
    Full_Adder FA_15639(s15639, c15639, in15639_1, in15639_2, c15278);
    wire[0:0] s15640, in15640_1, in15640_2;
    wire c15640;
    assign in15640_1 = {c15281};
    assign in15640_2 = {s15282[0]};
    Full_Adder FA_15640(s15640, c15640, in15640_1, in15640_2, c15280);
    wire[0:0] s15641, in15641_1, in15641_2;
    wire c15641;
    assign in15641_1 = {c15283};
    assign in15641_2 = {s15284[0]};
    Full_Adder FA_15641(s15641, c15641, in15641_1, in15641_2, c15282);
    wire[0:0] s15642, in15642_1, in15642_2;
    wire c15642;
    assign in15642_1 = {c15285};
    assign in15642_2 = {s15286[0]};
    Full_Adder FA_15642(s15642, c15642, in15642_1, in15642_2, c15284);
    wire[0:0] s15643, in15643_1, in15643_2;
    wire c15643;
    assign in15643_1 = {c15287};
    assign in15643_2 = {s15288[0]};
    Full_Adder FA_15643(s15643, c15643, in15643_1, in15643_2, c15286);
    wire[0:0] s15644, in15644_1, in15644_2;
    wire c15644;
    assign in15644_1 = {c15289};
    assign in15644_2 = {s15290[0]};
    Full_Adder FA_15644(s15644, c15644, in15644_1, in15644_2, c15288);
    wire[0:0] s15645, in15645_1, in15645_2;
    wire c15645;
    assign in15645_1 = {c15291};
    assign in15645_2 = {s15292[0]};
    Full_Adder FA_15645(s15645, c15645, in15645_1, in15645_2, c15290);
    wire[0:0] s15646, in15646_1, in15646_2;
    wire c15646;
    assign in15646_1 = {c15293};
    assign in15646_2 = {s15294[0]};
    Full_Adder FA_15646(s15646, c15646, in15646_1, in15646_2, c15292);
    wire[0:0] s15647, in15647_1, in15647_2;
    wire c15647;
    assign in15647_1 = {c15295};
    assign in15647_2 = {s15296[0]};
    Full_Adder FA_15647(s15647, c15647, in15647_1, in15647_2, c15294);
    wire[0:0] s15648, in15648_1, in15648_2;
    wire c15648;
    assign in15648_1 = {c15297};
    assign in15648_2 = {s15298[0]};
    Full_Adder FA_15648(s15648, c15648, in15648_1, in15648_2, c15296);
    wire[0:0] s15649, in15649_1, in15649_2;
    wire c15649;
    assign in15649_1 = {c15299};
    assign in15649_2 = {s15300[0]};
    Full_Adder FA_15649(s15649, c15649, in15649_1, in15649_2, c15298);
    wire[0:0] s15650, in15650_1, in15650_2;
    wire c15650;
    assign in15650_1 = {c15301};
    assign in15650_2 = {s15302[0]};
    Full_Adder FA_15650(s15650, c15650, in15650_1, in15650_2, c15300);
    wire[0:0] s15651, in15651_1, in15651_2;
    wire c15651;
    assign in15651_1 = {c15303};
    assign in15651_2 = {s15304[0]};
    Full_Adder FA_15651(s15651, c15651, in15651_1, in15651_2, c15302);
    wire[0:0] s15652, in15652_1, in15652_2;
    wire c15652;
    assign in15652_1 = {c15305};
    assign in15652_2 = {s15306[0]};
    Full_Adder FA_15652(s15652, c15652, in15652_1, in15652_2, c15304);
    wire[0:0] s15653, in15653_1, in15653_2;
    wire c15653;
    assign in15653_1 = {c15307};
    assign in15653_2 = {s15308[0]};
    Full_Adder FA_15653(s15653, c15653, in15653_1, in15653_2, c15306);
    wire[0:0] s15654, in15654_1, in15654_2;
    wire c15654;
    assign in15654_1 = {c15309};
    assign in15654_2 = {s15310[0]};
    Full_Adder FA_15654(s15654, c15654, in15654_1, in15654_2, c15308);
    wire[0:0] s15655, in15655_1, in15655_2;
    wire c15655;
    assign in15655_1 = {c15311};
    assign in15655_2 = {s15312[0]};
    Full_Adder FA_15655(s15655, c15655, in15655_1, in15655_2, c15310);
    wire[0:0] s15656, in15656_1, in15656_2;
    wire c15656;
    assign in15656_1 = {c15313};
    assign in15656_2 = {s15314[0]};
    Full_Adder FA_15656(s15656, c15656, in15656_1, in15656_2, c15312);
    wire[0:0] s15657, in15657_1, in15657_2;
    wire c15657;
    assign in15657_1 = {c15315};
    assign in15657_2 = {s15316[0]};
    Full_Adder FA_15657(s15657, c15657, in15657_1, in15657_2, c15314);
    wire[0:0] s15658, in15658_1, in15658_2;
    wire c15658;
    assign in15658_1 = {c15317};
    assign in15658_2 = {s15318[0]};
    Full_Adder FA_15658(s15658, c15658, in15658_1, in15658_2, c15316);
    wire[0:0] s15659, in15659_1, in15659_2;
    wire c15659;
    assign in15659_1 = {c15319};
    assign in15659_2 = {s15320[0]};
    Full_Adder FA_15659(s15659, c15659, in15659_1, in15659_2, c15318);
    wire[0:0] s15660, in15660_1, in15660_2;
    wire c15660;
    assign in15660_1 = {c15321};
    assign in15660_2 = {s15322[0]};
    Full_Adder FA_15660(s15660, c15660, in15660_1, in15660_2, c15320);
    wire[0:0] s15661, in15661_1, in15661_2;
    wire c15661;
    assign in15661_1 = {c15323};
    assign in15661_2 = {s15324[0]};
    Full_Adder FA_15661(s15661, c15661, in15661_1, in15661_2, c15322);
    wire[0:0] s15662, in15662_1, in15662_2;
    wire c15662;
    assign in15662_1 = {c15325};
    assign in15662_2 = {s15326[0]};
    Full_Adder FA_15662(s15662, c15662, in15662_1, in15662_2, c15324);
    wire[0:0] s15663, in15663_1, in15663_2;
    wire c15663;
    assign in15663_1 = {c15327};
    assign in15663_2 = {s15328[0]};
    Full_Adder FA_15663(s15663, c15663, in15663_1, in15663_2, c15326);
    wire[0:0] s15664, in15664_1, in15664_2;
    wire c15664;
    assign in15664_1 = {c15329};
    assign in15664_2 = {s15330[0]};
    Full_Adder FA_15664(s15664, c15664, in15664_1, in15664_2, c15328);
    wire[0:0] s15665, in15665_1, in15665_2;
    wire c15665;
    assign in15665_1 = {c15331};
    assign in15665_2 = {s15332[0]};
    Full_Adder FA_15665(s15665, c15665, in15665_1, in15665_2, c15330);
    wire[0:0] s15666, in15666_1, in15666_2;
    wire c15666;
    assign in15666_1 = {c15333};
    assign in15666_2 = {s15334[0]};
    Full_Adder FA_15666(s15666, c15666, in15666_1, in15666_2, c15332);
    wire[0:0] s15667, in15667_1, in15667_2;
    wire c15667;
    assign in15667_1 = {c15335};
    assign in15667_2 = {s15336[0]};
    Full_Adder FA_15667(s15667, c15667, in15667_1, in15667_2, c15334);
    wire[0:0] s15668, in15668_1, in15668_2;
    wire c15668;
    assign in15668_1 = {c15337};
    assign in15668_2 = {s15338[0]};
    Full_Adder FA_15668(s15668, c15668, in15668_1, in15668_2, c15336);
    wire[0:0] s15669, in15669_1, in15669_2;
    wire c15669;
    assign in15669_1 = {c15339};
    assign in15669_2 = {s15340[0]};
    Full_Adder FA_15669(s15669, c15669, in15669_1, in15669_2, c15338);
    wire[0:0] s15670, in15670_1, in15670_2;
    wire c15670;
    assign in15670_1 = {c15341};
    assign in15670_2 = {s15342[0]};
    Full_Adder FA_15670(s15670, c15670, in15670_1, in15670_2, c15340);
    wire[0:0] s15671, in15671_1, in15671_2;
    wire c15671;
    assign in15671_1 = {c15343};
    assign in15671_2 = {s15344[0]};
    Full_Adder FA_15671(s15671, c15671, in15671_1, in15671_2, c15342);
    wire[0:0] s15672, in15672_1, in15672_2;
    wire c15672;
    assign in15672_1 = {c15345};
    assign in15672_2 = {s15346[0]};
    Full_Adder FA_15672(s15672, c15672, in15672_1, in15672_2, c15344);
    wire[0:0] s15673, in15673_1, in15673_2;
    wire c15673;
    assign in15673_1 = {c15347};
    assign in15673_2 = {s15348[0]};
    Full_Adder FA_15673(s15673, c15673, in15673_1, in15673_2, c15346);
    wire[0:0] s15674, in15674_1, in15674_2;
    wire c15674;
    assign in15674_1 = {c15349};
    assign in15674_2 = {s15350[0]};
    Full_Adder FA_15674(s15674, c15674, in15674_1, in15674_2, c15348);
    wire[0:0] s15675, in15675_1, in15675_2;
    wire c15675;
    assign in15675_1 = {c15351};
    assign in15675_2 = {s15352[0]};
    Full_Adder FA_15675(s15675, c15675, in15675_1, in15675_2, c15350);
    wire[0:0] s15676, in15676_1, in15676_2;
    wire c15676;
    assign in15676_1 = {c15353};
    assign in15676_2 = {s15354[0]};
    Full_Adder FA_15676(s15676, c15676, in15676_1, in15676_2, c15352);
    wire[0:0] s15677, in15677_1, in15677_2;
    wire c15677;
    assign in15677_1 = {c15355};
    assign in15677_2 = {s15356[0]};
    Full_Adder FA_15677(s15677, c15677, in15677_1, in15677_2, c15354);
    wire[0:0] s15678, in15678_1, in15678_2;
    wire c15678;
    assign in15678_1 = {c15357};
    assign in15678_2 = {s15358[0]};
    Full_Adder FA_15678(s15678, c15678, in15678_1, in15678_2, c15356);
    wire[0:0] s15679, in15679_1, in15679_2;
    wire c15679;
    assign in15679_1 = {c15359};
    assign in15679_2 = {s15360[0]};
    Full_Adder FA_15679(s15679, c15679, in15679_1, in15679_2, c15358);
    wire[0:0] s15680, in15680_1, in15680_2;
    wire c15680;
    assign in15680_1 = {c15361};
    assign in15680_2 = {s15362[0]};
    Full_Adder FA_15680(s15680, c15680, in15680_1, in15680_2, c15360);
    wire[0:0] s15681, in15681_1, in15681_2;
    wire c15681;
    assign in15681_1 = {c15363};
    assign in15681_2 = {s15364[0]};
    Full_Adder FA_15681(s15681, c15681, in15681_1, in15681_2, c15362);
    wire[0:0] s15682, in15682_1, in15682_2;
    wire c15682;
    assign in15682_1 = {c15365};
    assign in15682_2 = {s15366[0]};
    Full_Adder FA_15682(s15682, c15682, in15682_1, in15682_2, c15364);
    wire[0:0] s15683, in15683_1, in15683_2;
    wire c15683;
    assign in15683_1 = {c15367};
    assign in15683_2 = {s15368[0]};
    Full_Adder FA_15683(s15683, c15683, in15683_1, in15683_2, c15366);
    wire[0:0] s15684, in15684_1, in15684_2;
    wire c15684;
    assign in15684_1 = {c15369};
    assign in15684_2 = {s15370[0]};
    Full_Adder FA_15684(s15684, c15684, in15684_1, in15684_2, c15368);
    wire[0:0] s15685, in15685_1, in15685_2;
    wire c15685;
    assign in15685_1 = {c15371};
    assign in15685_2 = {s15372[0]};
    Full_Adder FA_15685(s15685, c15685, in15685_1, in15685_2, c15370);
    wire[0:0] s15686, in15686_1, in15686_2;
    wire c15686;
    assign in15686_1 = {c15373};
    assign in15686_2 = {s15374[0]};
    Full_Adder FA_15686(s15686, c15686, in15686_1, in15686_2, c15372);
    wire[0:0] s15687, in15687_1, in15687_2;
    wire c15687;
    assign in15687_1 = {c15375};
    assign in15687_2 = {s15376[0]};
    Full_Adder FA_15687(s15687, c15687, in15687_1, in15687_2, c15374);
    wire[0:0] s15688, in15688_1, in15688_2;
    wire c15688;
    assign in15688_1 = {c15377};
    assign in15688_2 = {s15378[0]};
    Full_Adder FA_15688(s15688, c15688, in15688_1, in15688_2, c15376);
    wire[0:0] s15689, in15689_1, in15689_2;
    wire c15689;
    assign in15689_1 = {c15379};
    assign in15689_2 = {s15380[0]};
    Full_Adder FA_15689(s15689, c15689, in15689_1, in15689_2, c15378);
    wire[0:0] s15690, in15690_1, in15690_2;
    wire c15690;
    assign in15690_1 = {c15381};
    assign in15690_2 = {s15382[0]};
    Full_Adder FA_15690(s15690, c15690, in15690_1, in15690_2, c15380);
    wire[0:0] s15691, in15691_1, in15691_2;
    wire c15691;
    assign in15691_1 = {c15383};
    assign in15691_2 = {s15384[0]};
    Full_Adder FA_15691(s15691, c15691, in15691_1, in15691_2, c15382);
    wire[0:0] s15692, in15692_1, in15692_2;
    wire c15692;
    assign in15692_1 = {c15385};
    assign in15692_2 = {s15386[0]};
    Full_Adder FA_15692(s15692, c15692, in15692_1, in15692_2, c15384);
    wire[0:0] s15693, in15693_1, in15693_2;
    wire c15693;
    assign in15693_1 = {c15387};
    assign in15693_2 = {s15388[0]};
    Full_Adder FA_15693(s15693, c15693, in15693_1, in15693_2, c15386);
    wire[0:0] s15694, in15694_1, in15694_2;
    wire c15694;
    assign in15694_1 = {c15389};
    assign in15694_2 = {s15390[0]};
    Full_Adder FA_15694(s15694, c15694, in15694_1, in15694_2, c15388);
    wire[0:0] s15695, in15695_1, in15695_2;
    wire c15695;
    assign in15695_1 = {c15391};
    assign in15695_2 = {s15392[0]};
    Full_Adder FA_15695(s15695, c15695, in15695_1, in15695_2, c15390);
    wire[0:0] s15696, in15696_1, in15696_2;
    wire c15696;
    assign in15696_1 = {c15393};
    assign in15696_2 = {s15394[0]};
    Full_Adder FA_15696(s15696, c15696, in15696_1, in15696_2, c15392);
    wire[0:0] s15697, in15697_1, in15697_2;
    wire c15697;
    assign in15697_1 = {c15395};
    assign in15697_2 = {s15396[0]};
    Full_Adder FA_15697(s15697, c15697, in15697_1, in15697_2, c15394);
    wire[0:0] s15698, in15698_1, in15698_2;
    wire c15698;
    assign in15698_1 = {c15397};
    assign in15698_2 = {s15398[0]};
    Full_Adder FA_15698(s15698, c15698, in15698_1, in15698_2, c15396);
    wire[0:0] s15699, in15699_1, in15699_2;
    wire c15699;
    assign in15699_1 = {c15399};
    assign in15699_2 = {s15400[0]};
    Full_Adder FA_15699(s15699, c15699, in15699_1, in15699_2, c15398);
    wire[0:0] s15700, in15700_1, in15700_2;
    wire c15700;
    assign in15700_1 = {c15401};
    assign in15700_2 = {s15402[0]};
    Full_Adder FA_15700(s15700, c15700, in15700_1, in15700_2, c15400);
    wire[0:0] s15701, in15701_1, in15701_2;
    wire c15701;
    assign in15701_1 = {c15403};
    assign in15701_2 = {s15404[0]};
    Full_Adder FA_15701(s15701, c15701, in15701_1, in15701_2, c15402);
    wire[0:0] s15702, in15702_1, in15702_2;
    wire c15702;
    assign in15702_1 = {c15405};
    assign in15702_2 = {s15406[0]};
    Full_Adder FA_15702(s15702, c15702, in15702_1, in15702_2, c15404);
    wire[0:0] s15703, in15703_1, in15703_2;
    wire c15703;
    assign in15703_1 = {c15407};
    assign in15703_2 = {s15408[0]};
    Full_Adder FA_15703(s15703, c15703, in15703_1, in15703_2, c15406);
    wire[0:0] s15704, in15704_1, in15704_2;
    wire c15704;
    assign in15704_1 = {c15409};
    assign in15704_2 = {s15410[0]};
    Full_Adder FA_15704(s15704, c15704, in15704_1, in15704_2, c15408);
    wire[0:0] s15705, in15705_1, in15705_2;
    wire c15705;
    assign in15705_1 = {c15411};
    assign in15705_2 = {s15412[0]};
    Full_Adder FA_15705(s15705, c15705, in15705_1, in15705_2, c15410);
    wire[0:0] s15706, in15706_1, in15706_2;
    wire c15706;
    assign in15706_1 = {c15413};
    assign in15706_2 = {s15414[0]};
    Full_Adder FA_15706(s15706, c15706, in15706_1, in15706_2, c15412);
    wire[0:0] s15707, in15707_1, in15707_2;
    wire c15707;
    assign in15707_1 = {c15415};
    assign in15707_2 = {s15416[0]};
    Full_Adder FA_15707(s15707, c15707, in15707_1, in15707_2, c15414);
    wire[0:0] s15708, in15708_1, in15708_2;
    wire c15708;
    assign in15708_1 = {c15417};
    assign in15708_2 = {s15418[0]};
    Full_Adder FA_15708(s15708, c15708, in15708_1, in15708_2, c15416);
    wire[0:0] s15709, in15709_1, in15709_2;
    wire c15709;
    assign in15709_1 = {c15419};
    assign in15709_2 = {s15420[0]};
    Full_Adder FA_15709(s15709, c15709, in15709_1, in15709_2, c15418);
    wire[0:0] s15710, in15710_1, in15710_2;
    wire c15710;
    assign in15710_1 = {c15421};
    assign in15710_2 = {s15422[0]};
    Full_Adder FA_15710(s15710, c15710, in15710_1, in15710_2, c15420);
    wire[0:0] s15711, in15711_1, in15711_2;
    wire c15711;
    assign in15711_1 = {c15423};
    assign in15711_2 = {s15424[0]};
    Full_Adder FA_15711(s15711, c15711, in15711_1, in15711_2, c15422);
    wire[0:0] s15712, in15712_1, in15712_2;
    wire c15712;
    assign in15712_1 = {c15425};
    assign in15712_2 = {s15426[0]};
    Full_Adder FA_15712(s15712, c15712, in15712_1, in15712_2, c15424);
    wire[0:0] s15713, in15713_1, in15713_2;
    wire c15713;
    assign in15713_1 = {c15427};
    assign in15713_2 = {s15428[0]};
    Full_Adder FA_15713(s15713, c15713, in15713_1, in15713_2, c15426);
    wire[0:0] s15714, in15714_1, in15714_2;
    wire c15714;
    assign in15714_1 = {c15429};
    assign in15714_2 = {s15430[0]};
    Full_Adder FA_15714(s15714, c15714, in15714_1, in15714_2, c15428);
    wire[0:0] s15715, in15715_1, in15715_2;
    wire c15715;
    assign in15715_1 = {c15431};
    assign in15715_2 = {s15432[0]};
    Full_Adder FA_15715(s15715, c15715, in15715_1, in15715_2, c15430);
    wire[0:0] s15716, in15716_1, in15716_2;
    wire c15716;
    assign in15716_1 = {c15433};
    assign in15716_2 = {s15434[0]};
    Full_Adder FA_15716(s15716, c15716, in15716_1, in15716_2, c15432);
    wire[0:0] s15717, in15717_1, in15717_2;
    wire c15717;
    assign in15717_1 = {c15435};
    assign in15717_2 = {s15436[0]};
    Full_Adder FA_15717(s15717, c15717, in15717_1, in15717_2, c15434);
    wire[0:0] s15718, in15718_1, in15718_2;
    wire c15718;
    assign in15718_1 = {c15437};
    assign in15718_2 = {s15438[0]};
    Full_Adder FA_15718(s15718, c15718, in15718_1, in15718_2, c15436);
    wire[0:0] s15719, in15719_1, in15719_2;
    wire c15719;
    assign in15719_1 = {c15439};
    assign in15719_2 = {s15440[0]};
    Full_Adder FA_15719(s15719, c15719, in15719_1, in15719_2, c15438);
    wire[0:0] s15720, in15720_1, in15720_2;
    wire c15720;
    assign in15720_1 = {c15441};
    assign in15720_2 = {s15442[0]};
    Full_Adder FA_15720(s15720, c15720, in15720_1, in15720_2, c15440);
    wire[0:0] s15721, in15721_1, in15721_2;
    wire c15721;
    assign in15721_1 = {c15443};
    assign in15721_2 = {s15444[0]};
    Full_Adder FA_15721(s15721, c15721, in15721_1, in15721_2, c15442);
    wire[0:0] s15722, in15722_1, in15722_2;
    wire c15722;
    assign in15722_1 = {c15445};
    assign in15722_2 = {s15446[0]};
    Full_Adder FA_15722(s15722, c15722, in15722_1, in15722_2, c15444);
    wire[0:0] s15723, in15723_1, in15723_2;
    wire c15723;
    assign in15723_1 = {c15447};
    assign in15723_2 = {s15448[0]};
    Full_Adder FA_15723(s15723, c15723, in15723_1, in15723_2, c15446);
    wire[0:0] s15724, in15724_1, in15724_2;
    wire c15724;
    assign in15724_1 = {c15449};
    assign in15724_2 = {s15450[0]};
    Full_Adder FA_15724(s15724, c15724, in15724_1, in15724_2, c15448);
    wire[0:0] s15725, in15725_1, in15725_2;
    wire c15725;
    assign in15725_1 = {c15451};
    assign in15725_2 = {s15452[0]};
    Full_Adder FA_15725(s15725, c15725, in15725_1, in15725_2, c15450);
    wire[0:0] s15726, in15726_1, in15726_2;
    wire c15726;
    assign in15726_1 = {c15453};
    assign in15726_2 = {s15454[0]};
    Full_Adder FA_15726(s15726, c15726, in15726_1, in15726_2, c15452);
    wire[0:0] s15727, in15727_1, in15727_2;
    wire c15727;
    assign in15727_1 = {c15455};
    assign in15727_2 = {s15456[0]};
    Full_Adder FA_15727(s15727, c15727, in15727_1, in15727_2, c15454);
    wire[0:0] s15728, in15728_1, in15728_2;
    wire c15728;
    assign in15728_1 = {c15457};
    assign in15728_2 = {s15458[0]};
    Full_Adder FA_15728(s15728, c15728, in15728_1, in15728_2, c15456);
    wire[0:0] s15729, in15729_1, in15729_2;
    wire c15729;
    assign in15729_1 = {c15459};
    assign in15729_2 = {s15460[0]};
    Full_Adder FA_15729(s15729, c15729, in15729_1, in15729_2, c15458);
    wire[0:0] s15730, in15730_1, in15730_2;
    wire c15730;
    assign in15730_1 = {c15461};
    assign in15730_2 = {s15462[0]};
    Full_Adder FA_15730(s15730, c15730, in15730_1, in15730_2, c15460);
    wire[0:0] s15731, in15731_1, in15731_2;
    wire c15731;
    assign in15731_1 = {c15463};
    assign in15731_2 = {s15464[0]};
    Full_Adder FA_15731(s15731, c15731, in15731_1, in15731_2, c15462);
    wire[0:0] s15732, in15732_1, in15732_2;
    wire c15732;
    assign in15732_1 = {c15465};
    assign in15732_2 = {s15466[0]};
    Full_Adder FA_15732(s15732, c15732, in15732_1, in15732_2, c15464);
    wire[0:0] s15733, in15733_1, in15733_2;
    wire c15733;
    assign in15733_1 = {c15467};
    assign in15733_2 = {s15468[0]};
    Full_Adder FA_15733(s15733, c15733, in15733_1, in15733_2, c15466);
    wire[0:0] s15734, in15734_1, in15734_2;
    wire c15734;
    assign in15734_1 = {c15469};
    assign in15734_2 = {s15470[0]};
    Full_Adder FA_15734(s15734, c15734, in15734_1, in15734_2, c15468);
    wire[0:0] s15735, in15735_1, in15735_2;
    wire c15735;
    assign in15735_1 = {c15471};
    assign in15735_2 = {s15472[0]};
    Full_Adder FA_15735(s15735, c15735, in15735_1, in15735_2, c15470);
    wire[0:0] s15736, in15736_1, in15736_2;
    wire c15736;
    assign in15736_1 = {c15473};
    assign in15736_2 = {s15474[0]};
    Full_Adder FA_15736(s15736, c15736, in15736_1, in15736_2, c15472);
    wire[0:0] s15737, in15737_1, in15737_2;
    wire c15737;
    assign in15737_1 = {c15475};
    assign in15737_2 = {s15476[0]};
    Full_Adder FA_15737(s15737, c15737, in15737_1, in15737_2, c15474);
    wire[0:0] s15738, in15738_1, in15738_2;
    wire c15738;
    assign in15738_1 = {c15477};
    assign in15738_2 = {s15478[0]};
    Full_Adder FA_15738(s15738, c15738, in15738_1, in15738_2, c15476);
    wire[0:0] s15739, in15739_1, in15739_2;
    wire c15739;
    assign in15739_1 = {c15479};
    assign in15739_2 = {s15480[0]};
    Full_Adder FA_15739(s15739, c15739, in15739_1, in15739_2, c15478);
    wire[0:0] s15740, in15740_1, in15740_2;
    wire c15740;
    assign in15740_1 = {c15481};
    assign in15740_2 = {s15482[0]};
    Full_Adder FA_15740(s15740, c15740, in15740_1, in15740_2, c15480);
    wire[0:0] s15741, in15741_1, in15741_2;
    wire c15741;
    assign in15741_1 = {c15483};
    assign in15741_2 = {s15484[0]};
    Full_Adder FA_15741(s15741, c15741, in15741_1, in15741_2, c15482);
    wire[0:0] s15742, in15742_1, in15742_2;
    wire c15742;
    assign in15742_1 = {c15485};
    assign in15742_2 = {s15486[0]};
    Full_Adder FA_15742(s15742, c15742, in15742_1, in15742_2, c15484);
    wire[0:0] s15743, in15743_1, in15743_2;
    wire c15743;
    assign in15743_1 = {c15487};
    assign in15743_2 = {s15488[0]};
    Full_Adder FA_15743(s15743, c15743, in15743_1, in15743_2, c15486);
    wire[0:0] s15744, in15744_1, in15744_2;
    wire c15744;
    assign in15744_1 = {c15489};
    assign in15744_2 = {s15490[0]};
    Full_Adder FA_15744(s15744, c15744, in15744_1, in15744_2, c15488);
    wire[0:0] s15745, in15745_1, in15745_2;
    wire c15745;
    assign in15745_1 = {c15491};
    assign in15745_2 = {s15492[0]};
    Full_Adder FA_15745(s15745, c15745, in15745_1, in15745_2, c15490);
    wire[0:0] s15746, in15746_1, in15746_2;
    wire c15746;
    assign in15746_1 = {c15493};
    assign in15746_2 = {s15494[0]};
    Full_Adder FA_15746(s15746, c15746, in15746_1, in15746_2, c15492);
    wire[0:0] s15747, in15747_1, in15747_2;
    wire c15747;
    assign in15747_1 = {c15495};
    assign in15747_2 = {s15496[0]};
    Full_Adder FA_15747(s15747, c15747, in15747_1, in15747_2, c15494);
    wire[0:0] s15748, in15748_1, in15748_2;
    wire c15748;
    assign in15748_1 = {c15497};
    assign in15748_2 = {s15498[0]};
    Full_Adder FA_15748(s15748, c15748, in15748_1, in15748_2, c15496);
    wire[0:0] s15749, in15749_1, in15749_2;
    wire c15749;
    assign in15749_1 = {c15498};
    assign in15749_2 = {c15499};
    Full_Adder FA_15749(s15749, c15749, in15749_1, in15749_2, pp127[124]);
    wire[0:0] s15750, in15750_1, in15750_2;
    wire c15750;
    assign in15750_1 = {pp126[126]};
    assign in15750_2 = {pp127[125]};
    Full_Adder FA_15750(s15750, c15750, in15750_1, in15750_2, pp125[127]);

    /*Stage 11*/
    wire[0:0] s15751, in15751_1, in15751_2;
    wire c15751;
    assign in15751_1 = {pp0[2]};
    assign in15751_2 = {pp1[1]};
    Half_Adder HA_15751(s15751, c15751, in15751_1, in15751_2);
    wire[0:0] s15752, in15752_1, in15752_2;
    wire c15752;
    assign in15752_1 = {pp3[0]};
    assign in15752_2 = {s15501[0]};
    Full_Adder FA_15752(s15752, c15752, in15752_1, in15752_2, pp2[1]);
    wire[0:0] s15753, in15753_1, in15753_2;
    wire c15753;
    assign in15753_1 = {c15501};
    assign in15753_2 = {s15502[0]};
    Full_Adder FA_15753(s15753, c15753, in15753_1, in15753_2, s15007[0]);
    wire[0:0] s15754, in15754_1, in15754_2;
    wire c15754;
    assign in15754_1 = {c15502};
    assign in15754_2 = {s15503[0]};
    Full_Adder FA_15754(s15754, c15754, in15754_1, in15754_2, s15009[0]);
    wire[0:0] s15755, in15755_1, in15755_2;
    wire c15755;
    assign in15755_1 = {c15503};
    assign in15755_2 = {s15504[0]};
    Full_Adder FA_15755(s15755, c15755, in15755_1, in15755_2, s15011[0]);
    wire[0:0] s15756, in15756_1, in15756_2;
    wire c15756;
    assign in15756_1 = {c15504};
    assign in15756_2 = {s15505[0]};
    Full_Adder FA_15756(s15756, c15756, in15756_1, in15756_2, s15013[0]);
    wire[0:0] s15757, in15757_1, in15757_2;
    wire c15757;
    assign in15757_1 = {c15505};
    assign in15757_2 = {s15506[0]};
    Full_Adder FA_15757(s15757, c15757, in15757_1, in15757_2, s15015[0]);
    wire[0:0] s15758, in15758_1, in15758_2;
    wire c15758;
    assign in15758_1 = {c15506};
    assign in15758_2 = {s15507[0]};
    Full_Adder FA_15758(s15758, c15758, in15758_1, in15758_2, s15017[0]);
    wire[0:0] s15759, in15759_1, in15759_2;
    wire c15759;
    assign in15759_1 = {c15507};
    assign in15759_2 = {s15508[0]};
    Full_Adder FA_15759(s15759, c15759, in15759_1, in15759_2, s15019[0]);
    wire[0:0] s15760, in15760_1, in15760_2;
    wire c15760;
    assign in15760_1 = {c15508};
    assign in15760_2 = {s15509[0]};
    Full_Adder FA_15760(s15760, c15760, in15760_1, in15760_2, s15021[0]);
    wire[0:0] s15761, in15761_1, in15761_2;
    wire c15761;
    assign in15761_1 = {c15509};
    assign in15761_2 = {s15510[0]};
    Full_Adder FA_15761(s15761, c15761, in15761_1, in15761_2, s15023[0]);
    wire[0:0] s15762, in15762_1, in15762_2;
    wire c15762;
    assign in15762_1 = {c15510};
    assign in15762_2 = {s15511[0]};
    Full_Adder FA_15762(s15762, c15762, in15762_1, in15762_2, s15025[0]);
    wire[0:0] s15763, in15763_1, in15763_2;
    wire c15763;
    assign in15763_1 = {c15511};
    assign in15763_2 = {s15512[0]};
    Full_Adder FA_15763(s15763, c15763, in15763_1, in15763_2, s15027[0]);
    wire[0:0] s15764, in15764_1, in15764_2;
    wire c15764;
    assign in15764_1 = {c15512};
    assign in15764_2 = {s15513[0]};
    Full_Adder FA_15764(s15764, c15764, in15764_1, in15764_2, s15029[0]);
    wire[0:0] s15765, in15765_1, in15765_2;
    wire c15765;
    assign in15765_1 = {c15513};
    assign in15765_2 = {s15514[0]};
    Full_Adder FA_15765(s15765, c15765, in15765_1, in15765_2, s15031[0]);
    wire[0:0] s15766, in15766_1, in15766_2;
    wire c15766;
    assign in15766_1 = {c15514};
    assign in15766_2 = {s15515[0]};
    Full_Adder FA_15766(s15766, c15766, in15766_1, in15766_2, s15033[0]);
    wire[0:0] s15767, in15767_1, in15767_2;
    wire c15767;
    assign in15767_1 = {c15515};
    assign in15767_2 = {s15516[0]};
    Full_Adder FA_15767(s15767, c15767, in15767_1, in15767_2, s15035[0]);
    wire[0:0] s15768, in15768_1, in15768_2;
    wire c15768;
    assign in15768_1 = {c15516};
    assign in15768_2 = {s15517[0]};
    Full_Adder FA_15768(s15768, c15768, in15768_1, in15768_2, s15037[0]);
    wire[0:0] s15769, in15769_1, in15769_2;
    wire c15769;
    assign in15769_1 = {c15517};
    assign in15769_2 = {s15518[0]};
    Full_Adder FA_15769(s15769, c15769, in15769_1, in15769_2, s15039[0]);
    wire[0:0] s15770, in15770_1, in15770_2;
    wire c15770;
    assign in15770_1 = {c15518};
    assign in15770_2 = {s15519[0]};
    Full_Adder FA_15770(s15770, c15770, in15770_1, in15770_2, s15041[0]);
    wire[0:0] s15771, in15771_1, in15771_2;
    wire c15771;
    assign in15771_1 = {c15519};
    assign in15771_2 = {s15520[0]};
    Full_Adder FA_15771(s15771, c15771, in15771_1, in15771_2, s15043[0]);
    wire[0:0] s15772, in15772_1, in15772_2;
    wire c15772;
    assign in15772_1 = {c15520};
    assign in15772_2 = {s15521[0]};
    Full_Adder FA_15772(s15772, c15772, in15772_1, in15772_2, s15045[0]);
    wire[0:0] s15773, in15773_1, in15773_2;
    wire c15773;
    assign in15773_1 = {c15521};
    assign in15773_2 = {s15522[0]};
    Full_Adder FA_15773(s15773, c15773, in15773_1, in15773_2, s15047[0]);
    wire[0:0] s15774, in15774_1, in15774_2;
    wire c15774;
    assign in15774_1 = {c15522};
    assign in15774_2 = {s15523[0]};
    Full_Adder FA_15774(s15774, c15774, in15774_1, in15774_2, s15049[0]);
    wire[0:0] s15775, in15775_1, in15775_2;
    wire c15775;
    assign in15775_1 = {c15523};
    assign in15775_2 = {s15524[0]};
    Full_Adder FA_15775(s15775, c15775, in15775_1, in15775_2, s15051[0]);
    wire[0:0] s15776, in15776_1, in15776_2;
    wire c15776;
    assign in15776_1 = {c15524};
    assign in15776_2 = {s15525[0]};
    Full_Adder FA_15776(s15776, c15776, in15776_1, in15776_2, s15053[0]);
    wire[0:0] s15777, in15777_1, in15777_2;
    wire c15777;
    assign in15777_1 = {c15525};
    assign in15777_2 = {s15526[0]};
    Full_Adder FA_15777(s15777, c15777, in15777_1, in15777_2, s15055[0]);
    wire[0:0] s15778, in15778_1, in15778_2;
    wire c15778;
    assign in15778_1 = {c15526};
    assign in15778_2 = {s15527[0]};
    Full_Adder FA_15778(s15778, c15778, in15778_1, in15778_2, s15057[0]);
    wire[0:0] s15779, in15779_1, in15779_2;
    wire c15779;
    assign in15779_1 = {c15527};
    assign in15779_2 = {s15528[0]};
    Full_Adder FA_15779(s15779, c15779, in15779_1, in15779_2, s15059[0]);
    wire[0:0] s15780, in15780_1, in15780_2;
    wire c15780;
    assign in15780_1 = {c15528};
    assign in15780_2 = {s15529[0]};
    Full_Adder FA_15780(s15780, c15780, in15780_1, in15780_2, s15061[0]);
    wire[0:0] s15781, in15781_1, in15781_2;
    wire c15781;
    assign in15781_1 = {c15529};
    assign in15781_2 = {s15530[0]};
    Full_Adder FA_15781(s15781, c15781, in15781_1, in15781_2, s15063[0]);
    wire[0:0] s15782, in15782_1, in15782_2;
    wire c15782;
    assign in15782_1 = {c15530};
    assign in15782_2 = {s15531[0]};
    Full_Adder FA_15782(s15782, c15782, in15782_1, in15782_2, s15065[0]);
    wire[0:0] s15783, in15783_1, in15783_2;
    wire c15783;
    assign in15783_1 = {c15531};
    assign in15783_2 = {s15532[0]};
    Full_Adder FA_15783(s15783, c15783, in15783_1, in15783_2, s15067[0]);
    wire[0:0] s15784, in15784_1, in15784_2;
    wire c15784;
    assign in15784_1 = {c15532};
    assign in15784_2 = {s15533[0]};
    Full_Adder FA_15784(s15784, c15784, in15784_1, in15784_2, s15069[0]);
    wire[0:0] s15785, in15785_1, in15785_2;
    wire c15785;
    assign in15785_1 = {c15533};
    assign in15785_2 = {s15534[0]};
    Full_Adder FA_15785(s15785, c15785, in15785_1, in15785_2, s15071[0]);
    wire[0:0] s15786, in15786_1, in15786_2;
    wire c15786;
    assign in15786_1 = {c15534};
    assign in15786_2 = {s15535[0]};
    Full_Adder FA_15786(s15786, c15786, in15786_1, in15786_2, s15073[0]);
    wire[0:0] s15787, in15787_1, in15787_2;
    wire c15787;
    assign in15787_1 = {c15535};
    assign in15787_2 = {s15536[0]};
    Full_Adder FA_15787(s15787, c15787, in15787_1, in15787_2, s15075[0]);
    wire[0:0] s15788, in15788_1, in15788_2;
    wire c15788;
    assign in15788_1 = {c15536};
    assign in15788_2 = {s15537[0]};
    Full_Adder FA_15788(s15788, c15788, in15788_1, in15788_2, s15077[0]);
    wire[0:0] s15789, in15789_1, in15789_2;
    wire c15789;
    assign in15789_1 = {c15537};
    assign in15789_2 = {s15538[0]};
    Full_Adder FA_15789(s15789, c15789, in15789_1, in15789_2, s15079[0]);
    wire[0:0] s15790, in15790_1, in15790_2;
    wire c15790;
    assign in15790_1 = {c15538};
    assign in15790_2 = {s15539[0]};
    Full_Adder FA_15790(s15790, c15790, in15790_1, in15790_2, s15081[0]);
    wire[0:0] s15791, in15791_1, in15791_2;
    wire c15791;
    assign in15791_1 = {c15539};
    assign in15791_2 = {s15540[0]};
    Full_Adder FA_15791(s15791, c15791, in15791_1, in15791_2, s15083[0]);
    wire[0:0] s15792, in15792_1, in15792_2;
    wire c15792;
    assign in15792_1 = {c15540};
    assign in15792_2 = {s15541[0]};
    Full_Adder FA_15792(s15792, c15792, in15792_1, in15792_2, s15085[0]);
    wire[0:0] s15793, in15793_1, in15793_2;
    wire c15793;
    assign in15793_1 = {c15541};
    assign in15793_2 = {s15542[0]};
    Full_Adder FA_15793(s15793, c15793, in15793_1, in15793_2, s15087[0]);
    wire[0:0] s15794, in15794_1, in15794_2;
    wire c15794;
    assign in15794_1 = {c15542};
    assign in15794_2 = {s15543[0]};
    Full_Adder FA_15794(s15794, c15794, in15794_1, in15794_2, s15089[0]);
    wire[0:0] s15795, in15795_1, in15795_2;
    wire c15795;
    assign in15795_1 = {c15543};
    assign in15795_2 = {s15544[0]};
    Full_Adder FA_15795(s15795, c15795, in15795_1, in15795_2, s15091[0]);
    wire[0:0] s15796, in15796_1, in15796_2;
    wire c15796;
    assign in15796_1 = {c15544};
    assign in15796_2 = {s15545[0]};
    Full_Adder FA_15796(s15796, c15796, in15796_1, in15796_2, s15093[0]);
    wire[0:0] s15797, in15797_1, in15797_2;
    wire c15797;
    assign in15797_1 = {c15545};
    assign in15797_2 = {s15546[0]};
    Full_Adder FA_15797(s15797, c15797, in15797_1, in15797_2, s15095[0]);
    wire[0:0] s15798, in15798_1, in15798_2;
    wire c15798;
    assign in15798_1 = {c15546};
    assign in15798_2 = {s15547[0]};
    Full_Adder FA_15798(s15798, c15798, in15798_1, in15798_2, s15097[0]);
    wire[0:0] s15799, in15799_1, in15799_2;
    wire c15799;
    assign in15799_1 = {c15547};
    assign in15799_2 = {s15548[0]};
    Full_Adder FA_15799(s15799, c15799, in15799_1, in15799_2, s15099[0]);
    wire[0:0] s15800, in15800_1, in15800_2;
    wire c15800;
    assign in15800_1 = {c15548};
    assign in15800_2 = {s15549[0]};
    Full_Adder FA_15800(s15800, c15800, in15800_1, in15800_2, s15101[0]);
    wire[0:0] s15801, in15801_1, in15801_2;
    wire c15801;
    assign in15801_1 = {c15549};
    assign in15801_2 = {s15550[0]};
    Full_Adder FA_15801(s15801, c15801, in15801_1, in15801_2, s15103[0]);
    wire[0:0] s15802, in15802_1, in15802_2;
    wire c15802;
    assign in15802_1 = {c15550};
    assign in15802_2 = {s15551[0]};
    Full_Adder FA_15802(s15802, c15802, in15802_1, in15802_2, s15105[0]);
    wire[0:0] s15803, in15803_1, in15803_2;
    wire c15803;
    assign in15803_1 = {c15551};
    assign in15803_2 = {s15552[0]};
    Full_Adder FA_15803(s15803, c15803, in15803_1, in15803_2, s15107[0]);
    wire[0:0] s15804, in15804_1, in15804_2;
    wire c15804;
    assign in15804_1 = {c15552};
    assign in15804_2 = {s15553[0]};
    Full_Adder FA_15804(s15804, c15804, in15804_1, in15804_2, s15109[0]);
    wire[0:0] s15805, in15805_1, in15805_2;
    wire c15805;
    assign in15805_1 = {c15553};
    assign in15805_2 = {s15554[0]};
    Full_Adder FA_15805(s15805, c15805, in15805_1, in15805_2, s15111[0]);
    wire[0:0] s15806, in15806_1, in15806_2;
    wire c15806;
    assign in15806_1 = {c15554};
    assign in15806_2 = {s15555[0]};
    Full_Adder FA_15806(s15806, c15806, in15806_1, in15806_2, s15113[0]);
    wire[0:0] s15807, in15807_1, in15807_2;
    wire c15807;
    assign in15807_1 = {c15555};
    assign in15807_2 = {s15556[0]};
    Full_Adder FA_15807(s15807, c15807, in15807_1, in15807_2, s15115[0]);
    wire[0:0] s15808, in15808_1, in15808_2;
    wire c15808;
    assign in15808_1 = {c15556};
    assign in15808_2 = {s15557[0]};
    Full_Adder FA_15808(s15808, c15808, in15808_1, in15808_2, s15117[0]);
    wire[0:0] s15809, in15809_1, in15809_2;
    wire c15809;
    assign in15809_1 = {c15557};
    assign in15809_2 = {s15558[0]};
    Full_Adder FA_15809(s15809, c15809, in15809_1, in15809_2, s15119[0]);
    wire[0:0] s15810, in15810_1, in15810_2;
    wire c15810;
    assign in15810_1 = {c15558};
    assign in15810_2 = {s15559[0]};
    Full_Adder FA_15810(s15810, c15810, in15810_1, in15810_2, s15121[0]);
    wire[0:0] s15811, in15811_1, in15811_2;
    wire c15811;
    assign in15811_1 = {c15559};
    assign in15811_2 = {s15560[0]};
    Full_Adder FA_15811(s15811, c15811, in15811_1, in15811_2, s15123[0]);
    wire[0:0] s15812, in15812_1, in15812_2;
    wire c15812;
    assign in15812_1 = {c15560};
    assign in15812_2 = {s15561[0]};
    Full_Adder FA_15812(s15812, c15812, in15812_1, in15812_2, s15125[0]);
    wire[0:0] s15813, in15813_1, in15813_2;
    wire c15813;
    assign in15813_1 = {c15561};
    assign in15813_2 = {s15562[0]};
    Full_Adder FA_15813(s15813, c15813, in15813_1, in15813_2, s15127[0]);
    wire[0:0] s15814, in15814_1, in15814_2;
    wire c15814;
    assign in15814_1 = {c15562};
    assign in15814_2 = {s15563[0]};
    Full_Adder FA_15814(s15814, c15814, in15814_1, in15814_2, s15129[0]);
    wire[0:0] s15815, in15815_1, in15815_2;
    wire c15815;
    assign in15815_1 = {c15563};
    assign in15815_2 = {s15564[0]};
    Full_Adder FA_15815(s15815, c15815, in15815_1, in15815_2, s15131[0]);
    wire[0:0] s15816, in15816_1, in15816_2;
    wire c15816;
    assign in15816_1 = {c15564};
    assign in15816_2 = {s15565[0]};
    Full_Adder FA_15816(s15816, c15816, in15816_1, in15816_2, s15133[0]);
    wire[0:0] s15817, in15817_1, in15817_2;
    wire c15817;
    assign in15817_1 = {c15565};
    assign in15817_2 = {s15566[0]};
    Full_Adder FA_15817(s15817, c15817, in15817_1, in15817_2, s15135[0]);
    wire[0:0] s15818, in15818_1, in15818_2;
    wire c15818;
    assign in15818_1 = {c15566};
    assign in15818_2 = {s15567[0]};
    Full_Adder FA_15818(s15818, c15818, in15818_1, in15818_2, s15137[0]);
    wire[0:0] s15819, in15819_1, in15819_2;
    wire c15819;
    assign in15819_1 = {c15567};
    assign in15819_2 = {s15568[0]};
    Full_Adder FA_15819(s15819, c15819, in15819_1, in15819_2, s15139[0]);
    wire[0:0] s15820, in15820_1, in15820_2;
    wire c15820;
    assign in15820_1 = {c15568};
    assign in15820_2 = {s15569[0]};
    Full_Adder FA_15820(s15820, c15820, in15820_1, in15820_2, s15141[0]);
    wire[0:0] s15821, in15821_1, in15821_2;
    wire c15821;
    assign in15821_1 = {c15569};
    assign in15821_2 = {s15570[0]};
    Full_Adder FA_15821(s15821, c15821, in15821_1, in15821_2, s15143[0]);
    wire[0:0] s15822, in15822_1, in15822_2;
    wire c15822;
    assign in15822_1 = {c15570};
    assign in15822_2 = {s15571[0]};
    Full_Adder FA_15822(s15822, c15822, in15822_1, in15822_2, s15145[0]);
    wire[0:0] s15823, in15823_1, in15823_2;
    wire c15823;
    assign in15823_1 = {c15571};
    assign in15823_2 = {s15572[0]};
    Full_Adder FA_15823(s15823, c15823, in15823_1, in15823_2, s15147[0]);
    wire[0:0] s15824, in15824_1, in15824_2;
    wire c15824;
    assign in15824_1 = {c15572};
    assign in15824_2 = {s15573[0]};
    Full_Adder FA_15824(s15824, c15824, in15824_1, in15824_2, s15149[0]);
    wire[0:0] s15825, in15825_1, in15825_2;
    wire c15825;
    assign in15825_1 = {c15573};
    assign in15825_2 = {s15574[0]};
    Full_Adder FA_15825(s15825, c15825, in15825_1, in15825_2, s15151[0]);
    wire[0:0] s15826, in15826_1, in15826_2;
    wire c15826;
    assign in15826_1 = {c15574};
    assign in15826_2 = {s15575[0]};
    Full_Adder FA_15826(s15826, c15826, in15826_1, in15826_2, s15153[0]);
    wire[0:0] s15827, in15827_1, in15827_2;
    wire c15827;
    assign in15827_1 = {c15575};
    assign in15827_2 = {s15576[0]};
    Full_Adder FA_15827(s15827, c15827, in15827_1, in15827_2, s15155[0]);
    wire[0:0] s15828, in15828_1, in15828_2;
    wire c15828;
    assign in15828_1 = {c15576};
    assign in15828_2 = {s15577[0]};
    Full_Adder FA_15828(s15828, c15828, in15828_1, in15828_2, s15157[0]);
    wire[0:0] s15829, in15829_1, in15829_2;
    wire c15829;
    assign in15829_1 = {c15577};
    assign in15829_2 = {s15578[0]};
    Full_Adder FA_15829(s15829, c15829, in15829_1, in15829_2, s15159[0]);
    wire[0:0] s15830, in15830_1, in15830_2;
    wire c15830;
    assign in15830_1 = {c15578};
    assign in15830_2 = {s15579[0]};
    Full_Adder FA_15830(s15830, c15830, in15830_1, in15830_2, s15161[0]);
    wire[0:0] s15831, in15831_1, in15831_2;
    wire c15831;
    assign in15831_1 = {c15579};
    assign in15831_2 = {s15580[0]};
    Full_Adder FA_15831(s15831, c15831, in15831_1, in15831_2, s15163[0]);
    wire[0:0] s15832, in15832_1, in15832_2;
    wire c15832;
    assign in15832_1 = {c15580};
    assign in15832_2 = {s15581[0]};
    Full_Adder FA_15832(s15832, c15832, in15832_1, in15832_2, s15165[0]);
    wire[0:0] s15833, in15833_1, in15833_2;
    wire c15833;
    assign in15833_1 = {c15581};
    assign in15833_2 = {s15582[0]};
    Full_Adder FA_15833(s15833, c15833, in15833_1, in15833_2, s15167[0]);
    wire[0:0] s15834, in15834_1, in15834_2;
    wire c15834;
    assign in15834_1 = {c15582};
    assign in15834_2 = {s15583[0]};
    Full_Adder FA_15834(s15834, c15834, in15834_1, in15834_2, s15169[0]);
    wire[0:0] s15835, in15835_1, in15835_2;
    wire c15835;
    assign in15835_1 = {c15583};
    assign in15835_2 = {s15584[0]};
    Full_Adder FA_15835(s15835, c15835, in15835_1, in15835_2, s15171[0]);
    wire[0:0] s15836, in15836_1, in15836_2;
    wire c15836;
    assign in15836_1 = {c15584};
    assign in15836_2 = {s15585[0]};
    Full_Adder FA_15836(s15836, c15836, in15836_1, in15836_2, s15173[0]);
    wire[0:0] s15837, in15837_1, in15837_2;
    wire c15837;
    assign in15837_1 = {c15585};
    assign in15837_2 = {s15586[0]};
    Full_Adder FA_15837(s15837, c15837, in15837_1, in15837_2, s15175[0]);
    wire[0:0] s15838, in15838_1, in15838_2;
    wire c15838;
    assign in15838_1 = {c15586};
    assign in15838_2 = {s15587[0]};
    Full_Adder FA_15838(s15838, c15838, in15838_1, in15838_2, s15177[0]);
    wire[0:0] s15839, in15839_1, in15839_2;
    wire c15839;
    assign in15839_1 = {c15587};
    assign in15839_2 = {s15588[0]};
    Full_Adder FA_15839(s15839, c15839, in15839_1, in15839_2, s15179[0]);
    wire[0:0] s15840, in15840_1, in15840_2;
    wire c15840;
    assign in15840_1 = {c15588};
    assign in15840_2 = {s15589[0]};
    Full_Adder FA_15840(s15840, c15840, in15840_1, in15840_2, s15181[0]);
    wire[0:0] s15841, in15841_1, in15841_2;
    wire c15841;
    assign in15841_1 = {c15589};
    assign in15841_2 = {s15590[0]};
    Full_Adder FA_15841(s15841, c15841, in15841_1, in15841_2, s15183[0]);
    wire[0:0] s15842, in15842_1, in15842_2;
    wire c15842;
    assign in15842_1 = {c15590};
    assign in15842_2 = {s15591[0]};
    Full_Adder FA_15842(s15842, c15842, in15842_1, in15842_2, s15185[0]);
    wire[0:0] s15843, in15843_1, in15843_2;
    wire c15843;
    assign in15843_1 = {c15591};
    assign in15843_2 = {s15592[0]};
    Full_Adder FA_15843(s15843, c15843, in15843_1, in15843_2, s15187[0]);
    wire[0:0] s15844, in15844_1, in15844_2;
    wire c15844;
    assign in15844_1 = {c15592};
    assign in15844_2 = {s15593[0]};
    Full_Adder FA_15844(s15844, c15844, in15844_1, in15844_2, s15189[0]);
    wire[0:0] s15845, in15845_1, in15845_2;
    wire c15845;
    assign in15845_1 = {c15593};
    assign in15845_2 = {s15594[0]};
    Full_Adder FA_15845(s15845, c15845, in15845_1, in15845_2, s15191[0]);
    wire[0:0] s15846, in15846_1, in15846_2;
    wire c15846;
    assign in15846_1 = {c15594};
    assign in15846_2 = {s15595[0]};
    Full_Adder FA_15846(s15846, c15846, in15846_1, in15846_2, s15193[0]);
    wire[0:0] s15847, in15847_1, in15847_2;
    wire c15847;
    assign in15847_1 = {c15595};
    assign in15847_2 = {s15596[0]};
    Full_Adder FA_15847(s15847, c15847, in15847_1, in15847_2, s15195[0]);
    wire[0:0] s15848, in15848_1, in15848_2;
    wire c15848;
    assign in15848_1 = {c15596};
    assign in15848_2 = {s15597[0]};
    Full_Adder FA_15848(s15848, c15848, in15848_1, in15848_2, s15197[0]);
    wire[0:0] s15849, in15849_1, in15849_2;
    wire c15849;
    assign in15849_1 = {c15597};
    assign in15849_2 = {s15598[0]};
    Full_Adder FA_15849(s15849, c15849, in15849_1, in15849_2, s15199[0]);
    wire[0:0] s15850, in15850_1, in15850_2;
    wire c15850;
    assign in15850_1 = {c15598};
    assign in15850_2 = {s15599[0]};
    Full_Adder FA_15850(s15850, c15850, in15850_1, in15850_2, s15201[0]);
    wire[0:0] s15851, in15851_1, in15851_2;
    wire c15851;
    assign in15851_1 = {c15599};
    assign in15851_2 = {s15600[0]};
    Full_Adder FA_15851(s15851, c15851, in15851_1, in15851_2, s15203[0]);
    wire[0:0] s15852, in15852_1, in15852_2;
    wire c15852;
    assign in15852_1 = {c15600};
    assign in15852_2 = {s15601[0]};
    Full_Adder FA_15852(s15852, c15852, in15852_1, in15852_2, s15205[0]);
    wire[0:0] s15853, in15853_1, in15853_2;
    wire c15853;
    assign in15853_1 = {c15601};
    assign in15853_2 = {s15602[0]};
    Full_Adder FA_15853(s15853, c15853, in15853_1, in15853_2, s15207[0]);
    wire[0:0] s15854, in15854_1, in15854_2;
    wire c15854;
    assign in15854_1 = {c15602};
    assign in15854_2 = {s15603[0]};
    Full_Adder FA_15854(s15854, c15854, in15854_1, in15854_2, s15209[0]);
    wire[0:0] s15855, in15855_1, in15855_2;
    wire c15855;
    assign in15855_1 = {c15603};
    assign in15855_2 = {s15604[0]};
    Full_Adder FA_15855(s15855, c15855, in15855_1, in15855_2, s15211[0]);
    wire[0:0] s15856, in15856_1, in15856_2;
    wire c15856;
    assign in15856_1 = {c15604};
    assign in15856_2 = {s15605[0]};
    Full_Adder FA_15856(s15856, c15856, in15856_1, in15856_2, s15213[0]);
    wire[0:0] s15857, in15857_1, in15857_2;
    wire c15857;
    assign in15857_1 = {c15605};
    assign in15857_2 = {s15606[0]};
    Full_Adder FA_15857(s15857, c15857, in15857_1, in15857_2, s15215[0]);
    wire[0:0] s15858, in15858_1, in15858_2;
    wire c15858;
    assign in15858_1 = {c15606};
    assign in15858_2 = {s15607[0]};
    Full_Adder FA_15858(s15858, c15858, in15858_1, in15858_2, s15217[0]);
    wire[0:0] s15859, in15859_1, in15859_2;
    wire c15859;
    assign in15859_1 = {c15607};
    assign in15859_2 = {s15608[0]};
    Full_Adder FA_15859(s15859, c15859, in15859_1, in15859_2, s15219[0]);
    wire[0:0] s15860, in15860_1, in15860_2;
    wire c15860;
    assign in15860_1 = {c15608};
    assign in15860_2 = {s15609[0]};
    Full_Adder FA_15860(s15860, c15860, in15860_1, in15860_2, s15221[0]);
    wire[0:0] s15861, in15861_1, in15861_2;
    wire c15861;
    assign in15861_1 = {c15609};
    assign in15861_2 = {s15610[0]};
    Full_Adder FA_15861(s15861, c15861, in15861_1, in15861_2, s15223[0]);
    wire[0:0] s15862, in15862_1, in15862_2;
    wire c15862;
    assign in15862_1 = {c15610};
    assign in15862_2 = {s15611[0]};
    Full_Adder FA_15862(s15862, c15862, in15862_1, in15862_2, s15225[0]);
    wire[0:0] s15863, in15863_1, in15863_2;
    wire c15863;
    assign in15863_1 = {c15611};
    assign in15863_2 = {s15612[0]};
    Full_Adder FA_15863(s15863, c15863, in15863_1, in15863_2, s15227[0]);
    wire[0:0] s15864, in15864_1, in15864_2;
    wire c15864;
    assign in15864_1 = {c15612};
    assign in15864_2 = {s15613[0]};
    Full_Adder FA_15864(s15864, c15864, in15864_1, in15864_2, s15229[0]);
    wire[0:0] s15865, in15865_1, in15865_2;
    wire c15865;
    assign in15865_1 = {c15613};
    assign in15865_2 = {s15614[0]};
    Full_Adder FA_15865(s15865, c15865, in15865_1, in15865_2, s15231[0]);
    wire[0:0] s15866, in15866_1, in15866_2;
    wire c15866;
    assign in15866_1 = {c15614};
    assign in15866_2 = {s15615[0]};
    Full_Adder FA_15866(s15866, c15866, in15866_1, in15866_2, s15233[0]);
    wire[0:0] s15867, in15867_1, in15867_2;
    wire c15867;
    assign in15867_1 = {c15615};
    assign in15867_2 = {s15616[0]};
    Full_Adder FA_15867(s15867, c15867, in15867_1, in15867_2, s15235[0]);
    wire[0:0] s15868, in15868_1, in15868_2;
    wire c15868;
    assign in15868_1 = {c15616};
    assign in15868_2 = {s15617[0]};
    Full_Adder FA_15868(s15868, c15868, in15868_1, in15868_2, s15237[0]);
    wire[0:0] s15869, in15869_1, in15869_2;
    wire c15869;
    assign in15869_1 = {c15617};
    assign in15869_2 = {s15618[0]};
    Full_Adder FA_15869(s15869, c15869, in15869_1, in15869_2, s15239[0]);
    wire[0:0] s15870, in15870_1, in15870_2;
    wire c15870;
    assign in15870_1 = {c15618};
    assign in15870_2 = {s15619[0]};
    Full_Adder FA_15870(s15870, c15870, in15870_1, in15870_2, s15241[0]);
    wire[0:0] s15871, in15871_1, in15871_2;
    wire c15871;
    assign in15871_1 = {c15619};
    assign in15871_2 = {s15620[0]};
    Full_Adder FA_15871(s15871, c15871, in15871_1, in15871_2, s15243[0]);
    wire[0:0] s15872, in15872_1, in15872_2;
    wire c15872;
    assign in15872_1 = {c15620};
    assign in15872_2 = {s15621[0]};
    Full_Adder FA_15872(s15872, c15872, in15872_1, in15872_2, s15245[0]);
    wire[0:0] s15873, in15873_1, in15873_2;
    wire c15873;
    assign in15873_1 = {c15621};
    assign in15873_2 = {s15622[0]};
    Full_Adder FA_15873(s15873, c15873, in15873_1, in15873_2, s15247[0]);
    wire[0:0] s15874, in15874_1, in15874_2;
    wire c15874;
    assign in15874_1 = {c15622};
    assign in15874_2 = {s15623[0]};
    Full_Adder FA_15874(s15874, c15874, in15874_1, in15874_2, s15249[0]);
    wire[0:0] s15875, in15875_1, in15875_2;
    wire c15875;
    assign in15875_1 = {c15623};
    assign in15875_2 = {s15624[0]};
    Full_Adder FA_15875(s15875, c15875, in15875_1, in15875_2, s15251[0]);
    wire[0:0] s15876, in15876_1, in15876_2;
    wire c15876;
    assign in15876_1 = {c15624};
    assign in15876_2 = {s15625[0]};
    Full_Adder FA_15876(s15876, c15876, in15876_1, in15876_2, s15253[0]);
    wire[0:0] s15877, in15877_1, in15877_2;
    wire c15877;
    assign in15877_1 = {c15625};
    assign in15877_2 = {s15626[0]};
    Full_Adder FA_15877(s15877, c15877, in15877_1, in15877_2, s15255[0]);
    wire[0:0] s15878, in15878_1, in15878_2;
    wire c15878;
    assign in15878_1 = {c15626};
    assign in15878_2 = {s15627[0]};
    Full_Adder FA_15878(s15878, c15878, in15878_1, in15878_2, s15257[0]);
    wire[0:0] s15879, in15879_1, in15879_2;
    wire c15879;
    assign in15879_1 = {c15627};
    assign in15879_2 = {s15628[0]};
    Full_Adder FA_15879(s15879, c15879, in15879_1, in15879_2, s15259[0]);
    wire[0:0] s15880, in15880_1, in15880_2;
    wire c15880;
    assign in15880_1 = {c15628};
    assign in15880_2 = {s15629[0]};
    Full_Adder FA_15880(s15880, c15880, in15880_1, in15880_2, s15261[0]);
    wire[0:0] s15881, in15881_1, in15881_2;
    wire c15881;
    assign in15881_1 = {c15629};
    assign in15881_2 = {s15630[0]};
    Full_Adder FA_15881(s15881, c15881, in15881_1, in15881_2, s15263[0]);
    wire[0:0] s15882, in15882_1, in15882_2;
    wire c15882;
    assign in15882_1 = {c15630};
    assign in15882_2 = {s15631[0]};
    Full_Adder FA_15882(s15882, c15882, in15882_1, in15882_2, s15265[0]);
    wire[0:0] s15883, in15883_1, in15883_2;
    wire c15883;
    assign in15883_1 = {c15631};
    assign in15883_2 = {s15632[0]};
    Full_Adder FA_15883(s15883, c15883, in15883_1, in15883_2, s15267[0]);
    wire[0:0] s15884, in15884_1, in15884_2;
    wire c15884;
    assign in15884_1 = {c15632};
    assign in15884_2 = {s15633[0]};
    Full_Adder FA_15884(s15884, c15884, in15884_1, in15884_2, s15269[0]);
    wire[0:0] s15885, in15885_1, in15885_2;
    wire c15885;
    assign in15885_1 = {c15633};
    assign in15885_2 = {s15634[0]};
    Full_Adder FA_15885(s15885, c15885, in15885_1, in15885_2, s15271[0]);
    wire[0:0] s15886, in15886_1, in15886_2;
    wire c15886;
    assign in15886_1 = {c15634};
    assign in15886_2 = {s15635[0]};
    Full_Adder FA_15886(s15886, c15886, in15886_1, in15886_2, s15273[0]);
    wire[0:0] s15887, in15887_1, in15887_2;
    wire c15887;
    assign in15887_1 = {c15635};
    assign in15887_2 = {s15636[0]};
    Full_Adder FA_15887(s15887, c15887, in15887_1, in15887_2, s15275[0]);
    wire[0:0] s15888, in15888_1, in15888_2;
    wire c15888;
    assign in15888_1 = {c15636};
    assign in15888_2 = {s15637[0]};
    Full_Adder FA_15888(s15888, c15888, in15888_1, in15888_2, s15277[0]);
    wire[0:0] s15889, in15889_1, in15889_2;
    wire c15889;
    assign in15889_1 = {c15637};
    assign in15889_2 = {s15638[0]};
    Full_Adder FA_15889(s15889, c15889, in15889_1, in15889_2, s15279[0]);
    wire[0:0] s15890, in15890_1, in15890_2;
    wire c15890;
    assign in15890_1 = {c15638};
    assign in15890_2 = {s15639[0]};
    Full_Adder FA_15890(s15890, c15890, in15890_1, in15890_2, s15281[0]);
    wire[0:0] s15891, in15891_1, in15891_2;
    wire c15891;
    assign in15891_1 = {c15639};
    assign in15891_2 = {s15640[0]};
    Full_Adder FA_15891(s15891, c15891, in15891_1, in15891_2, s15283[0]);
    wire[0:0] s15892, in15892_1, in15892_2;
    wire c15892;
    assign in15892_1 = {c15640};
    assign in15892_2 = {s15641[0]};
    Full_Adder FA_15892(s15892, c15892, in15892_1, in15892_2, s15285[0]);
    wire[0:0] s15893, in15893_1, in15893_2;
    wire c15893;
    assign in15893_1 = {c15641};
    assign in15893_2 = {s15642[0]};
    Full_Adder FA_15893(s15893, c15893, in15893_1, in15893_2, s15287[0]);
    wire[0:0] s15894, in15894_1, in15894_2;
    wire c15894;
    assign in15894_1 = {c15642};
    assign in15894_2 = {s15643[0]};
    Full_Adder FA_15894(s15894, c15894, in15894_1, in15894_2, s15289[0]);
    wire[0:0] s15895, in15895_1, in15895_2;
    wire c15895;
    assign in15895_1 = {c15643};
    assign in15895_2 = {s15644[0]};
    Full_Adder FA_15895(s15895, c15895, in15895_1, in15895_2, s15291[0]);
    wire[0:0] s15896, in15896_1, in15896_2;
    wire c15896;
    assign in15896_1 = {c15644};
    assign in15896_2 = {s15645[0]};
    Full_Adder FA_15896(s15896, c15896, in15896_1, in15896_2, s15293[0]);
    wire[0:0] s15897, in15897_1, in15897_2;
    wire c15897;
    assign in15897_1 = {c15645};
    assign in15897_2 = {s15646[0]};
    Full_Adder FA_15897(s15897, c15897, in15897_1, in15897_2, s15295[0]);
    wire[0:0] s15898, in15898_1, in15898_2;
    wire c15898;
    assign in15898_1 = {c15646};
    assign in15898_2 = {s15647[0]};
    Full_Adder FA_15898(s15898, c15898, in15898_1, in15898_2, s15297[0]);
    wire[0:0] s15899, in15899_1, in15899_2;
    wire c15899;
    assign in15899_1 = {c15647};
    assign in15899_2 = {s15648[0]};
    Full_Adder FA_15899(s15899, c15899, in15899_1, in15899_2, s15299[0]);
    wire[0:0] s15900, in15900_1, in15900_2;
    wire c15900;
    assign in15900_1 = {c15648};
    assign in15900_2 = {s15649[0]};
    Full_Adder FA_15900(s15900, c15900, in15900_1, in15900_2, s15301[0]);
    wire[0:0] s15901, in15901_1, in15901_2;
    wire c15901;
    assign in15901_1 = {c15649};
    assign in15901_2 = {s15650[0]};
    Full_Adder FA_15901(s15901, c15901, in15901_1, in15901_2, s15303[0]);
    wire[0:0] s15902, in15902_1, in15902_2;
    wire c15902;
    assign in15902_1 = {c15650};
    assign in15902_2 = {s15651[0]};
    Full_Adder FA_15902(s15902, c15902, in15902_1, in15902_2, s15305[0]);
    wire[0:0] s15903, in15903_1, in15903_2;
    wire c15903;
    assign in15903_1 = {c15651};
    assign in15903_2 = {s15652[0]};
    Full_Adder FA_15903(s15903, c15903, in15903_1, in15903_2, s15307[0]);
    wire[0:0] s15904, in15904_1, in15904_2;
    wire c15904;
    assign in15904_1 = {c15652};
    assign in15904_2 = {s15653[0]};
    Full_Adder FA_15904(s15904, c15904, in15904_1, in15904_2, s15309[0]);
    wire[0:0] s15905, in15905_1, in15905_2;
    wire c15905;
    assign in15905_1 = {c15653};
    assign in15905_2 = {s15654[0]};
    Full_Adder FA_15905(s15905, c15905, in15905_1, in15905_2, s15311[0]);
    wire[0:0] s15906, in15906_1, in15906_2;
    wire c15906;
    assign in15906_1 = {c15654};
    assign in15906_2 = {s15655[0]};
    Full_Adder FA_15906(s15906, c15906, in15906_1, in15906_2, s15313[0]);
    wire[0:0] s15907, in15907_1, in15907_2;
    wire c15907;
    assign in15907_1 = {c15655};
    assign in15907_2 = {s15656[0]};
    Full_Adder FA_15907(s15907, c15907, in15907_1, in15907_2, s15315[0]);
    wire[0:0] s15908, in15908_1, in15908_2;
    wire c15908;
    assign in15908_1 = {c15656};
    assign in15908_2 = {s15657[0]};
    Full_Adder FA_15908(s15908, c15908, in15908_1, in15908_2, s15317[0]);
    wire[0:0] s15909, in15909_1, in15909_2;
    wire c15909;
    assign in15909_1 = {c15657};
    assign in15909_2 = {s15658[0]};
    Full_Adder FA_15909(s15909, c15909, in15909_1, in15909_2, s15319[0]);
    wire[0:0] s15910, in15910_1, in15910_2;
    wire c15910;
    assign in15910_1 = {c15658};
    assign in15910_2 = {s15659[0]};
    Full_Adder FA_15910(s15910, c15910, in15910_1, in15910_2, s15321[0]);
    wire[0:0] s15911, in15911_1, in15911_2;
    wire c15911;
    assign in15911_1 = {c15659};
    assign in15911_2 = {s15660[0]};
    Full_Adder FA_15911(s15911, c15911, in15911_1, in15911_2, s15323[0]);
    wire[0:0] s15912, in15912_1, in15912_2;
    wire c15912;
    assign in15912_1 = {c15660};
    assign in15912_2 = {s15661[0]};
    Full_Adder FA_15912(s15912, c15912, in15912_1, in15912_2, s15325[0]);
    wire[0:0] s15913, in15913_1, in15913_2;
    wire c15913;
    assign in15913_1 = {c15661};
    assign in15913_2 = {s15662[0]};
    Full_Adder FA_15913(s15913, c15913, in15913_1, in15913_2, s15327[0]);
    wire[0:0] s15914, in15914_1, in15914_2;
    wire c15914;
    assign in15914_1 = {c15662};
    assign in15914_2 = {s15663[0]};
    Full_Adder FA_15914(s15914, c15914, in15914_1, in15914_2, s15329[0]);
    wire[0:0] s15915, in15915_1, in15915_2;
    wire c15915;
    assign in15915_1 = {c15663};
    assign in15915_2 = {s15664[0]};
    Full_Adder FA_15915(s15915, c15915, in15915_1, in15915_2, s15331[0]);
    wire[0:0] s15916, in15916_1, in15916_2;
    wire c15916;
    assign in15916_1 = {c15664};
    assign in15916_2 = {s15665[0]};
    Full_Adder FA_15916(s15916, c15916, in15916_1, in15916_2, s15333[0]);
    wire[0:0] s15917, in15917_1, in15917_2;
    wire c15917;
    assign in15917_1 = {c15665};
    assign in15917_2 = {s15666[0]};
    Full_Adder FA_15917(s15917, c15917, in15917_1, in15917_2, s15335[0]);
    wire[0:0] s15918, in15918_1, in15918_2;
    wire c15918;
    assign in15918_1 = {c15666};
    assign in15918_2 = {s15667[0]};
    Full_Adder FA_15918(s15918, c15918, in15918_1, in15918_2, s15337[0]);
    wire[0:0] s15919, in15919_1, in15919_2;
    wire c15919;
    assign in15919_1 = {c15667};
    assign in15919_2 = {s15668[0]};
    Full_Adder FA_15919(s15919, c15919, in15919_1, in15919_2, s15339[0]);
    wire[0:0] s15920, in15920_1, in15920_2;
    wire c15920;
    assign in15920_1 = {c15668};
    assign in15920_2 = {s15669[0]};
    Full_Adder FA_15920(s15920, c15920, in15920_1, in15920_2, s15341[0]);
    wire[0:0] s15921, in15921_1, in15921_2;
    wire c15921;
    assign in15921_1 = {c15669};
    assign in15921_2 = {s15670[0]};
    Full_Adder FA_15921(s15921, c15921, in15921_1, in15921_2, s15343[0]);
    wire[0:0] s15922, in15922_1, in15922_2;
    wire c15922;
    assign in15922_1 = {c15670};
    assign in15922_2 = {s15671[0]};
    Full_Adder FA_15922(s15922, c15922, in15922_1, in15922_2, s15345[0]);
    wire[0:0] s15923, in15923_1, in15923_2;
    wire c15923;
    assign in15923_1 = {c15671};
    assign in15923_2 = {s15672[0]};
    Full_Adder FA_15923(s15923, c15923, in15923_1, in15923_2, s15347[0]);
    wire[0:0] s15924, in15924_1, in15924_2;
    wire c15924;
    assign in15924_1 = {c15672};
    assign in15924_2 = {s15673[0]};
    Full_Adder FA_15924(s15924, c15924, in15924_1, in15924_2, s15349[0]);
    wire[0:0] s15925, in15925_1, in15925_2;
    wire c15925;
    assign in15925_1 = {c15673};
    assign in15925_2 = {s15674[0]};
    Full_Adder FA_15925(s15925, c15925, in15925_1, in15925_2, s15351[0]);
    wire[0:0] s15926, in15926_1, in15926_2;
    wire c15926;
    assign in15926_1 = {c15674};
    assign in15926_2 = {s15675[0]};
    Full_Adder FA_15926(s15926, c15926, in15926_1, in15926_2, s15353[0]);
    wire[0:0] s15927, in15927_1, in15927_2;
    wire c15927;
    assign in15927_1 = {c15675};
    assign in15927_2 = {s15676[0]};
    Full_Adder FA_15927(s15927, c15927, in15927_1, in15927_2, s15355[0]);
    wire[0:0] s15928, in15928_1, in15928_2;
    wire c15928;
    assign in15928_1 = {c15676};
    assign in15928_2 = {s15677[0]};
    Full_Adder FA_15928(s15928, c15928, in15928_1, in15928_2, s15357[0]);
    wire[0:0] s15929, in15929_1, in15929_2;
    wire c15929;
    assign in15929_1 = {c15677};
    assign in15929_2 = {s15678[0]};
    Full_Adder FA_15929(s15929, c15929, in15929_1, in15929_2, s15359[0]);
    wire[0:0] s15930, in15930_1, in15930_2;
    wire c15930;
    assign in15930_1 = {c15678};
    assign in15930_2 = {s15679[0]};
    Full_Adder FA_15930(s15930, c15930, in15930_1, in15930_2, s15361[0]);
    wire[0:0] s15931, in15931_1, in15931_2;
    wire c15931;
    assign in15931_1 = {c15679};
    assign in15931_2 = {s15680[0]};
    Full_Adder FA_15931(s15931, c15931, in15931_1, in15931_2, s15363[0]);
    wire[0:0] s15932, in15932_1, in15932_2;
    wire c15932;
    assign in15932_1 = {c15680};
    assign in15932_2 = {s15681[0]};
    Full_Adder FA_15932(s15932, c15932, in15932_1, in15932_2, s15365[0]);
    wire[0:0] s15933, in15933_1, in15933_2;
    wire c15933;
    assign in15933_1 = {c15681};
    assign in15933_2 = {s15682[0]};
    Full_Adder FA_15933(s15933, c15933, in15933_1, in15933_2, s15367[0]);
    wire[0:0] s15934, in15934_1, in15934_2;
    wire c15934;
    assign in15934_1 = {c15682};
    assign in15934_2 = {s15683[0]};
    Full_Adder FA_15934(s15934, c15934, in15934_1, in15934_2, s15369[0]);
    wire[0:0] s15935, in15935_1, in15935_2;
    wire c15935;
    assign in15935_1 = {c15683};
    assign in15935_2 = {s15684[0]};
    Full_Adder FA_15935(s15935, c15935, in15935_1, in15935_2, s15371[0]);
    wire[0:0] s15936, in15936_1, in15936_2;
    wire c15936;
    assign in15936_1 = {c15684};
    assign in15936_2 = {s15685[0]};
    Full_Adder FA_15936(s15936, c15936, in15936_1, in15936_2, s15373[0]);
    wire[0:0] s15937, in15937_1, in15937_2;
    wire c15937;
    assign in15937_1 = {c15685};
    assign in15937_2 = {s15686[0]};
    Full_Adder FA_15937(s15937, c15937, in15937_1, in15937_2, s15375[0]);
    wire[0:0] s15938, in15938_1, in15938_2;
    wire c15938;
    assign in15938_1 = {c15686};
    assign in15938_2 = {s15687[0]};
    Full_Adder FA_15938(s15938, c15938, in15938_1, in15938_2, s15377[0]);
    wire[0:0] s15939, in15939_1, in15939_2;
    wire c15939;
    assign in15939_1 = {c15687};
    assign in15939_2 = {s15688[0]};
    Full_Adder FA_15939(s15939, c15939, in15939_1, in15939_2, s15379[0]);
    wire[0:0] s15940, in15940_1, in15940_2;
    wire c15940;
    assign in15940_1 = {c15688};
    assign in15940_2 = {s15689[0]};
    Full_Adder FA_15940(s15940, c15940, in15940_1, in15940_2, s15381[0]);
    wire[0:0] s15941, in15941_1, in15941_2;
    wire c15941;
    assign in15941_1 = {c15689};
    assign in15941_2 = {s15690[0]};
    Full_Adder FA_15941(s15941, c15941, in15941_1, in15941_2, s15383[0]);
    wire[0:0] s15942, in15942_1, in15942_2;
    wire c15942;
    assign in15942_1 = {c15690};
    assign in15942_2 = {s15691[0]};
    Full_Adder FA_15942(s15942, c15942, in15942_1, in15942_2, s15385[0]);
    wire[0:0] s15943, in15943_1, in15943_2;
    wire c15943;
    assign in15943_1 = {c15691};
    assign in15943_2 = {s15692[0]};
    Full_Adder FA_15943(s15943, c15943, in15943_1, in15943_2, s15387[0]);
    wire[0:0] s15944, in15944_1, in15944_2;
    wire c15944;
    assign in15944_1 = {c15692};
    assign in15944_2 = {s15693[0]};
    Full_Adder FA_15944(s15944, c15944, in15944_1, in15944_2, s15389[0]);
    wire[0:0] s15945, in15945_1, in15945_2;
    wire c15945;
    assign in15945_1 = {c15693};
    assign in15945_2 = {s15694[0]};
    Full_Adder FA_15945(s15945, c15945, in15945_1, in15945_2, s15391[0]);
    wire[0:0] s15946, in15946_1, in15946_2;
    wire c15946;
    assign in15946_1 = {c15694};
    assign in15946_2 = {s15695[0]};
    Full_Adder FA_15946(s15946, c15946, in15946_1, in15946_2, s15393[0]);
    wire[0:0] s15947, in15947_1, in15947_2;
    wire c15947;
    assign in15947_1 = {c15695};
    assign in15947_2 = {s15696[0]};
    Full_Adder FA_15947(s15947, c15947, in15947_1, in15947_2, s15395[0]);
    wire[0:0] s15948, in15948_1, in15948_2;
    wire c15948;
    assign in15948_1 = {c15696};
    assign in15948_2 = {s15697[0]};
    Full_Adder FA_15948(s15948, c15948, in15948_1, in15948_2, s15397[0]);
    wire[0:0] s15949, in15949_1, in15949_2;
    wire c15949;
    assign in15949_1 = {c15697};
    assign in15949_2 = {s15698[0]};
    Full_Adder FA_15949(s15949, c15949, in15949_1, in15949_2, s15399[0]);
    wire[0:0] s15950, in15950_1, in15950_2;
    wire c15950;
    assign in15950_1 = {c15698};
    assign in15950_2 = {s15699[0]};
    Full_Adder FA_15950(s15950, c15950, in15950_1, in15950_2, s15401[0]);
    wire[0:0] s15951, in15951_1, in15951_2;
    wire c15951;
    assign in15951_1 = {c15699};
    assign in15951_2 = {s15700[0]};
    Full_Adder FA_15951(s15951, c15951, in15951_1, in15951_2, s15403[0]);
    wire[0:0] s15952, in15952_1, in15952_2;
    wire c15952;
    assign in15952_1 = {c15700};
    assign in15952_2 = {s15701[0]};
    Full_Adder FA_15952(s15952, c15952, in15952_1, in15952_2, s15405[0]);
    wire[0:0] s15953, in15953_1, in15953_2;
    wire c15953;
    assign in15953_1 = {c15701};
    assign in15953_2 = {s15702[0]};
    Full_Adder FA_15953(s15953, c15953, in15953_1, in15953_2, s15407[0]);
    wire[0:0] s15954, in15954_1, in15954_2;
    wire c15954;
    assign in15954_1 = {c15702};
    assign in15954_2 = {s15703[0]};
    Full_Adder FA_15954(s15954, c15954, in15954_1, in15954_2, s15409[0]);
    wire[0:0] s15955, in15955_1, in15955_2;
    wire c15955;
    assign in15955_1 = {c15703};
    assign in15955_2 = {s15704[0]};
    Full_Adder FA_15955(s15955, c15955, in15955_1, in15955_2, s15411[0]);
    wire[0:0] s15956, in15956_1, in15956_2;
    wire c15956;
    assign in15956_1 = {c15704};
    assign in15956_2 = {s15705[0]};
    Full_Adder FA_15956(s15956, c15956, in15956_1, in15956_2, s15413[0]);
    wire[0:0] s15957, in15957_1, in15957_2;
    wire c15957;
    assign in15957_1 = {c15705};
    assign in15957_2 = {s15706[0]};
    Full_Adder FA_15957(s15957, c15957, in15957_1, in15957_2, s15415[0]);
    wire[0:0] s15958, in15958_1, in15958_2;
    wire c15958;
    assign in15958_1 = {c15706};
    assign in15958_2 = {s15707[0]};
    Full_Adder FA_15958(s15958, c15958, in15958_1, in15958_2, s15417[0]);
    wire[0:0] s15959, in15959_1, in15959_2;
    wire c15959;
    assign in15959_1 = {c15707};
    assign in15959_2 = {s15708[0]};
    Full_Adder FA_15959(s15959, c15959, in15959_1, in15959_2, s15419[0]);
    wire[0:0] s15960, in15960_1, in15960_2;
    wire c15960;
    assign in15960_1 = {c15708};
    assign in15960_2 = {s15709[0]};
    Full_Adder FA_15960(s15960, c15960, in15960_1, in15960_2, s15421[0]);
    wire[0:0] s15961, in15961_1, in15961_2;
    wire c15961;
    assign in15961_1 = {c15709};
    assign in15961_2 = {s15710[0]};
    Full_Adder FA_15961(s15961, c15961, in15961_1, in15961_2, s15423[0]);
    wire[0:0] s15962, in15962_1, in15962_2;
    wire c15962;
    assign in15962_1 = {c15710};
    assign in15962_2 = {s15711[0]};
    Full_Adder FA_15962(s15962, c15962, in15962_1, in15962_2, s15425[0]);
    wire[0:0] s15963, in15963_1, in15963_2;
    wire c15963;
    assign in15963_1 = {c15711};
    assign in15963_2 = {s15712[0]};
    Full_Adder FA_15963(s15963, c15963, in15963_1, in15963_2, s15427[0]);
    wire[0:0] s15964, in15964_1, in15964_2;
    wire c15964;
    assign in15964_1 = {c15712};
    assign in15964_2 = {s15713[0]};
    Full_Adder FA_15964(s15964, c15964, in15964_1, in15964_2, s15429[0]);
    wire[0:0] s15965, in15965_1, in15965_2;
    wire c15965;
    assign in15965_1 = {c15713};
    assign in15965_2 = {s15714[0]};
    Full_Adder FA_15965(s15965, c15965, in15965_1, in15965_2, s15431[0]);
    wire[0:0] s15966, in15966_1, in15966_2;
    wire c15966;
    assign in15966_1 = {c15714};
    assign in15966_2 = {s15715[0]};
    Full_Adder FA_15966(s15966, c15966, in15966_1, in15966_2, s15433[0]);
    wire[0:0] s15967, in15967_1, in15967_2;
    wire c15967;
    assign in15967_1 = {c15715};
    assign in15967_2 = {s15716[0]};
    Full_Adder FA_15967(s15967, c15967, in15967_1, in15967_2, s15435[0]);
    wire[0:0] s15968, in15968_1, in15968_2;
    wire c15968;
    assign in15968_1 = {c15716};
    assign in15968_2 = {s15717[0]};
    Full_Adder FA_15968(s15968, c15968, in15968_1, in15968_2, s15437[0]);
    wire[0:0] s15969, in15969_1, in15969_2;
    wire c15969;
    assign in15969_1 = {c15717};
    assign in15969_2 = {s15718[0]};
    Full_Adder FA_15969(s15969, c15969, in15969_1, in15969_2, s15439[0]);
    wire[0:0] s15970, in15970_1, in15970_2;
    wire c15970;
    assign in15970_1 = {c15718};
    assign in15970_2 = {s15719[0]};
    Full_Adder FA_15970(s15970, c15970, in15970_1, in15970_2, s15441[0]);
    wire[0:0] s15971, in15971_1, in15971_2;
    wire c15971;
    assign in15971_1 = {c15719};
    assign in15971_2 = {s15720[0]};
    Full_Adder FA_15971(s15971, c15971, in15971_1, in15971_2, s15443[0]);
    wire[0:0] s15972, in15972_1, in15972_2;
    wire c15972;
    assign in15972_1 = {c15720};
    assign in15972_2 = {s15721[0]};
    Full_Adder FA_15972(s15972, c15972, in15972_1, in15972_2, s15445[0]);
    wire[0:0] s15973, in15973_1, in15973_2;
    wire c15973;
    assign in15973_1 = {c15721};
    assign in15973_2 = {s15722[0]};
    Full_Adder FA_15973(s15973, c15973, in15973_1, in15973_2, s15447[0]);
    wire[0:0] s15974, in15974_1, in15974_2;
    wire c15974;
    assign in15974_1 = {c15722};
    assign in15974_2 = {s15723[0]};
    Full_Adder FA_15974(s15974, c15974, in15974_1, in15974_2, s15449[0]);
    wire[0:0] s15975, in15975_1, in15975_2;
    wire c15975;
    assign in15975_1 = {c15723};
    assign in15975_2 = {s15724[0]};
    Full_Adder FA_15975(s15975, c15975, in15975_1, in15975_2, s15451[0]);
    wire[0:0] s15976, in15976_1, in15976_2;
    wire c15976;
    assign in15976_1 = {c15724};
    assign in15976_2 = {s15725[0]};
    Full_Adder FA_15976(s15976, c15976, in15976_1, in15976_2, s15453[0]);
    wire[0:0] s15977, in15977_1, in15977_2;
    wire c15977;
    assign in15977_1 = {c15725};
    assign in15977_2 = {s15726[0]};
    Full_Adder FA_15977(s15977, c15977, in15977_1, in15977_2, s15455[0]);
    wire[0:0] s15978, in15978_1, in15978_2;
    wire c15978;
    assign in15978_1 = {c15726};
    assign in15978_2 = {s15727[0]};
    Full_Adder FA_15978(s15978, c15978, in15978_1, in15978_2, s15457[0]);
    wire[0:0] s15979, in15979_1, in15979_2;
    wire c15979;
    assign in15979_1 = {c15727};
    assign in15979_2 = {s15728[0]};
    Full_Adder FA_15979(s15979, c15979, in15979_1, in15979_2, s15459[0]);
    wire[0:0] s15980, in15980_1, in15980_2;
    wire c15980;
    assign in15980_1 = {c15728};
    assign in15980_2 = {s15729[0]};
    Full_Adder FA_15980(s15980, c15980, in15980_1, in15980_2, s15461[0]);
    wire[0:0] s15981, in15981_1, in15981_2;
    wire c15981;
    assign in15981_1 = {c15729};
    assign in15981_2 = {s15730[0]};
    Full_Adder FA_15981(s15981, c15981, in15981_1, in15981_2, s15463[0]);
    wire[0:0] s15982, in15982_1, in15982_2;
    wire c15982;
    assign in15982_1 = {c15730};
    assign in15982_2 = {s15731[0]};
    Full_Adder FA_15982(s15982, c15982, in15982_1, in15982_2, s15465[0]);
    wire[0:0] s15983, in15983_1, in15983_2;
    wire c15983;
    assign in15983_1 = {c15731};
    assign in15983_2 = {s15732[0]};
    Full_Adder FA_15983(s15983, c15983, in15983_1, in15983_2, s15467[0]);
    wire[0:0] s15984, in15984_1, in15984_2;
    wire c15984;
    assign in15984_1 = {c15732};
    assign in15984_2 = {s15733[0]};
    Full_Adder FA_15984(s15984, c15984, in15984_1, in15984_2, s15469[0]);
    wire[0:0] s15985, in15985_1, in15985_2;
    wire c15985;
    assign in15985_1 = {c15733};
    assign in15985_2 = {s15734[0]};
    Full_Adder FA_15985(s15985, c15985, in15985_1, in15985_2, s15471[0]);
    wire[0:0] s15986, in15986_1, in15986_2;
    wire c15986;
    assign in15986_1 = {c15734};
    assign in15986_2 = {s15735[0]};
    Full_Adder FA_15986(s15986, c15986, in15986_1, in15986_2, s15473[0]);
    wire[0:0] s15987, in15987_1, in15987_2;
    wire c15987;
    assign in15987_1 = {c15735};
    assign in15987_2 = {s15736[0]};
    Full_Adder FA_15987(s15987, c15987, in15987_1, in15987_2, s15475[0]);
    wire[0:0] s15988, in15988_1, in15988_2;
    wire c15988;
    assign in15988_1 = {c15736};
    assign in15988_2 = {s15737[0]};
    Full_Adder FA_15988(s15988, c15988, in15988_1, in15988_2, s15477[0]);
    wire[0:0] s15989, in15989_1, in15989_2;
    wire c15989;
    assign in15989_1 = {c15737};
    assign in15989_2 = {s15738[0]};
    Full_Adder FA_15989(s15989, c15989, in15989_1, in15989_2, s15479[0]);
    wire[0:0] s15990, in15990_1, in15990_2;
    wire c15990;
    assign in15990_1 = {c15738};
    assign in15990_2 = {s15739[0]};
    Full_Adder FA_15990(s15990, c15990, in15990_1, in15990_2, s15481[0]);
    wire[0:0] s15991, in15991_1, in15991_2;
    wire c15991;
    assign in15991_1 = {c15739};
    assign in15991_2 = {s15740[0]};
    Full_Adder FA_15991(s15991, c15991, in15991_1, in15991_2, s15483[0]);
    wire[0:0] s15992, in15992_1, in15992_2;
    wire c15992;
    assign in15992_1 = {c15740};
    assign in15992_2 = {s15741[0]};
    Full_Adder FA_15992(s15992, c15992, in15992_1, in15992_2, s15485[0]);
    wire[0:0] s15993, in15993_1, in15993_2;
    wire c15993;
    assign in15993_1 = {c15741};
    assign in15993_2 = {s15742[0]};
    Full_Adder FA_15993(s15993, c15993, in15993_1, in15993_2, s15487[0]);
    wire[0:0] s15994, in15994_1, in15994_2;
    wire c15994;
    assign in15994_1 = {c15742};
    assign in15994_2 = {s15743[0]};
    Full_Adder FA_15994(s15994, c15994, in15994_1, in15994_2, s15489[0]);
    wire[0:0] s15995, in15995_1, in15995_2;
    wire c15995;
    assign in15995_1 = {c15743};
    assign in15995_2 = {s15744[0]};
    Full_Adder FA_15995(s15995, c15995, in15995_1, in15995_2, s15491[0]);
    wire[0:0] s15996, in15996_1, in15996_2;
    wire c15996;
    assign in15996_1 = {c15744};
    assign in15996_2 = {s15745[0]};
    Full_Adder FA_15996(s15996, c15996, in15996_1, in15996_2, s15493[0]);
    wire[0:0] s15997, in15997_1, in15997_2;
    wire c15997;
    assign in15997_1 = {c15745};
    assign in15997_2 = {s15746[0]};
    Full_Adder FA_15997(s15997, c15997, in15997_1, in15997_2, s15495[0]);
    wire[0:0] s15998, in15998_1, in15998_2;
    wire c15998;
    assign in15998_1 = {c15746};
    assign in15998_2 = {s15747[0]};
    Full_Adder FA_15998(s15998, c15998, in15998_1, in15998_2, s15497[0]);
    wire[0:0] s15999, in15999_1, in15999_2;
    wire c15999;
    assign in15999_1 = {c15747};
    assign in15999_2 = {s15748[0]};
    Full_Adder FA_15999(s15999, c15999, in15999_1, in15999_2, s15499[0]);
    wire[0:0] s16000, in16000_1, in16000_2;
    wire c16000;
    assign in16000_1 = {c15748};
    assign in16000_2 = {s15749[0]};
    Full_Adder FA_16000(s16000, c16000, in16000_1, in16000_2, s15500[0]);
    wire[0:0] s16001, in16001_1, in16001_2;
    wire c16001;
    assign in16001_1 = {c15749};
    assign in16001_2 = {s15750[0]};
    Full_Adder FA_16001(s16001, c16001, in16001_1, in16001_2, c15500);
    wire[0:0] s16002, in16002_1, in16002_2;
    wire c16002;
    assign in16002_1 = {pp127[126]};
    assign in16002_2 = {c15750};
    Full_Adder FA_16002(s16002, c16002, in16002_1, in16002_2, pp126[127]);


    /*Final Stage 11*/
    wire[253:0] s, in_1, in_2;
    wire c;
    assign in_1 = {pp0[1],pp2[0],c15751,c15752,c15753,c15754,c15755,c15756,c15757,c15758,c15759,c15760,c15761,c15762,c15763,c15764,c15765,c15766,c15767,c15768,c15769,c15770,c15771,c15772,c15773,c15774,c15775,c15776,c15777,c15778,c15779,c15780,c15781,c15782,c15783,c15784,c15785,c15786,c15787,c15788,c15789,c15790,c15791,c15792,c15793,c15794,c15795,c15796,c15797,c15798,c15799,c15800,c15801,c15802,c15803,c15804,c15805,c15806,c15807,c15808,c15809,c15810,c15811,c15812,c15813,c15814,c15815,c15816,c15817,c15818,c15819,c15820,c15821,c15822,c15823,c15824,c15825,c15826,c15827,c15828,c15829,c15830,c15831,c15832,c15833,c15834,c15835,c15836,c15837,c15838,c15839,c15840,c15841,c15842,c15843,c15844,c15845,c15846,c15847,c15848,c15849,c15850,c15851,c15852,c15853,c15854,c15855,c15856,c15857,c15858,c15859,c15860,c15861,c15862,c15863,c15864,c15865,c15866,c15867,c15868,c15869,c15870,c15871,c15872,c15873,c15874,c15875,c15876,c15877,c15878,c15879,c15880,c15881,c15882,c15883,c15884,c15885,c15886,c15887,c15888,c15889,c15890,c15891,c15892,c15893,c15894,c15895,c15896,c15897,c15898,c15899,c15900,c15901,c15902,c15903,c15904,c15905,c15906,c15907,c15908,c15909,c15910,c15911,c15912,c15913,c15914,c15915,c15916,c15917,c15918,c15919,c15920,c15921,c15922,c15923,c15924,c15925,c15926,c15927,c15928,c15929,c15930,c15931,c15932,c15933,c15934,c15935,c15936,c15937,c15938,c15939,c15940,c15941,c15942,c15943,c15944,c15945,c15946,c15947,c15948,c15949,c15950,c15951,c15952,c15953,c15954,c15955,c15956,c15957,c15958,c15959,c15960,c15961,c15962,c15963,c15964,c15965,c15966,c15967,c15968,c15969,c15970,c15971,c15972,c15973,c15974,c15975,c15976,c15977,c15978,c15979,c15980,c15981,c15982,c15983,c15984,c15985,c15986,c15987,c15988,c15989,c15990,c15991,c15992,c15993,c15994,c15995,c15996,c15997,c15998,c15999,c16000,c16001,pp127[127]};
    assign in_2 = {pp1[0],s15751[0],s15752[0],s15753[0],s15754[0],s15755[0],s15756[0],s15757[0],s15758[0],s15759[0],s15760[0],s15761[0],s15762[0],s15763[0],s15764[0],s15765[0],s15766[0],s15767[0],s15768[0],s15769[0],s15770[0],s15771[0],s15772[0],s15773[0],s15774[0],s15775[0],s15776[0],s15777[0],s15778[0],s15779[0],s15780[0],s15781[0],s15782[0],s15783[0],s15784[0],s15785[0],s15786[0],s15787[0],s15788[0],s15789[0],s15790[0],s15791[0],s15792[0],s15793[0],s15794[0],s15795[0],s15796[0],s15797[0],s15798[0],s15799[0],s15800[0],s15801[0],s15802[0],s15803[0],s15804[0],s15805[0],s15806[0],s15807[0],s15808[0],s15809[0],s15810[0],s15811[0],s15812[0],s15813[0],s15814[0],s15815[0],s15816[0],s15817[0],s15818[0],s15819[0],s15820[0],s15821[0],s15822[0],s15823[0],s15824[0],s15825[0],s15826[0],s15827[0],s15828[0],s15829[0],s15830[0],s15831[0],s15832[0],s15833[0],s15834[0],s15835[0],s15836[0],s15837[0],s15838[0],s15839[0],s15840[0],s15841[0],s15842[0],s15843[0],s15844[0],s15845[0],s15846[0],s15847[0],s15848[0],s15849[0],s15850[0],s15851[0],s15852[0],s15853[0],s15854[0],s15855[0],s15856[0],s15857[0],s15858[0],s15859[0],s15860[0],s15861[0],s15862[0],s15863[0],s15864[0],s15865[0],s15866[0],s15867[0],s15868[0],s15869[0],s15870[0],s15871[0],s15872[0],s15873[0],s15874[0],s15875[0],s15876[0],s15877[0],s15878[0],s15879[0],s15880[0],s15881[0],s15882[0],s15883[0],s15884[0],s15885[0],s15886[0],s15887[0],s15888[0],s15889[0],s15890[0],s15891[0],s15892[0],s15893[0],s15894[0],s15895[0],s15896[0],s15897[0],s15898[0],s15899[0],s15900[0],s15901[0],s15902[0],s15903[0],s15904[0],s15905[0],s15906[0],s15907[0],s15908[0],s15909[0],s15910[0],s15911[0],s15912[0],s15913[0],s15914[0],s15915[0],s15916[0],s15917[0],s15918[0],s15919[0],s15920[0],s15921[0],s15922[0],s15923[0],s15924[0],s15925[0],s15926[0],s15927[0],s15928[0],s15929[0],s15930[0],s15931[0],s15932[0],s15933[0],s15934[0],s15935[0],s15936[0],s15937[0],s15938[0],s15939[0],s15940[0],s15941[0],s15942[0],s15943[0],s15944[0],s15945[0],s15946[0],s15947[0],s15948[0],s15949[0],s15950[0],s15951[0],s15952[0],s15953[0],s15954[0],s15955[0],s15956[0],s15957[0],s15958[0],s15959[0],s15960[0],s15961[0],s15962[0],s15963[0],s15964[0],s15965[0],s15966[0],s15967[0],s15968[0],s15969[0],s15970[0],s15971[0],s15972[0],s15973[0],s15974[0],s15975[0],s15976[0],s15977[0],s15978[0],s15979[0],s15980[0],s15981[0],s15982[0],s15983[0],s15984[0],s15985[0],s15986[0],s15987[0],s15988[0],s15989[0],s15990[0],s15991[0],s15992[0],s15993[0],s15994[0],s15995[0],s15996[0],s15997[0],s15998[0],s15999[0],s16000[0],s16001[0],s16002[0],c16002};
    CLA_254(s, c, in_1, in_2);

    assign product[0] = pp0[0];
    assign product[1] = s[0];
    assign product[2] = s[1];
    assign product[3] = s[2];
    assign product[4] = s[3];
    assign product[5] = s[4];
    assign product[6] = s[5];
    assign product[7] = s[6];
    assign product[8] = s[7];
    assign product[9] = s[8];
    assign product[10] = s[9];
    assign product[11] = s[10];
    assign product[12] = s[11];
    assign product[13] = s[12];
    assign product[14] = s[13];
    assign product[15] = s[14];
    assign product[16] = s[15];
    assign product[17] = s[16];
    assign product[18] = s[17];
    assign product[19] = s[18];
    assign product[20] = s[19];
    assign product[21] = s[20];
    assign product[22] = s[21];
    assign product[23] = s[22];
    assign product[24] = s[23];
    assign product[25] = s[24];
    assign product[26] = s[25];
    assign product[27] = s[26];
    assign product[28] = s[27];
    assign product[29] = s[28];
    assign product[30] = s[29];
    assign product[31] = s[30];
    assign product[32] = s[31];
    assign product[33] = s[32];
    assign product[34] = s[33];
    assign product[35] = s[34];
    assign product[36] = s[35];
    assign product[37] = s[36];
    assign product[38] = s[37];
    assign product[39] = s[38];
    assign product[40] = s[39];
    assign product[41] = s[40];
    assign product[42] = s[41];
    assign product[43] = s[42];
    assign product[44] = s[43];
    assign product[45] = s[44];
    assign product[46] = s[45];
    assign product[47] = s[46];
    assign product[48] = s[47];
    assign product[49] = s[48];
    assign product[50] = s[49];
    assign product[51] = s[50];
    assign product[52] = s[51];
    assign product[53] = s[52];
    assign product[54] = s[53];
    assign product[55] = s[54];
    assign product[56] = s[55];
    assign product[57] = s[56];
    assign product[58] = s[57];
    assign product[59] = s[58];
    assign product[60] = s[59];
    assign product[61] = s[60];
    assign product[62] = s[61];
    assign product[63] = s[62];
    assign product[64] = s[63];
    assign product[65] = s[64];
    assign product[66] = s[65];
    assign product[67] = s[66];
    assign product[68] = s[67];
    assign product[69] = s[68];
    assign product[70] = s[69];
    assign product[71] = s[70];
    assign product[72] = s[71];
    assign product[73] = s[72];
    assign product[74] = s[73];
    assign product[75] = s[74];
    assign product[76] = s[75];
    assign product[77] = s[76];
    assign product[78] = s[77];
    assign product[79] = s[78];
    assign product[80] = s[79];
    assign product[81] = s[80];
    assign product[82] = s[81];
    assign product[83] = s[82];
    assign product[84] = s[83];
    assign product[85] = s[84];
    assign product[86] = s[85];
    assign product[87] = s[86];
    assign product[88] = s[87];
    assign product[89] = s[88];
    assign product[90] = s[89];
    assign product[91] = s[90];
    assign product[92] = s[91];
    assign product[93] = s[92];
    assign product[94] = s[93];
    assign product[95] = s[94];
    assign product[96] = s[95];
    assign product[97] = s[96];
    assign product[98] = s[97];
    assign product[99] = s[98];
    assign product[100] = s[99];
    assign product[101] = s[100];
    assign product[102] = s[101];
    assign product[103] = s[102];
    assign product[104] = s[103];
    assign product[105] = s[104];
    assign product[106] = s[105];
    assign product[107] = s[106];
    assign product[108] = s[107];
    assign product[109] = s[108];
    assign product[110] = s[109];
    assign product[111] = s[110];
    assign product[112] = s[111];
    assign product[113] = s[112];
    assign product[114] = s[113];
    assign product[115] = s[114];
    assign product[116] = s[115];
    assign product[117] = s[116];
    assign product[118] = s[117];
    assign product[119] = s[118];
    assign product[120] = s[119];
    assign product[121] = s[120];
    assign product[122] = s[121];
    assign product[123] = s[122];
    assign product[124] = s[123];
    assign product[125] = s[124];
    assign product[126] = s[125];
    assign product[127] = s[126];
    assign product[128] = s[127];
    assign product[129] = s[128];
    assign product[130] = s[129];
    assign product[131] = s[130];
    assign product[132] = s[131];
    assign product[133] = s[132];
    assign product[134] = s[133];
    assign product[135] = s[134];
    assign product[136] = s[135];
    assign product[137] = s[136];
    assign product[138] = s[137];
    assign product[139] = s[138];
    assign product[140] = s[139];
    assign product[141] = s[140];
    assign product[142] = s[141];
    assign product[143] = s[142];
    assign product[144] = s[143];
    assign product[145] = s[144];
    assign product[146] = s[145];
    assign product[147] = s[146];
    assign product[148] = s[147];
    assign product[149] = s[148];
    assign product[150] = s[149];
    assign product[151] = s[150];
    assign product[152] = s[151];
    assign product[153] = s[152];
    assign product[154] = s[153];
    assign product[155] = s[154];
    assign product[156] = s[155];
    assign product[157] = s[156];
    assign product[158] = s[157];
    assign product[159] = s[158];
    assign product[160] = s[159];
    assign product[161] = s[160];
    assign product[162] = s[161];
    assign product[163] = s[162];
    assign product[164] = s[163];
    assign product[165] = s[164];
    assign product[166] = s[165];
    assign product[167] = s[166];
    assign product[168] = s[167];
    assign product[169] = s[168];
    assign product[170] = s[169];
    assign product[171] = s[170];
    assign product[172] = s[171];
    assign product[173] = s[172];
    assign product[174] = s[173];
    assign product[175] = s[174];
    assign product[176] = s[175];
    assign product[177] = s[176];
    assign product[178] = s[177];
    assign product[179] = s[178];
    assign product[180] = s[179];
    assign product[181] = s[180];
    assign product[182] = s[181];
    assign product[183] = s[182];
    assign product[184] = s[183];
    assign product[185] = s[184];
    assign product[186] = s[185];
    assign product[187] = s[186];
    assign product[188] = s[187];
    assign product[189] = s[188];
    assign product[190] = s[189];
    assign product[191] = s[190];
    assign product[192] = s[191];
    assign product[193] = s[192];
    assign product[194] = s[193];
    assign product[195] = s[194];
    assign product[196] = s[195];
    assign product[197] = s[196];
    assign product[198] = s[197];
    assign product[199] = s[198];
    assign product[200] = s[199];
    assign product[201] = s[200];
    assign product[202] = s[201];
    assign product[203] = s[202];
    assign product[204] = s[203];
    assign product[205] = s[204];
    assign product[206] = s[205];
    assign product[207] = s[206];
    assign product[208] = s[207];
    assign product[209] = s[208];
    assign product[210] = s[209];
    assign product[211] = s[210];
    assign product[212] = s[211];
    assign product[213] = s[212];
    assign product[214] = s[213];
    assign product[215] = s[214];
    assign product[216] = s[215];
    assign product[217] = s[216];
    assign product[218] = s[217];
    assign product[219] = s[218];
    assign product[220] = s[219];
    assign product[221] = s[220];
    assign product[222] = s[221];
    assign product[223] = s[222];
    assign product[224] = s[223];
    assign product[225] = s[224];
    assign product[226] = s[225];
    assign product[227] = s[226];
    assign product[228] = s[227];
    assign product[229] = s[228];
    assign product[230] = s[229];
    assign product[231] = s[230];
    assign product[232] = s[231];
    assign product[233] = s[232];
    assign product[234] = s[233];
    assign product[235] = s[234];
    assign product[236] = s[235];
    assign product[237] = s[236];
    assign product[238] = s[237];
    assign product[239] = s[238];
    assign product[240] = s[239];
    assign product[241] = s[240];
    assign product[242] = s[241];
    assign product[243] = s[242];
    assign product[244] = s[243];
    assign product[245] = s[244];
    assign product[246] = s[245];
    assign product[247] = s[246];
    assign product[248] = s[247];
    assign product[249] = s[248];
    assign product[250] = s[249];
    assign product[251] = s[250];
    assign product[252] = s[251];
    assign product[253] = s[252];
    assign product[254] = s[253];
    assign product[255] = c;
endmodule

module Half_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2);
    xor(sum, in1, in2);
    and(cout, in1, in2);
endmodule

module Full_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2,
                  input wire cin);
    wire temp1;
    wire temp2;
    wire temp3;
    xor(sum, in1, in2, cin);
    and(temp1,in1,in2);
    and(temp2,in1,cin);
    and(temp3,in2,cin);
    or(cout,temp1,temp2,temp3);
endmodule


module CLA_254(output [253:0] sum, output cout, input [253:0] in1, input [253:0] in2);

    wire[253:0] G;
    wire[253:0] C;
    wire[253:0] P;

    assign G[0] = in1[253] & in2[253];
    assign P[0] = in1[253] ^ in2[253];
    assign G[1] = in1[252] & in2[252];
    assign P[1] = in1[252] ^ in2[252];
    assign G[2] = in1[251] & in2[251];
    assign P[2] = in1[251] ^ in2[251];
    assign G[3] = in1[250] & in2[250];
    assign P[3] = in1[250] ^ in2[250];
    assign G[4] = in1[249] & in2[249];
    assign P[4] = in1[249] ^ in2[249];
    assign G[5] = in1[248] & in2[248];
    assign P[5] = in1[248] ^ in2[248];
    assign G[6] = in1[247] & in2[247];
    assign P[6] = in1[247] ^ in2[247];
    assign G[7] = in1[246] & in2[246];
    assign P[7] = in1[246] ^ in2[246];
    assign G[8] = in1[245] & in2[245];
    assign P[8] = in1[245] ^ in2[245];
    assign G[9] = in1[244] & in2[244];
    assign P[9] = in1[244] ^ in2[244];
    assign G[10] = in1[243] & in2[243];
    assign P[10] = in1[243] ^ in2[243];
    assign G[11] = in1[242] & in2[242];
    assign P[11] = in1[242] ^ in2[242];
    assign G[12] = in1[241] & in2[241];
    assign P[12] = in1[241] ^ in2[241];
    assign G[13] = in1[240] & in2[240];
    assign P[13] = in1[240] ^ in2[240];
    assign G[14] = in1[239] & in2[239];
    assign P[14] = in1[239] ^ in2[239];
    assign G[15] = in1[238] & in2[238];
    assign P[15] = in1[238] ^ in2[238];
    assign G[16] = in1[237] & in2[237];
    assign P[16] = in1[237] ^ in2[237];
    assign G[17] = in1[236] & in2[236];
    assign P[17] = in1[236] ^ in2[236];
    assign G[18] = in1[235] & in2[235];
    assign P[18] = in1[235] ^ in2[235];
    assign G[19] = in1[234] & in2[234];
    assign P[19] = in1[234] ^ in2[234];
    assign G[20] = in1[233] & in2[233];
    assign P[20] = in1[233] ^ in2[233];
    assign G[21] = in1[232] & in2[232];
    assign P[21] = in1[232] ^ in2[232];
    assign G[22] = in1[231] & in2[231];
    assign P[22] = in1[231] ^ in2[231];
    assign G[23] = in1[230] & in2[230];
    assign P[23] = in1[230] ^ in2[230];
    assign G[24] = in1[229] & in2[229];
    assign P[24] = in1[229] ^ in2[229];
    assign G[25] = in1[228] & in2[228];
    assign P[25] = in1[228] ^ in2[228];
    assign G[26] = in1[227] & in2[227];
    assign P[26] = in1[227] ^ in2[227];
    assign G[27] = in1[226] & in2[226];
    assign P[27] = in1[226] ^ in2[226];
    assign G[28] = in1[225] & in2[225];
    assign P[28] = in1[225] ^ in2[225];
    assign G[29] = in1[224] & in2[224];
    assign P[29] = in1[224] ^ in2[224];
    assign G[30] = in1[223] & in2[223];
    assign P[30] = in1[223] ^ in2[223];
    assign G[31] = in1[222] & in2[222];
    assign P[31] = in1[222] ^ in2[222];
    assign G[32] = in1[221] & in2[221];
    assign P[32] = in1[221] ^ in2[221];
    assign G[33] = in1[220] & in2[220];
    assign P[33] = in1[220] ^ in2[220];
    assign G[34] = in1[219] & in2[219];
    assign P[34] = in1[219] ^ in2[219];
    assign G[35] = in1[218] & in2[218];
    assign P[35] = in1[218] ^ in2[218];
    assign G[36] = in1[217] & in2[217];
    assign P[36] = in1[217] ^ in2[217];
    assign G[37] = in1[216] & in2[216];
    assign P[37] = in1[216] ^ in2[216];
    assign G[38] = in1[215] & in2[215];
    assign P[38] = in1[215] ^ in2[215];
    assign G[39] = in1[214] & in2[214];
    assign P[39] = in1[214] ^ in2[214];
    assign G[40] = in1[213] & in2[213];
    assign P[40] = in1[213] ^ in2[213];
    assign G[41] = in1[212] & in2[212];
    assign P[41] = in1[212] ^ in2[212];
    assign G[42] = in1[211] & in2[211];
    assign P[42] = in1[211] ^ in2[211];
    assign G[43] = in1[210] & in2[210];
    assign P[43] = in1[210] ^ in2[210];
    assign G[44] = in1[209] & in2[209];
    assign P[44] = in1[209] ^ in2[209];
    assign G[45] = in1[208] & in2[208];
    assign P[45] = in1[208] ^ in2[208];
    assign G[46] = in1[207] & in2[207];
    assign P[46] = in1[207] ^ in2[207];
    assign G[47] = in1[206] & in2[206];
    assign P[47] = in1[206] ^ in2[206];
    assign G[48] = in1[205] & in2[205];
    assign P[48] = in1[205] ^ in2[205];
    assign G[49] = in1[204] & in2[204];
    assign P[49] = in1[204] ^ in2[204];
    assign G[50] = in1[203] & in2[203];
    assign P[50] = in1[203] ^ in2[203];
    assign G[51] = in1[202] & in2[202];
    assign P[51] = in1[202] ^ in2[202];
    assign G[52] = in1[201] & in2[201];
    assign P[52] = in1[201] ^ in2[201];
    assign G[53] = in1[200] & in2[200];
    assign P[53] = in1[200] ^ in2[200];
    assign G[54] = in1[199] & in2[199];
    assign P[54] = in1[199] ^ in2[199];
    assign G[55] = in1[198] & in2[198];
    assign P[55] = in1[198] ^ in2[198];
    assign G[56] = in1[197] & in2[197];
    assign P[56] = in1[197] ^ in2[197];
    assign G[57] = in1[196] & in2[196];
    assign P[57] = in1[196] ^ in2[196];
    assign G[58] = in1[195] & in2[195];
    assign P[58] = in1[195] ^ in2[195];
    assign G[59] = in1[194] & in2[194];
    assign P[59] = in1[194] ^ in2[194];
    assign G[60] = in1[193] & in2[193];
    assign P[60] = in1[193] ^ in2[193];
    assign G[61] = in1[192] & in2[192];
    assign P[61] = in1[192] ^ in2[192];
    assign G[62] = in1[191] & in2[191];
    assign P[62] = in1[191] ^ in2[191];
    assign G[63] = in1[190] & in2[190];
    assign P[63] = in1[190] ^ in2[190];
    assign G[64] = in1[189] & in2[189];
    assign P[64] = in1[189] ^ in2[189];
    assign G[65] = in1[188] & in2[188];
    assign P[65] = in1[188] ^ in2[188];
    assign G[66] = in1[187] & in2[187];
    assign P[66] = in1[187] ^ in2[187];
    assign G[67] = in1[186] & in2[186];
    assign P[67] = in1[186] ^ in2[186];
    assign G[68] = in1[185] & in2[185];
    assign P[68] = in1[185] ^ in2[185];
    assign G[69] = in1[184] & in2[184];
    assign P[69] = in1[184] ^ in2[184];
    assign G[70] = in1[183] & in2[183];
    assign P[70] = in1[183] ^ in2[183];
    assign G[71] = in1[182] & in2[182];
    assign P[71] = in1[182] ^ in2[182];
    assign G[72] = in1[181] & in2[181];
    assign P[72] = in1[181] ^ in2[181];
    assign G[73] = in1[180] & in2[180];
    assign P[73] = in1[180] ^ in2[180];
    assign G[74] = in1[179] & in2[179];
    assign P[74] = in1[179] ^ in2[179];
    assign G[75] = in1[178] & in2[178];
    assign P[75] = in1[178] ^ in2[178];
    assign G[76] = in1[177] & in2[177];
    assign P[76] = in1[177] ^ in2[177];
    assign G[77] = in1[176] & in2[176];
    assign P[77] = in1[176] ^ in2[176];
    assign G[78] = in1[175] & in2[175];
    assign P[78] = in1[175] ^ in2[175];
    assign G[79] = in1[174] & in2[174];
    assign P[79] = in1[174] ^ in2[174];
    assign G[80] = in1[173] & in2[173];
    assign P[80] = in1[173] ^ in2[173];
    assign G[81] = in1[172] & in2[172];
    assign P[81] = in1[172] ^ in2[172];
    assign G[82] = in1[171] & in2[171];
    assign P[82] = in1[171] ^ in2[171];
    assign G[83] = in1[170] & in2[170];
    assign P[83] = in1[170] ^ in2[170];
    assign G[84] = in1[169] & in2[169];
    assign P[84] = in1[169] ^ in2[169];
    assign G[85] = in1[168] & in2[168];
    assign P[85] = in1[168] ^ in2[168];
    assign G[86] = in1[167] & in2[167];
    assign P[86] = in1[167] ^ in2[167];
    assign G[87] = in1[166] & in2[166];
    assign P[87] = in1[166] ^ in2[166];
    assign G[88] = in1[165] & in2[165];
    assign P[88] = in1[165] ^ in2[165];
    assign G[89] = in1[164] & in2[164];
    assign P[89] = in1[164] ^ in2[164];
    assign G[90] = in1[163] & in2[163];
    assign P[90] = in1[163] ^ in2[163];
    assign G[91] = in1[162] & in2[162];
    assign P[91] = in1[162] ^ in2[162];
    assign G[92] = in1[161] & in2[161];
    assign P[92] = in1[161] ^ in2[161];
    assign G[93] = in1[160] & in2[160];
    assign P[93] = in1[160] ^ in2[160];
    assign G[94] = in1[159] & in2[159];
    assign P[94] = in1[159] ^ in2[159];
    assign G[95] = in1[158] & in2[158];
    assign P[95] = in1[158] ^ in2[158];
    assign G[96] = in1[157] & in2[157];
    assign P[96] = in1[157] ^ in2[157];
    assign G[97] = in1[156] & in2[156];
    assign P[97] = in1[156] ^ in2[156];
    assign G[98] = in1[155] & in2[155];
    assign P[98] = in1[155] ^ in2[155];
    assign G[99] = in1[154] & in2[154];
    assign P[99] = in1[154] ^ in2[154];
    assign G[100] = in1[153] & in2[153];
    assign P[100] = in1[153] ^ in2[153];
    assign G[101] = in1[152] & in2[152];
    assign P[101] = in1[152] ^ in2[152];
    assign G[102] = in1[151] & in2[151];
    assign P[102] = in1[151] ^ in2[151];
    assign G[103] = in1[150] & in2[150];
    assign P[103] = in1[150] ^ in2[150];
    assign G[104] = in1[149] & in2[149];
    assign P[104] = in1[149] ^ in2[149];
    assign G[105] = in1[148] & in2[148];
    assign P[105] = in1[148] ^ in2[148];
    assign G[106] = in1[147] & in2[147];
    assign P[106] = in1[147] ^ in2[147];
    assign G[107] = in1[146] & in2[146];
    assign P[107] = in1[146] ^ in2[146];
    assign G[108] = in1[145] & in2[145];
    assign P[108] = in1[145] ^ in2[145];
    assign G[109] = in1[144] & in2[144];
    assign P[109] = in1[144] ^ in2[144];
    assign G[110] = in1[143] & in2[143];
    assign P[110] = in1[143] ^ in2[143];
    assign G[111] = in1[142] & in2[142];
    assign P[111] = in1[142] ^ in2[142];
    assign G[112] = in1[141] & in2[141];
    assign P[112] = in1[141] ^ in2[141];
    assign G[113] = in1[140] & in2[140];
    assign P[113] = in1[140] ^ in2[140];
    assign G[114] = in1[139] & in2[139];
    assign P[114] = in1[139] ^ in2[139];
    assign G[115] = in1[138] & in2[138];
    assign P[115] = in1[138] ^ in2[138];
    assign G[116] = in1[137] & in2[137];
    assign P[116] = in1[137] ^ in2[137];
    assign G[117] = in1[136] & in2[136];
    assign P[117] = in1[136] ^ in2[136];
    assign G[118] = in1[135] & in2[135];
    assign P[118] = in1[135] ^ in2[135];
    assign G[119] = in1[134] & in2[134];
    assign P[119] = in1[134] ^ in2[134];
    assign G[120] = in1[133] & in2[133];
    assign P[120] = in1[133] ^ in2[133];
    assign G[121] = in1[132] & in2[132];
    assign P[121] = in1[132] ^ in2[132];
    assign G[122] = in1[131] & in2[131];
    assign P[122] = in1[131] ^ in2[131];
    assign G[123] = in1[130] & in2[130];
    assign P[123] = in1[130] ^ in2[130];
    assign G[124] = in1[129] & in2[129];
    assign P[124] = in1[129] ^ in2[129];
    assign G[125] = in1[128] & in2[128];
    assign P[125] = in1[128] ^ in2[128];
    assign G[126] = in1[127] & in2[127];
    assign P[126] = in1[127] ^ in2[127];
    assign G[127] = in1[126] & in2[126];
    assign P[127] = in1[126] ^ in2[126];
    assign G[128] = in1[125] & in2[125];
    assign P[128] = in1[125] ^ in2[125];
    assign G[129] = in1[124] & in2[124];
    assign P[129] = in1[124] ^ in2[124];
    assign G[130] = in1[123] & in2[123];
    assign P[130] = in1[123] ^ in2[123];
    assign G[131] = in1[122] & in2[122];
    assign P[131] = in1[122] ^ in2[122];
    assign G[132] = in1[121] & in2[121];
    assign P[132] = in1[121] ^ in2[121];
    assign G[133] = in1[120] & in2[120];
    assign P[133] = in1[120] ^ in2[120];
    assign G[134] = in1[119] & in2[119];
    assign P[134] = in1[119] ^ in2[119];
    assign G[135] = in1[118] & in2[118];
    assign P[135] = in1[118] ^ in2[118];
    assign G[136] = in1[117] & in2[117];
    assign P[136] = in1[117] ^ in2[117];
    assign G[137] = in1[116] & in2[116];
    assign P[137] = in1[116] ^ in2[116];
    assign G[138] = in1[115] & in2[115];
    assign P[138] = in1[115] ^ in2[115];
    assign G[139] = in1[114] & in2[114];
    assign P[139] = in1[114] ^ in2[114];
    assign G[140] = in1[113] & in2[113];
    assign P[140] = in1[113] ^ in2[113];
    assign G[141] = in1[112] & in2[112];
    assign P[141] = in1[112] ^ in2[112];
    assign G[142] = in1[111] & in2[111];
    assign P[142] = in1[111] ^ in2[111];
    assign G[143] = in1[110] & in2[110];
    assign P[143] = in1[110] ^ in2[110];
    assign G[144] = in1[109] & in2[109];
    assign P[144] = in1[109] ^ in2[109];
    assign G[145] = in1[108] & in2[108];
    assign P[145] = in1[108] ^ in2[108];
    assign G[146] = in1[107] & in2[107];
    assign P[146] = in1[107] ^ in2[107];
    assign G[147] = in1[106] & in2[106];
    assign P[147] = in1[106] ^ in2[106];
    assign G[148] = in1[105] & in2[105];
    assign P[148] = in1[105] ^ in2[105];
    assign G[149] = in1[104] & in2[104];
    assign P[149] = in1[104] ^ in2[104];
    assign G[150] = in1[103] & in2[103];
    assign P[150] = in1[103] ^ in2[103];
    assign G[151] = in1[102] & in2[102];
    assign P[151] = in1[102] ^ in2[102];
    assign G[152] = in1[101] & in2[101];
    assign P[152] = in1[101] ^ in2[101];
    assign G[153] = in1[100] & in2[100];
    assign P[153] = in1[100] ^ in2[100];
    assign G[154] = in1[99] & in2[99];
    assign P[154] = in1[99] ^ in2[99];
    assign G[155] = in1[98] & in2[98];
    assign P[155] = in1[98] ^ in2[98];
    assign G[156] = in1[97] & in2[97];
    assign P[156] = in1[97] ^ in2[97];
    assign G[157] = in1[96] & in2[96];
    assign P[157] = in1[96] ^ in2[96];
    assign G[158] = in1[95] & in2[95];
    assign P[158] = in1[95] ^ in2[95];
    assign G[159] = in1[94] & in2[94];
    assign P[159] = in1[94] ^ in2[94];
    assign G[160] = in1[93] & in2[93];
    assign P[160] = in1[93] ^ in2[93];
    assign G[161] = in1[92] & in2[92];
    assign P[161] = in1[92] ^ in2[92];
    assign G[162] = in1[91] & in2[91];
    assign P[162] = in1[91] ^ in2[91];
    assign G[163] = in1[90] & in2[90];
    assign P[163] = in1[90] ^ in2[90];
    assign G[164] = in1[89] & in2[89];
    assign P[164] = in1[89] ^ in2[89];
    assign G[165] = in1[88] & in2[88];
    assign P[165] = in1[88] ^ in2[88];
    assign G[166] = in1[87] & in2[87];
    assign P[166] = in1[87] ^ in2[87];
    assign G[167] = in1[86] & in2[86];
    assign P[167] = in1[86] ^ in2[86];
    assign G[168] = in1[85] & in2[85];
    assign P[168] = in1[85] ^ in2[85];
    assign G[169] = in1[84] & in2[84];
    assign P[169] = in1[84] ^ in2[84];
    assign G[170] = in1[83] & in2[83];
    assign P[170] = in1[83] ^ in2[83];
    assign G[171] = in1[82] & in2[82];
    assign P[171] = in1[82] ^ in2[82];
    assign G[172] = in1[81] & in2[81];
    assign P[172] = in1[81] ^ in2[81];
    assign G[173] = in1[80] & in2[80];
    assign P[173] = in1[80] ^ in2[80];
    assign G[174] = in1[79] & in2[79];
    assign P[174] = in1[79] ^ in2[79];
    assign G[175] = in1[78] & in2[78];
    assign P[175] = in1[78] ^ in2[78];
    assign G[176] = in1[77] & in2[77];
    assign P[176] = in1[77] ^ in2[77];
    assign G[177] = in1[76] & in2[76];
    assign P[177] = in1[76] ^ in2[76];
    assign G[178] = in1[75] & in2[75];
    assign P[178] = in1[75] ^ in2[75];
    assign G[179] = in1[74] & in2[74];
    assign P[179] = in1[74] ^ in2[74];
    assign G[180] = in1[73] & in2[73];
    assign P[180] = in1[73] ^ in2[73];
    assign G[181] = in1[72] & in2[72];
    assign P[181] = in1[72] ^ in2[72];
    assign G[182] = in1[71] & in2[71];
    assign P[182] = in1[71] ^ in2[71];
    assign G[183] = in1[70] & in2[70];
    assign P[183] = in1[70] ^ in2[70];
    assign G[184] = in1[69] & in2[69];
    assign P[184] = in1[69] ^ in2[69];
    assign G[185] = in1[68] & in2[68];
    assign P[185] = in1[68] ^ in2[68];
    assign G[186] = in1[67] & in2[67];
    assign P[186] = in1[67] ^ in2[67];
    assign G[187] = in1[66] & in2[66];
    assign P[187] = in1[66] ^ in2[66];
    assign G[188] = in1[65] & in2[65];
    assign P[188] = in1[65] ^ in2[65];
    assign G[189] = in1[64] & in2[64];
    assign P[189] = in1[64] ^ in2[64];
    assign G[190] = in1[63] & in2[63];
    assign P[190] = in1[63] ^ in2[63];
    assign G[191] = in1[62] & in2[62];
    assign P[191] = in1[62] ^ in2[62];
    assign G[192] = in1[61] & in2[61];
    assign P[192] = in1[61] ^ in2[61];
    assign G[193] = in1[60] & in2[60];
    assign P[193] = in1[60] ^ in2[60];
    assign G[194] = in1[59] & in2[59];
    assign P[194] = in1[59] ^ in2[59];
    assign G[195] = in1[58] & in2[58];
    assign P[195] = in1[58] ^ in2[58];
    assign G[196] = in1[57] & in2[57];
    assign P[196] = in1[57] ^ in2[57];
    assign G[197] = in1[56] & in2[56];
    assign P[197] = in1[56] ^ in2[56];
    assign G[198] = in1[55] & in2[55];
    assign P[198] = in1[55] ^ in2[55];
    assign G[199] = in1[54] & in2[54];
    assign P[199] = in1[54] ^ in2[54];
    assign G[200] = in1[53] & in2[53];
    assign P[200] = in1[53] ^ in2[53];
    assign G[201] = in1[52] & in2[52];
    assign P[201] = in1[52] ^ in2[52];
    assign G[202] = in1[51] & in2[51];
    assign P[202] = in1[51] ^ in2[51];
    assign G[203] = in1[50] & in2[50];
    assign P[203] = in1[50] ^ in2[50];
    assign G[204] = in1[49] & in2[49];
    assign P[204] = in1[49] ^ in2[49];
    assign G[205] = in1[48] & in2[48];
    assign P[205] = in1[48] ^ in2[48];
    assign G[206] = in1[47] & in2[47];
    assign P[206] = in1[47] ^ in2[47];
    assign G[207] = in1[46] & in2[46];
    assign P[207] = in1[46] ^ in2[46];
    assign G[208] = in1[45] & in2[45];
    assign P[208] = in1[45] ^ in2[45];
    assign G[209] = in1[44] & in2[44];
    assign P[209] = in1[44] ^ in2[44];
    assign G[210] = in1[43] & in2[43];
    assign P[210] = in1[43] ^ in2[43];
    assign G[211] = in1[42] & in2[42];
    assign P[211] = in1[42] ^ in2[42];
    assign G[212] = in1[41] & in2[41];
    assign P[212] = in1[41] ^ in2[41];
    assign G[213] = in1[40] & in2[40];
    assign P[213] = in1[40] ^ in2[40];
    assign G[214] = in1[39] & in2[39];
    assign P[214] = in1[39] ^ in2[39];
    assign G[215] = in1[38] & in2[38];
    assign P[215] = in1[38] ^ in2[38];
    assign G[216] = in1[37] & in2[37];
    assign P[216] = in1[37] ^ in2[37];
    assign G[217] = in1[36] & in2[36];
    assign P[217] = in1[36] ^ in2[36];
    assign G[218] = in1[35] & in2[35];
    assign P[218] = in1[35] ^ in2[35];
    assign G[219] = in1[34] & in2[34];
    assign P[219] = in1[34] ^ in2[34];
    assign G[220] = in1[33] & in2[33];
    assign P[220] = in1[33] ^ in2[33];
    assign G[221] = in1[32] & in2[32];
    assign P[221] = in1[32] ^ in2[32];
    assign G[222] = in1[31] & in2[31];
    assign P[222] = in1[31] ^ in2[31];
    assign G[223] = in1[30] & in2[30];
    assign P[223] = in1[30] ^ in2[30];
    assign G[224] = in1[29] & in2[29];
    assign P[224] = in1[29] ^ in2[29];
    assign G[225] = in1[28] & in2[28];
    assign P[225] = in1[28] ^ in2[28];
    assign G[226] = in1[27] & in2[27];
    assign P[226] = in1[27] ^ in2[27];
    assign G[227] = in1[26] & in2[26];
    assign P[227] = in1[26] ^ in2[26];
    assign G[228] = in1[25] & in2[25];
    assign P[228] = in1[25] ^ in2[25];
    assign G[229] = in1[24] & in2[24];
    assign P[229] = in1[24] ^ in2[24];
    assign G[230] = in1[23] & in2[23];
    assign P[230] = in1[23] ^ in2[23];
    assign G[231] = in1[22] & in2[22];
    assign P[231] = in1[22] ^ in2[22];
    assign G[232] = in1[21] & in2[21];
    assign P[232] = in1[21] ^ in2[21];
    assign G[233] = in1[20] & in2[20];
    assign P[233] = in1[20] ^ in2[20];
    assign G[234] = in1[19] & in2[19];
    assign P[234] = in1[19] ^ in2[19];
    assign G[235] = in1[18] & in2[18];
    assign P[235] = in1[18] ^ in2[18];
    assign G[236] = in1[17] & in2[17];
    assign P[236] = in1[17] ^ in2[17];
    assign G[237] = in1[16] & in2[16];
    assign P[237] = in1[16] ^ in2[16];
    assign G[238] = in1[15] & in2[15];
    assign P[238] = in1[15] ^ in2[15];
    assign G[239] = in1[14] & in2[14];
    assign P[239] = in1[14] ^ in2[14];
    assign G[240] = in1[13] & in2[13];
    assign P[240] = in1[13] ^ in2[13];
    assign G[241] = in1[12] & in2[12];
    assign P[241] = in1[12] ^ in2[12];
    assign G[242] = in1[11] & in2[11];
    assign P[242] = in1[11] ^ in2[11];
    assign G[243] = in1[10] & in2[10];
    assign P[243] = in1[10] ^ in2[10];
    assign G[244] = in1[9] & in2[9];
    assign P[244] = in1[9] ^ in2[9];
    assign G[245] = in1[8] & in2[8];
    assign P[245] = in1[8] ^ in2[8];
    assign G[246] = in1[7] & in2[7];
    assign P[246] = in1[7] ^ in2[7];
    assign G[247] = in1[6] & in2[6];
    assign P[247] = in1[6] ^ in2[6];
    assign G[248] = in1[5] & in2[5];
    assign P[248] = in1[5] ^ in2[5];
    assign G[249] = in1[4] & in2[4];
    assign P[249] = in1[4] ^ in2[4];
    assign G[250] = in1[3] & in2[3];
    assign P[250] = in1[3] ^ in2[3];
    assign G[251] = in1[2] & in2[2];
    assign P[251] = in1[2] ^ in2[2];
    assign G[252] = in1[1] & in2[1];
    assign P[252] = in1[1] ^ in2[1];
    assign G[253] = in1[0] & in2[0];
    assign P[253] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign C[243] = G[242] | (P[242] & C[242]);
    assign C[244] = G[243] | (P[243] & C[243]);
    assign C[245] = G[244] | (P[244] & C[244]);
    assign C[246] = G[245] | (P[245] & C[245]);
    assign C[247] = G[246] | (P[246] & C[246]);
    assign C[248] = G[247] | (P[247] & C[247]);
    assign C[249] = G[248] | (P[248] & C[248]);
    assign C[250] = G[249] | (P[249] & C[249]);
    assign C[251] = G[250] | (P[250] & C[250]);
    assign C[252] = G[251] | (P[251] & C[251]);
    assign C[253] = G[252] | (P[252] & C[252]);
    assign cout = G[253] | (P[253] & C[253]);
    assign sum = P ^ C;
endmodule


